magic
tech sky130A
magscale 1 2
timestamp 1768990256
<< error_s >>
rect 3300 7342 10218 7346
rect 3300 5334 3330 7342
rect 3366 7276 3732 7280
rect 3794 7276 4160 7280
rect 4222 7276 4588 7280
rect 4650 7276 5016 7280
rect 5078 7276 5444 7280
rect 5506 7276 5872 7280
rect 5934 7276 6300 7280
rect 6362 7276 6728 7280
rect 6790 7276 7156 7280
rect 7218 7276 7584 7280
rect 7646 7276 8012 7280
rect 8074 7276 8440 7280
rect 8502 7276 8868 7280
rect 8930 7276 9296 7280
rect 9358 7276 9724 7280
rect 9786 7276 10152 7280
rect 3366 5400 3396 7276
rect 10122 5400 10152 7276
rect 10188 5334 10218 7342
rect 12200 6762 19118 6766
rect 12200 4634 12230 6762
rect 12266 6696 12632 6700
rect 12694 6696 13060 6700
rect 13122 6696 13488 6700
rect 13550 6696 13916 6700
rect 13978 6696 14344 6700
rect 14406 6696 14772 6700
rect 14834 6696 15200 6700
rect 15262 6696 15628 6700
rect 15690 6696 16056 6700
rect 16118 6696 16484 6700
rect 16546 6696 16912 6700
rect 16974 6696 17340 6700
rect 17402 6696 17768 6700
rect 17830 6696 18196 6700
rect 18258 6696 18624 6700
rect 18686 6696 19052 6700
rect 12266 4700 12296 6696
rect 19022 4700 19052 6696
rect 19088 4634 19118 6762
<< locali >>
rect 4000 4000 10100 4300
rect 4000 500 4300 4000
rect 6900 500 7300 4000
rect 9800 500 10100 4000
rect 1200 200 12800 500
rect 1200 -1800 1500 200
rect 12500 -1800 12800 200
rect 1200 -2100 12800 -1800
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__cap_mim_m3_1_RK594X  sky130_fd_pr__cap_mim_m3_1_RK594X_0
timestamp 1768989049
transform 1 0 -6508 0 1 3320
box -5492 -5320 5492 5320
use sky130_fd_pr__cap_mim_m3_1_RK594X  sky130_fd_pr__cap_mim_m3_1_RK594X_1
timestamp 1768989049
transform 1 0 23492 0 1 3320
box -5492 -5320 5492 5320
use sky130_fd_pr__nfet_g5v0d10v5_B9VV4Y  sky130_fd_pr__nfet_g5v0d10v5_B9VV4Y_0
timestamp 1768990256
transform 1 0 5525 0 1 3428
box -525 -528 525 528
use sky130_fd_pr__nfet_g5v0d10v5_B9VV4Y  sky130_fd_pr__nfet_g5v0d10v5_B9VV4Y_1
timestamp 1768990256
transform 1 0 8525 0 1 3428
box -525 -528 525 528
use sky130_fd_pr__nfet_g5v0d10v5_TJAW4Y  sky130_fd_pr__nfet_g5v0d10v5_TJAW4Y_0
timestamp 1768990256
transform 1 0 8525 0 1 1428
box -525 -528 525 528
use sky130_fd_pr__pfet_g5v0d10v5_HCTFFM  XM2
timestamp 1768990256
transform 1 0 6759 0 1 6304
box -3459 -1004 3459 1042
use sky130_fd_pr__nfet_g5v0d10v5_TJAW4Y  XM3
timestamp 1768990256
transform 1 0 5525 0 1 1428
box -525 -528 525 528
use sky130_fd_pr__nfet_g5v0d10v5_23PDXH  XM5
timestamp 1768990256
transform 1 0 7005 0 1 -793
box -5105 -807 5105 807
use sky130_fd_pr__pfet_g5v0d10v5_H6T99K  XM7
timestamp 1768990256
transform 1 0 15659 0 1 5664
box -3459 -1064 3459 1102
use sky130_fd_pr__pfet_g5v0d10v5_X45ZZ5  XM9
timestamp 1768989049
transform 1 0 17705 0 1 -4203
box -705 -797 705 797
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VP
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VN
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 IBIAS
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VSS
port 5 nsew
<< end >>
