magic
tech sky130A
magscale 1 2
timestamp 1769590285
<< pwell >>
rect -615 -471 615 471
<< mvnmos >>
rect -387 -213 -237 213
rect -179 -213 -29 213
rect 29 -213 179 213
rect 237 -213 387 213
<< mvndiff >>
rect -445 201 -387 213
rect -445 -201 -433 201
rect -399 -201 -387 201
rect -445 -213 -387 -201
rect -237 201 -179 213
rect -237 -201 -225 201
rect -191 -201 -179 201
rect -237 -213 -179 -201
rect -29 201 29 213
rect -29 -201 -17 201
rect 17 -201 29 201
rect -29 -213 29 -201
rect 179 201 237 213
rect 179 -201 191 201
rect 225 -201 237 201
rect 179 -213 237 -201
rect 387 201 445 213
rect 387 -201 399 201
rect 433 -201 445 201
rect 387 -213 445 -201
<< mvndiffc >>
rect -433 -201 -399 201
rect -225 -201 -191 201
rect -17 -201 17 201
rect 191 -201 225 201
rect 399 -201 433 201
<< mvpsubdiff >>
rect -579 423 579 435
rect -579 389 -471 423
rect 471 389 579 423
rect -579 377 579 389
rect -579 327 -521 377
rect -579 -327 -567 327
rect -533 -327 -521 327
rect 521 327 579 377
rect -579 -377 -521 -327
rect 521 -327 533 327
rect 567 -327 579 327
rect 521 -377 579 -327
rect -579 -389 579 -377
rect -579 -423 -471 -389
rect 471 -423 579 -389
rect -579 -435 579 -423
<< mvpsubdiffcont >>
rect -471 389 471 423
rect -567 -327 -533 327
rect 533 -327 567 327
rect -471 -423 471 -389
<< poly >>
rect -387 285 -237 301
rect -387 251 -371 285
rect -253 251 -237 285
rect -387 213 -237 251
rect -179 285 -29 301
rect -179 251 -163 285
rect -45 251 -29 285
rect -179 213 -29 251
rect 29 285 179 301
rect 29 251 45 285
rect 163 251 179 285
rect 29 213 179 251
rect 237 285 387 301
rect 237 251 253 285
rect 371 251 387 285
rect 237 213 387 251
rect -387 -251 -237 -213
rect -387 -285 -371 -251
rect -253 -285 -237 -251
rect -387 -301 -237 -285
rect -179 -251 -29 -213
rect -179 -285 -163 -251
rect -45 -285 -29 -251
rect -179 -301 -29 -285
rect 29 -251 179 -213
rect 29 -285 45 -251
rect 163 -285 179 -251
rect 29 -301 179 -285
rect 237 -251 387 -213
rect 237 -285 253 -251
rect 371 -285 387 -251
rect 237 -301 387 -285
<< polycont >>
rect -371 251 -253 285
rect -163 251 -45 285
rect 45 251 163 285
rect 253 251 371 285
rect -371 -285 -253 -251
rect -163 -285 -45 -251
rect 45 -285 163 -251
rect 253 -285 371 -251
<< locali >>
rect -567 389 -471 423
rect 471 389 567 423
rect -567 327 -533 389
rect 533 327 567 389
rect -387 251 -371 285
rect -253 251 -237 285
rect -179 251 -163 285
rect -45 251 -29 285
rect 29 251 45 285
rect 163 251 179 285
rect 237 251 253 285
rect 371 251 387 285
rect -433 201 -399 217
rect -433 -217 -399 -201
rect -225 201 -191 217
rect -225 -217 -191 -201
rect -17 201 17 217
rect -17 -217 17 -201
rect 191 201 225 217
rect 191 -217 225 -201
rect 399 201 433 217
rect 399 -217 433 -201
rect -387 -285 -371 -251
rect -253 -285 -237 -251
rect -179 -285 -163 -251
rect -45 -285 -29 -251
rect 29 -285 45 -251
rect 163 -285 179 -251
rect 237 -285 253 -251
rect 371 -285 387 -251
rect -567 -389 -533 -327
rect 533 -389 567 -327
rect -567 -423 -471 -389
rect 471 -423 567 -389
<< viali >>
rect -371 251 -253 285
rect -163 251 -45 285
rect 45 251 163 285
rect 253 251 371 285
rect -433 -201 -399 201
rect -225 -201 -191 201
rect -17 -201 17 201
rect 191 -201 225 201
rect 399 -201 433 201
rect -371 -285 -253 -251
rect -163 -285 -45 -251
rect 45 -285 163 -251
rect 253 -285 371 -251
<< metal1 >>
rect -383 285 -241 291
rect -383 251 -371 285
rect -253 251 -241 285
rect -383 245 -241 251
rect -175 285 -33 291
rect -175 251 -163 285
rect -45 251 -33 285
rect -175 245 -33 251
rect 33 285 175 291
rect 33 251 45 285
rect 163 251 175 285
rect 33 245 175 251
rect 241 285 383 291
rect 241 251 253 285
rect 371 251 383 285
rect 241 245 383 251
rect -439 201 -393 213
rect -439 -201 -433 201
rect -399 -201 -393 201
rect -439 -213 -393 -201
rect -231 201 -185 213
rect -231 -201 -225 201
rect -191 -201 -185 201
rect -231 -213 -185 -201
rect -23 201 23 213
rect -23 -201 -17 201
rect 17 -201 23 201
rect -23 -213 23 -201
rect 185 201 231 213
rect 185 -201 191 201
rect 225 -201 231 201
rect 185 -213 231 -201
rect 393 201 439 213
rect 393 -201 399 201
rect 433 -201 439 201
rect 393 -213 439 -201
rect -383 -251 -241 -245
rect -383 -285 -371 -251
rect -253 -285 -241 -251
rect -383 -291 -241 -285
rect -175 -251 -33 -245
rect -175 -285 -163 -251
rect -45 -285 -33 -251
rect -175 -291 -33 -285
rect 33 -251 175 -245
rect 33 -285 45 -251
rect 163 -285 175 -251
rect 33 -291 175 -285
rect 241 -251 383 -245
rect 241 -285 253 -251
rect 371 -285 383 -251
rect 241 -291 383 -285
<< properties >>
string FIXED_BBOX -550 -406 550 406
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.125 l 0.75 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
