magic
tech sky130A
magscale 1 2
timestamp 1770105080
<< pwell >>
rect -815 -1758 815 1758
<< mvnmos >>
rect -587 -1500 -337 1500
rect -279 -1500 -29 1500
rect 29 -1500 279 1500
rect 337 -1500 587 1500
<< mvndiff >>
rect -645 1488 -587 1500
rect -645 -1488 -633 1488
rect -599 -1488 -587 1488
rect -645 -1500 -587 -1488
rect -337 1488 -279 1500
rect -337 -1488 -325 1488
rect -291 -1488 -279 1488
rect -337 -1500 -279 -1488
rect -29 1488 29 1500
rect -29 -1488 -17 1488
rect 17 -1488 29 1488
rect -29 -1500 29 -1488
rect 279 1488 337 1500
rect 279 -1488 291 1488
rect 325 -1488 337 1488
rect 279 -1500 337 -1488
rect 587 1488 645 1500
rect 587 -1488 599 1488
rect 633 -1488 645 1488
rect 587 -1500 645 -1488
<< mvndiffc >>
rect -633 -1488 -599 1488
rect -325 -1488 -291 1488
rect -17 -1488 17 1488
rect 291 -1488 325 1488
rect 599 -1488 633 1488
<< mvpsubdiff >>
rect -779 1710 779 1722
rect -779 1676 -671 1710
rect 671 1676 779 1710
rect -779 1664 779 1676
rect -779 1614 -721 1664
rect -779 -1614 -767 1614
rect -733 -1614 -721 1614
rect 721 1614 779 1664
rect -779 -1664 -721 -1614
rect 721 -1614 733 1614
rect 767 -1614 779 1614
rect 721 -1664 779 -1614
rect -779 -1676 779 -1664
rect -779 -1710 -671 -1676
rect 671 -1710 779 -1676
rect -779 -1722 779 -1710
<< mvpsubdiffcont >>
rect -671 1676 671 1710
rect -767 -1614 -733 1614
rect 733 -1614 767 1614
rect -671 -1710 671 -1676
<< poly >>
rect -587 1572 -337 1588
rect -587 1538 -571 1572
rect -353 1538 -337 1572
rect -587 1500 -337 1538
rect -279 1572 -29 1588
rect -279 1538 -263 1572
rect -45 1538 -29 1572
rect -279 1500 -29 1538
rect 29 1572 279 1588
rect 29 1538 45 1572
rect 263 1538 279 1572
rect 29 1500 279 1538
rect 337 1572 587 1588
rect 337 1538 353 1572
rect 571 1538 587 1572
rect 337 1500 587 1538
rect -587 -1538 -337 -1500
rect -587 -1572 -571 -1538
rect -353 -1572 -337 -1538
rect -587 -1588 -337 -1572
rect -279 -1538 -29 -1500
rect -279 -1572 -263 -1538
rect -45 -1572 -29 -1538
rect -279 -1588 -29 -1572
rect 29 -1538 279 -1500
rect 29 -1572 45 -1538
rect 263 -1572 279 -1538
rect 29 -1588 279 -1572
rect 337 -1538 587 -1500
rect 337 -1572 353 -1538
rect 571 -1572 587 -1538
rect 337 -1588 587 -1572
<< polycont >>
rect -571 1538 -353 1572
rect -263 1538 -45 1572
rect 45 1538 263 1572
rect 353 1538 571 1572
rect -571 -1572 -353 -1538
rect -263 -1572 -45 -1538
rect 45 -1572 263 -1538
rect 353 -1572 571 -1538
<< locali >>
rect -767 1676 -671 1710
rect 671 1676 767 1710
rect -767 1614 -733 1676
rect 733 1614 767 1676
rect -587 1538 -571 1572
rect -353 1538 -337 1572
rect -279 1538 -263 1572
rect -45 1538 -29 1572
rect 29 1538 45 1572
rect 263 1538 279 1572
rect 337 1538 353 1572
rect 571 1538 587 1572
rect -633 1488 -599 1504
rect -633 -1504 -599 -1488
rect -325 1488 -291 1504
rect -325 -1504 -291 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 291 1488 325 1504
rect 291 -1504 325 -1488
rect 599 1488 633 1504
rect 599 -1504 633 -1488
rect -587 -1572 -571 -1538
rect -353 -1572 -337 -1538
rect -279 -1572 -263 -1538
rect -45 -1572 -29 -1538
rect 29 -1572 45 -1538
rect 263 -1572 279 -1538
rect 337 -1572 353 -1538
rect 571 -1572 587 -1538
rect -767 -1676 -733 -1614
rect 733 -1676 767 -1614
rect -767 -1710 -671 -1676
rect 671 -1710 767 -1676
<< viali >>
rect -571 1538 -353 1572
rect -263 1538 -45 1572
rect 45 1538 263 1572
rect 353 1538 571 1572
rect -633 -1488 -599 1488
rect -325 -1488 -291 1488
rect -17 -1488 17 1488
rect 291 -1488 325 1488
rect 599 -1488 633 1488
rect -571 -1572 -353 -1538
rect -263 -1572 -45 -1538
rect 45 -1572 263 -1538
rect 353 -1572 571 -1538
<< metal1 >>
rect -583 1572 -341 1578
rect -583 1538 -571 1572
rect -353 1538 -341 1572
rect -583 1532 -341 1538
rect -275 1572 -33 1578
rect -275 1538 -263 1572
rect -45 1538 -33 1572
rect -275 1532 -33 1538
rect 33 1572 275 1578
rect 33 1538 45 1572
rect 263 1538 275 1572
rect 33 1532 275 1538
rect 341 1572 583 1578
rect 341 1538 353 1572
rect 571 1538 583 1572
rect 341 1532 583 1538
rect -639 1488 -593 1500
rect -639 -1488 -633 1488
rect -599 -1488 -593 1488
rect -639 -1500 -593 -1488
rect -331 1488 -285 1500
rect -331 -1488 -325 1488
rect -291 -1488 -285 1488
rect -331 -1500 -285 -1488
rect -23 1488 23 1500
rect -23 -1488 -17 1488
rect 17 -1488 23 1488
rect -23 -1500 23 -1488
rect 285 1488 331 1500
rect 285 -1488 291 1488
rect 325 -1488 331 1488
rect 285 -1500 331 -1488
rect 593 1488 639 1500
rect 593 -1488 599 1488
rect 633 -1488 639 1488
rect 593 -1500 639 -1488
rect -583 -1538 -341 -1532
rect -583 -1572 -571 -1538
rect -353 -1572 -341 -1538
rect -583 -1578 -341 -1572
rect -275 -1538 -33 -1532
rect -275 -1572 -263 -1538
rect -45 -1572 -33 -1538
rect -275 -1578 -33 -1572
rect 33 -1538 275 -1532
rect 33 -1572 45 -1538
rect 263 -1572 275 -1538
rect 33 -1578 275 -1572
rect 341 -1538 583 -1532
rect 341 -1572 353 -1538
rect 571 -1572 583 -1538
rect 341 -1578 583 -1572
<< properties >>
string FIXED_BBOX -750 -1693 750 1693
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 15.0 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
