magic
tech sky130A
magscale 1 2
timestamp 1770035380
<< error_p >>
rect -2559 1098 2559 1102
rect -2559 -1030 -2529 1098
rect -2493 1032 2493 1036
rect -2493 -964 -2463 1032
rect 2463 -964 2493 1032
rect -2344 -1011 -2276 -1005
rect -2036 -1011 -1968 -1005
rect -1728 -1011 -1660 -1005
rect -1420 -1011 -1352 -1005
rect -1112 -1011 -1044 -1005
rect -804 -1011 -736 -1005
rect -496 -1011 -428 -1005
rect -188 -1011 -120 -1005
rect 428 -1011 496 -1005
rect 736 -1011 804 -1005
rect 1044 -1011 1112 -1005
rect 1352 -1011 1420 -1005
rect 1660 -1011 1728 -1005
rect 1968 -1011 2036 -1005
rect 2276 -1011 2344 -1005
rect -2344 -1045 -2332 -1011
rect -2036 -1045 -2024 -1011
rect -1728 -1045 -1716 -1011
rect -1420 -1045 -1408 -1011
rect -1112 -1045 -1100 -1011
rect -804 -1045 -792 -1011
rect -496 -1045 -484 -1011
rect -188 -1045 -176 -1011
rect 428 -1045 440 -1011
rect 736 -1045 748 -1011
rect 1044 -1045 1056 -1011
rect 1352 -1045 1364 -1011
rect 1660 -1045 1672 -1011
rect 1968 -1045 1980 -1011
rect 2276 -1045 2288 -1011
rect 2529 -1030 2559 1098
rect -2344 -1051 -2276 -1045
rect -2036 -1051 -1968 -1045
rect -1728 -1051 -1660 -1045
rect -1420 -1051 -1352 -1045
rect -1112 -1051 -1044 -1045
rect -804 -1051 -736 -1045
rect -496 -1051 -428 -1045
rect -188 -1051 -120 -1045
rect 428 -1051 496 -1045
rect 736 -1051 804 -1045
rect 1044 -1051 1112 -1045
rect 1352 -1051 1420 -1045
rect 1660 -1051 1728 -1045
rect 1968 -1051 2036 -1045
rect 2276 -1051 2344 -1045
<< nwell >>
rect -2529 -1064 2529 1098
<< mvpmos >>
rect -2435 -964 -2185 1036
rect -2127 -964 -1877 1036
rect -1819 -964 -1569 1036
rect -1511 -964 -1261 1036
rect -1203 -964 -953 1036
rect -895 -964 -645 1036
rect -587 -964 -337 1036
rect -279 -964 -29 1036
rect 29 -964 279 1036
rect 337 -964 587 1036
rect 645 -964 895 1036
rect 953 -964 1203 1036
rect 1261 -964 1511 1036
rect 1569 -964 1819 1036
rect 1877 -964 2127 1036
rect 2185 -964 2435 1036
<< mvpdiff >>
rect -2493 1024 -2435 1036
rect -2493 -952 -2481 1024
rect -2447 -952 -2435 1024
rect -2493 -964 -2435 -952
rect -2185 1024 -2127 1036
rect -2185 -952 -2173 1024
rect -2139 -952 -2127 1024
rect -2185 -964 -2127 -952
rect -1877 1024 -1819 1036
rect -1877 -952 -1865 1024
rect -1831 -952 -1819 1024
rect -1877 -964 -1819 -952
rect -1569 1024 -1511 1036
rect -1569 -952 -1557 1024
rect -1523 -952 -1511 1024
rect -1569 -964 -1511 -952
rect -1261 1024 -1203 1036
rect -1261 -952 -1249 1024
rect -1215 -952 -1203 1024
rect -1261 -964 -1203 -952
rect -953 1024 -895 1036
rect -953 -952 -941 1024
rect -907 -952 -895 1024
rect -953 -964 -895 -952
rect -645 1024 -587 1036
rect -645 -952 -633 1024
rect -599 -952 -587 1024
rect -645 -964 -587 -952
rect -337 1024 -279 1036
rect -337 -952 -325 1024
rect -291 -952 -279 1024
rect -337 -964 -279 -952
rect -29 1024 29 1036
rect -29 -952 -17 1024
rect 17 -952 29 1024
rect -29 -964 29 -952
rect 279 1024 337 1036
rect 279 -952 291 1024
rect 325 -952 337 1024
rect 279 -964 337 -952
rect 587 1024 645 1036
rect 587 -952 599 1024
rect 633 -952 645 1024
rect 587 -964 645 -952
rect 895 1024 953 1036
rect 895 -952 907 1024
rect 941 -952 953 1024
rect 895 -964 953 -952
rect 1203 1024 1261 1036
rect 1203 -952 1215 1024
rect 1249 -952 1261 1024
rect 1203 -964 1261 -952
rect 1511 1024 1569 1036
rect 1511 -952 1523 1024
rect 1557 -952 1569 1024
rect 1511 -964 1569 -952
rect 1819 1024 1877 1036
rect 1819 -952 1831 1024
rect 1865 -952 1877 1024
rect 1819 -964 1877 -952
rect 2127 1024 2185 1036
rect 2127 -952 2139 1024
rect 2173 -952 2185 1024
rect 2127 -964 2185 -952
rect 2435 1024 2493 1036
rect 2435 -952 2447 1024
rect 2481 -952 2493 1024
rect 2435 -964 2493 -952
<< mvpdiffc >>
rect -2481 -952 -2447 1024
rect -2173 -952 -2139 1024
rect -1865 -952 -1831 1024
rect -1557 -952 -1523 1024
rect -1249 -952 -1215 1024
rect -941 -952 -907 1024
rect -633 -952 -599 1024
rect -325 -952 -291 1024
rect -17 -952 17 1024
rect 291 -952 325 1024
rect 599 -952 633 1024
rect 907 -952 941 1024
rect 1215 -952 1249 1024
rect 1523 -952 1557 1024
rect 1831 -952 1865 1024
rect 2139 -952 2173 1024
rect 2447 -952 2481 1024
<< poly >>
rect -2435 1036 -2185 1062
rect -2127 1036 -1877 1062
rect -1819 1036 -1569 1062
rect -1511 1036 -1261 1062
rect -1203 1036 -953 1062
rect -895 1036 -645 1062
rect -587 1036 -337 1062
rect -279 1036 -29 1062
rect 29 1036 279 1062
rect 337 1036 587 1062
rect 645 1036 895 1062
rect 953 1036 1203 1062
rect 1261 1036 1511 1062
rect 1569 1036 1819 1062
rect 1877 1036 2127 1062
rect 2185 1036 2435 1062
rect -2435 -1011 -2185 -964
rect -2435 -1028 -2332 -1011
rect -2348 -1045 -2332 -1028
rect -2288 -1028 -2185 -1011
rect -2127 -1011 -1877 -964
rect -2127 -1028 -2024 -1011
rect -2288 -1045 -2272 -1028
rect -2348 -1061 -2272 -1045
rect -2040 -1045 -2024 -1028
rect -1980 -1028 -1877 -1011
rect -1819 -1011 -1569 -964
rect -1819 -1028 -1716 -1011
rect -1980 -1045 -1964 -1028
rect -2040 -1061 -1964 -1045
rect -1732 -1045 -1716 -1028
rect -1672 -1028 -1569 -1011
rect -1511 -1011 -1261 -964
rect -1511 -1028 -1408 -1011
rect -1672 -1045 -1656 -1028
rect -1732 -1061 -1656 -1045
rect -1424 -1045 -1408 -1028
rect -1364 -1028 -1261 -1011
rect -1203 -1011 -953 -964
rect -1203 -1028 -1100 -1011
rect -1364 -1045 -1348 -1028
rect -1424 -1061 -1348 -1045
rect -1116 -1045 -1100 -1028
rect -1056 -1028 -953 -1011
rect -895 -1011 -645 -964
rect -895 -1028 -792 -1011
rect -1056 -1045 -1040 -1028
rect -1116 -1061 -1040 -1045
rect -808 -1045 -792 -1028
rect -748 -1028 -645 -1011
rect -587 -1011 -337 -964
rect -587 -1028 -484 -1011
rect -748 -1045 -732 -1028
rect -808 -1061 -732 -1045
rect -500 -1045 -484 -1028
rect -440 -1028 -337 -1011
rect -279 -1011 -29 -964
rect -279 -1028 -176 -1011
rect -440 -1045 -424 -1028
rect -500 -1061 -424 -1045
rect -192 -1045 -176 -1028
rect -132 -1028 -29 -1011
rect 29 -1011 279 -964
rect 29 -1028 132 -1011
rect -132 -1045 -116 -1028
rect -192 -1061 -116 -1045
rect 116 -1045 132 -1028
rect 176 -1028 279 -1011
rect 337 -1011 587 -964
rect 337 -1028 440 -1011
rect 176 -1045 192 -1028
rect 116 -1061 192 -1045
rect 424 -1045 440 -1028
rect 484 -1028 587 -1011
rect 645 -1011 895 -964
rect 645 -1028 748 -1011
rect 484 -1045 500 -1028
rect 424 -1061 500 -1045
rect 732 -1045 748 -1028
rect 792 -1028 895 -1011
rect 953 -1011 1203 -964
rect 953 -1028 1056 -1011
rect 792 -1045 808 -1028
rect 732 -1061 808 -1045
rect 1040 -1045 1056 -1028
rect 1100 -1028 1203 -1011
rect 1261 -1011 1511 -964
rect 1261 -1028 1364 -1011
rect 1100 -1045 1116 -1028
rect 1040 -1061 1116 -1045
rect 1348 -1045 1364 -1028
rect 1408 -1028 1511 -1011
rect 1569 -1011 1819 -964
rect 1569 -1028 1672 -1011
rect 1408 -1045 1424 -1028
rect 1348 -1061 1424 -1045
rect 1656 -1045 1672 -1028
rect 1716 -1028 1819 -1011
rect 1877 -1011 2127 -964
rect 1877 -1028 1980 -1011
rect 1716 -1045 1732 -1028
rect 1656 -1061 1732 -1045
rect 1964 -1045 1980 -1028
rect 2024 -1028 2127 -1011
rect 2185 -1011 2435 -964
rect 2185 -1028 2288 -1011
rect 2024 -1045 2040 -1028
rect 1964 -1061 2040 -1045
rect 2272 -1045 2288 -1028
rect 2332 -1028 2435 -1011
rect 2332 -1045 2348 -1028
rect 2272 -1061 2348 -1045
<< polycont >>
rect -2332 -1045 -2288 -1011
rect -2024 -1045 -1980 -1011
rect -1716 -1045 -1672 -1011
rect -1408 -1045 -1364 -1011
rect -1100 -1045 -1056 -1011
rect -792 -1045 -748 -1011
rect -484 -1045 -440 -1011
rect -176 -1045 -132 -1011
rect 132 -1045 176 -1011
rect 440 -1045 484 -1011
rect 748 -1045 792 -1011
rect 1056 -1045 1100 -1011
rect 1364 -1045 1408 -1011
rect 1672 -1045 1716 -1011
rect 1980 -1045 2024 -1011
rect 2288 -1045 2332 -1011
<< locali >>
rect -2481 1024 -2447 1040
rect -2481 -968 -2447 -952
rect -2173 1024 -2139 1040
rect -2173 -968 -2139 -952
rect -1865 1024 -1831 1040
rect -1865 -968 -1831 -952
rect -1557 1024 -1523 1040
rect -1557 -968 -1523 -952
rect -1249 1024 -1215 1040
rect -1249 -968 -1215 -952
rect -941 1024 -907 1040
rect -941 -968 -907 -952
rect -633 1024 -599 1040
rect -633 -968 -599 -952
rect -325 1024 -291 1040
rect -325 -968 -291 -952
rect -17 1024 17 1040
rect -17 -968 17 -952
rect 291 1024 325 1040
rect 291 -968 325 -952
rect 599 1024 633 1040
rect 599 -968 633 -952
rect 907 1024 941 1040
rect 907 -968 941 -952
rect 1215 1024 1249 1040
rect 1215 -968 1249 -952
rect 1523 1024 1557 1040
rect 1523 -968 1557 -952
rect 1831 1024 1865 1040
rect 1831 -968 1865 -952
rect 2139 1024 2173 1040
rect 2139 -968 2173 -952
rect 2447 1024 2481 1040
rect 2447 -968 2481 -952
rect -2348 -1045 -2332 -1011
rect -2288 -1045 -2272 -1011
rect -2040 -1045 -2024 -1011
rect -1980 -1045 -1964 -1011
rect -1732 -1045 -1716 -1011
rect -1672 -1045 -1656 -1011
rect -1424 -1045 -1408 -1011
rect -1364 -1045 -1348 -1011
rect -1116 -1045 -1100 -1011
rect -1056 -1045 -1040 -1011
rect -808 -1045 -792 -1011
rect -748 -1045 -732 -1011
rect -500 -1045 -484 -1011
rect -440 -1045 -424 -1011
rect -192 -1045 -176 -1011
rect -132 -1045 -116 -1011
rect 116 -1045 132 -1011
rect 176 -1045 192 -1011
rect 424 -1045 440 -1011
rect 484 -1045 500 -1011
rect 732 -1045 748 -1011
rect 792 -1045 808 -1011
rect 1040 -1045 1056 -1011
rect 1100 -1045 1116 -1011
rect 1348 -1045 1364 -1011
rect 1408 -1045 1424 -1011
rect 1656 -1045 1672 -1011
rect 1716 -1045 1732 -1011
rect 1964 -1045 1980 -1011
rect 2024 -1045 2040 -1011
rect 2272 -1045 2288 -1011
rect 2332 -1045 2348 -1011
<< viali >>
rect -2481 -952 -2447 1024
rect -2173 -952 -2139 1024
rect -1865 -952 -1831 1024
rect -1557 -952 -1523 1024
rect -1249 -952 -1215 1024
rect -941 -952 -907 1024
rect -633 -952 -599 1024
rect -325 -952 -291 1024
rect -17 -952 17 1024
rect 291 -952 325 1024
rect 599 -952 633 1024
rect 907 -952 941 1024
rect 1215 -952 1249 1024
rect 1523 -952 1557 1024
rect 1831 -952 1865 1024
rect 2139 -952 2173 1024
rect 2447 -952 2481 1024
rect -2332 -1045 -2288 -1011
rect -2024 -1045 -1980 -1011
rect -1716 -1045 -1672 -1011
rect -1408 -1045 -1364 -1011
rect -1100 -1045 -1056 -1011
rect -792 -1045 -748 -1011
rect -484 -1045 -440 -1011
rect -176 -1045 -132 -1011
rect 132 -1045 176 -1011
rect 440 -1045 484 -1011
rect 748 -1045 792 -1011
rect 1056 -1045 1100 -1011
rect 1364 -1045 1408 -1011
rect 1672 -1045 1716 -1011
rect 1980 -1045 2024 -1011
rect 2288 -1045 2332 -1011
<< metal1 >>
rect -2487 1024 -2441 1036
rect -2487 -952 -2481 1024
rect -2447 -952 -2441 1024
rect -2487 -964 -2441 -952
rect -2179 1024 -2133 1036
rect -2179 -952 -2173 1024
rect -2139 -952 -2133 1024
rect -2179 -964 -2133 -952
rect -1871 1024 -1825 1036
rect -1871 -952 -1865 1024
rect -1831 -952 -1825 1024
rect -1871 -964 -1825 -952
rect -1563 1024 -1517 1036
rect -1563 -952 -1557 1024
rect -1523 -952 -1517 1024
rect -1563 -964 -1517 -952
rect -1255 1024 -1209 1036
rect -1255 -952 -1249 1024
rect -1215 -952 -1209 1024
rect -1255 -964 -1209 -952
rect -947 1024 -901 1036
rect -947 -952 -941 1024
rect -907 -952 -901 1024
rect -947 -964 -901 -952
rect -639 1024 -593 1036
rect -639 -952 -633 1024
rect -599 -952 -593 1024
rect -639 -964 -593 -952
rect -331 1024 -285 1036
rect -331 -952 -325 1024
rect -291 -952 -285 1024
rect -331 -964 -285 -952
rect -23 1024 23 1036
rect -23 -952 -17 1024
rect 17 200 23 1024
rect 285 1024 331 1036
rect 17 0 200 200
rect 17 -200 23 0
rect 17 -400 200 -200
rect 17 -600 23 -400
rect 17 -800 200 -600
rect 17 -952 23 -800
rect -23 -964 23 -952
rect 285 -952 291 1024
rect 325 -952 331 1024
rect 285 -964 331 -952
rect 593 1024 639 1036
rect 593 -952 599 1024
rect 633 -952 639 1024
rect 593 -964 639 -952
rect 901 1024 947 1036
rect 901 -952 907 1024
rect 941 -952 947 1024
rect 901 -964 947 -952
rect 1209 1024 1255 1036
rect 1209 -952 1215 1024
rect 1249 -952 1255 1024
rect 1209 -964 1255 -952
rect 1517 1024 1563 1036
rect 1517 -952 1523 1024
rect 1557 -952 1563 1024
rect 1517 -964 1563 -952
rect 1825 1024 1871 1036
rect 1825 -952 1831 1024
rect 1865 -952 1871 1024
rect 1825 -964 1871 -952
rect 2133 1024 2179 1036
rect 2133 -952 2139 1024
rect 2173 -952 2179 1024
rect 2133 -964 2179 -952
rect 2441 1024 2487 1036
rect 2441 -952 2447 1024
rect 2481 -952 2487 1024
rect 2441 -964 2487 -952
rect -2344 -1011 -2276 -1005
rect -2344 -1045 -2332 -1011
rect -2288 -1045 -2276 -1011
rect -2344 -1051 -2276 -1045
rect -2036 -1011 -1968 -1005
rect -2036 -1045 -2024 -1011
rect -1980 -1045 -1968 -1011
rect -2036 -1051 -1968 -1045
rect -1728 -1011 -1660 -1005
rect -1728 -1045 -1716 -1011
rect -1672 -1045 -1660 -1011
rect -1728 -1051 -1660 -1045
rect -1420 -1011 -1352 -1005
rect -1420 -1045 -1408 -1011
rect -1364 -1045 -1352 -1011
rect -1420 -1051 -1352 -1045
rect -1112 -1011 -1044 -1005
rect -1112 -1045 -1100 -1011
rect -1056 -1045 -1044 -1011
rect -1112 -1051 -1044 -1045
rect -804 -1011 -736 -1005
rect -804 -1045 -792 -1011
rect -748 -1045 -736 -1011
rect -804 -1051 -736 -1045
rect -496 -1011 -428 -1005
rect -496 -1045 -484 -1011
rect -440 -1045 -428 -1011
rect -496 -1051 -428 -1045
rect -188 -1011 -120 -1005
rect -188 -1045 -176 -1011
rect -132 -1045 -120 -1011
rect -188 -1051 -120 -1045
rect 0 -1011 200 -1000
rect 0 -1045 132 -1011
rect 176 -1045 200 -1011
rect 0 -1200 200 -1045
rect 428 -1011 496 -1005
rect 428 -1045 440 -1011
rect 484 -1045 496 -1011
rect 428 -1051 496 -1045
rect 736 -1011 804 -1005
rect 736 -1045 748 -1011
rect 792 -1045 804 -1011
rect 736 -1051 804 -1045
rect 1044 -1011 1112 -1005
rect 1044 -1045 1056 -1011
rect 1100 -1045 1112 -1011
rect 1044 -1051 1112 -1045
rect 1352 -1011 1420 -1005
rect 1352 -1045 1364 -1011
rect 1408 -1045 1420 -1011
rect 1352 -1051 1420 -1045
rect 1660 -1011 1728 -1005
rect 1660 -1045 1672 -1011
rect 1716 -1045 1728 -1011
rect 1660 -1051 1728 -1045
rect 1968 -1011 2036 -1005
rect 1968 -1045 1980 -1011
rect 2024 -1045 2036 -1011
rect 1968 -1051 2036 -1045
rect 2276 -1011 2344 -1005
rect 2276 -1045 2288 -1011
rect 2332 -1045 2344 -1011
rect 2276 -1051 2344 -1045
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
rect 0 -8800 200 -8600
rect 0 -9200 200 -9000
rect 0 -9600 200 -9400
rect 0 -10000 200 -9800
rect 0 -10400 200 -10200
rect 0 -10800 200 -10600
rect 0 -11200 200 -11000
rect 0 -11600 200 -11400
rect 0 -12000 200 -11800
rect 0 -12400 200 -12200
rect 0 -12800 200 -12600
rect 0 -13200 200 -13000
rect 0 -13600 200 -13400
rect 0 -14000 200 -13800
rect 0 -14400 200 -14200
rect 0 -14800 200 -14600
rect 0 -15200 200 -15000
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X0
timestamp 0
transform 1 0 -2271 0 1 -13998
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X1
timestamp 0
transform 1 0 -1600 0 1 -14093
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X2
timestamp 0
transform 1 0 -929 0 1 -14188
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X3
timestamp 0
transform 1 0 -258 0 1 -14283
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X4
timestamp 0
transform 1 0 413 0 1 -14378
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X5
timestamp 0
transform 1 0 1084 0 1 -14473
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X6
timestamp 0
transform 1 0 1755 0 1 -14568
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X7
timestamp 0
transform 1 0 2426 0 1 -14663
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_XJB3AQ  X8
timestamp 0
transform 1 0 3097 0 1 -14758
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X9
timestamp 0
transform 1 0 3768 0 1 -14853
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X10
timestamp 0
transform 1 0 4439 0 1 -14948
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_UUE6JB  X11
timestamp 0
transform 1 0 5110 0 1 -15043
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X12
timestamp 0
transform 1 0 5781 0 1 -15138
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X13
timestamp 0
transform 1 0 6452 0 1 -15233
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X14
timestamp 0
transform 1 0 7123 0 1 -15328
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_Y5UTF8  X15
timestamp 0
transform 1 0 7794 0 1 -15423
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 a_2127_n964#
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 a_n2493_n964#
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 a_n2127_n1028#
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 {}
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 a_587_n964#
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 a_1569_n1028#
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 a_1203_n964#
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 a_n1877_n964#
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 a_953_n1028#
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 a_337_n1028#
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 a_n279_n1028#
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 a_n895_n1028#
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 a_n1819_n1028#
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 a_n337_n964#
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 a_n1203_n1028#
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 a_n953_n964#
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 a_2185_n1028#
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 {}
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 a_29_n1028#
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 w_n2529_n1064#
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 256 0 0 0 a_2435_n964#
port 21 nsew
flabel metal1 0 -8800 200 -8600 0 FreeSans 256 0 0 0 a_n2185_n964#
port 22 nsew
flabel metal1 0 -9200 200 -9000 0 FreeSans 256 0 0 0 a_n2435_n1028#
port 23 nsew
flabel metal1 0 -9600 200 -9400 0 FreeSans 256 0 0 0 a_279_n964#
port 24 nsew
flabel metal1 0 -10000 200 -9800 0 FreeSans 256 0 0 0 {}
port 25 nsew
flabel metal1 0 -10400 200 -10200 0 FreeSans 256 0 0 0 a_1877_n1028#
port 26 nsew
flabel metal1 0 -10800 200 -10600 0 FreeSans 256 0 0 0 a_895_n964#
port 27 nsew
flabel metal1 0 -11200 200 -11000 0 FreeSans 256 0 0 0 a_1261_n1028#
port 28 nsew
flabel metal1 0 -11600 200 -11400 0 FreeSans 256 0 0 0 a_n1261_n964#
port 29 nsew
flabel metal1 0 -12000 200 -11800 0 FreeSans 256 0 0 0 a_1511_n964#
port 30 nsew
flabel metal1 0 -12400 200 -12200 0 FreeSans 256 0 0 0 a_n1569_n964#
port 31 nsew
flabel metal1 0 -12800 200 -12600 0 FreeSans 256 0 0 0 {}
port 32 nsew
flabel metal1 0 -13200 200 -13000 0 FreeSans 256 0 0 0 a_1819_n964#
port 33 nsew
flabel metal1 0 -13600 200 -13400 0 FreeSans 256 0 0 0 a_645_n1028#
port 34 nsew
flabel metal1 0 -14000 200 -13800 0 FreeSans 256 0 0 0 a_n587_n1028#
port 35 nsew
flabel metal1 0 -14400 200 -14200 0 FreeSans 256 0 0 0 a_n645_n964#
port 36 nsew
flabel metal1 0 -14800 200 -14600 0 FreeSans 256 0 0 0 a_n1511_n1028#
port 37 nsew
flabel metal1 0 -15200 200 -15000 0 FreeSans 256 0 0 0 a_n29_n964#
port 38 nsew
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 1.25 m 1 nf 16 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
