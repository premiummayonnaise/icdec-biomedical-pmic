magic
tech sky130A
magscale 1 2
timestamp 1768759254
<< error_p >>
rect -891 -309 -861 309
rect -825 -243 -795 243
rect 795 -243 825 243
rect 861 -309 891 309
<< nwell >>
rect -861 -343 861 343
<< mvpmos >>
rect -767 -243 -517 243
rect -339 -243 -89 243
rect 89 -243 339 243
rect 517 -243 767 243
<< mvpdiff >>
rect -825 231 -767 243
rect -825 -231 -813 231
rect -779 -231 -767 231
rect -825 -243 -767 -231
rect -517 231 -459 243
rect -517 -231 -505 231
rect -471 -231 -459 231
rect -517 -243 -459 -231
rect -397 231 -339 243
rect -397 -231 -385 231
rect -351 -231 -339 231
rect -397 -243 -339 -231
rect -89 231 -31 243
rect -89 -231 -77 231
rect -43 -231 -31 231
rect -89 -243 -31 -231
rect 31 231 89 243
rect 31 -231 43 231
rect 77 -231 89 231
rect 31 -243 89 -231
rect 339 231 397 243
rect 339 -231 351 231
rect 385 -231 397 231
rect 339 -243 397 -231
rect 459 231 517 243
rect 459 -231 471 231
rect 505 -231 517 231
rect 459 -243 517 -231
rect 767 231 825 243
rect 767 -231 779 231
rect 813 -231 825 231
rect 767 -243 825 -231
<< mvpdiffc >>
rect -813 -231 -779 231
rect -505 -231 -471 231
rect -385 -231 -351 231
rect -77 -231 -43 231
rect 43 -231 77 231
rect 351 -231 385 231
rect 471 -231 505 231
rect 779 -231 813 231
<< poly >>
rect -767 324 -517 340
rect -767 290 -751 324
rect -533 290 -517 324
rect -767 243 -517 290
rect -339 324 -89 340
rect -339 290 -323 324
rect -105 290 -89 324
rect -339 243 -89 290
rect 89 324 339 340
rect 89 290 105 324
rect 323 290 339 324
rect 89 243 339 290
rect 517 324 767 340
rect 517 290 533 324
rect 751 290 767 324
rect 517 243 767 290
rect -767 -290 -517 -243
rect -767 -324 -751 -290
rect -533 -324 -517 -290
rect -767 -340 -517 -324
rect -339 -290 -89 -243
rect -339 -324 -323 -290
rect -105 -324 -89 -290
rect -339 -340 -89 -324
rect 89 -290 339 -243
rect 89 -324 105 -290
rect 323 -324 339 -290
rect 89 -340 339 -324
rect 517 -290 767 -243
rect 517 -324 533 -290
rect 751 -324 767 -290
rect 517 -340 767 -324
<< polycont >>
rect -751 290 -533 324
rect -323 290 -105 324
rect 105 290 323 324
rect 533 290 751 324
rect -751 -324 -533 -290
rect -323 -324 -105 -290
rect 105 -324 323 -290
rect 533 -324 751 -290
<< locali >>
rect -767 290 -751 324
rect -533 290 -517 324
rect -339 290 -323 324
rect -105 290 -89 324
rect 89 290 105 324
rect 323 290 339 324
rect 517 290 533 324
rect 751 290 767 324
rect -813 231 -779 247
rect -813 -247 -779 -231
rect -505 231 -471 247
rect -505 -247 -471 -231
rect -385 231 -351 247
rect -385 -247 -351 -231
rect -77 231 -43 247
rect -77 -247 -43 -231
rect 43 231 77 247
rect 43 -247 77 -231
rect 351 231 385 247
rect 351 -247 385 -231
rect 471 231 505 247
rect 471 -247 505 -231
rect 779 231 813 247
rect 779 -247 813 -231
rect -767 -324 -751 -290
rect -533 -324 -517 -290
rect -339 -324 -323 -290
rect -105 -324 -89 -290
rect 89 -324 105 -290
rect 323 -324 339 -290
rect 517 -324 533 -290
rect 751 -324 767 -290
<< viali >>
rect -751 290 -533 324
rect -323 290 -105 324
rect 105 290 323 324
rect 533 290 751 324
rect -813 -231 -779 231
rect -505 -231 -471 231
rect -385 -231 -351 231
rect -77 -231 -43 231
rect 43 -231 77 231
rect 351 -231 385 231
rect 471 -231 505 231
rect 779 -231 813 231
rect -751 -324 -533 -290
rect -323 -324 -105 -290
rect 105 -324 323 -290
rect 533 -324 751 -290
<< metal1 >>
rect -763 324 -521 330
rect -763 290 -751 324
rect -533 290 -521 324
rect -763 284 -521 290
rect -335 324 -93 330
rect -335 290 -323 324
rect -105 290 -93 324
rect -335 284 -93 290
rect 93 324 335 330
rect 93 290 105 324
rect 323 290 335 324
rect 93 284 335 290
rect 521 324 763 330
rect 521 290 533 324
rect 751 290 763 324
rect 521 284 763 290
rect -819 231 -773 243
rect -819 -231 -813 231
rect -779 -231 -773 231
rect -819 -243 -773 -231
rect -511 231 -465 243
rect -511 -231 -505 231
rect -471 -231 -465 231
rect -511 -243 -465 -231
rect -391 231 -345 243
rect -391 -231 -385 231
rect -351 -231 -345 231
rect -391 -243 -345 -231
rect -83 231 -37 243
rect -83 -231 -77 231
rect -43 -231 -37 231
rect -83 -243 -37 -231
rect 37 231 83 243
rect 37 -231 43 231
rect 77 -231 83 231
rect 37 -243 83 -231
rect 345 231 391 243
rect 345 -231 351 231
rect 385 -231 391 231
rect 345 -243 391 -231
rect 465 231 511 243
rect 465 -231 471 231
rect 505 -231 511 231
rect 465 -243 511 -231
rect 773 231 819 243
rect 773 -231 779 231
rect 813 -231 819 231
rect 773 -243 819 -231
rect -763 -290 -521 -284
rect -763 -324 -751 -290
rect -533 -324 -521 -290
rect -763 -330 -521 -324
rect -335 -290 -93 -284
rect -335 -324 -323 -290
rect -105 -324 -93 -290
rect -335 -330 -93 -324
rect 93 -290 335 -284
rect 93 -324 105 -290
rect 323 -324 335 -290
rect 93 -330 335 -324
rect 521 -290 763 -284
rect 521 -324 533 -290
rect 751 -324 763 -290
rect 521 -330 763 -324
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.425 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
