magic
tech sky130A
magscale 1 2
timestamp 1770003475
<< pwell >>
rect 2100 -900 8100 1100
<< psubdiff >>
rect 2100 1080 8100 1100
rect 2100 1020 2220 1080
rect 7980 1020 8100 1080
rect 2100 1000 8100 1020
rect 2100 980 2200 1000
rect 2100 -780 2120 980
rect 2180 -780 2200 980
rect 2100 -800 2200 -780
rect 8000 980 8100 1000
rect 8000 -780 8020 980
rect 8080 -780 8100 980
rect 8000 -800 8100 -780
rect 2100 -820 8100 -800
rect 2100 -880 2220 -820
rect 7980 -880 8100 -820
rect 2100 -900 8100 -880
<< psubdiffcont >>
rect 2220 1020 7980 1080
rect 2120 -780 2180 980
rect 8020 -780 8080 980
rect 2220 -880 7980 -820
<< locali >>
rect 2100 1080 8100 1100
rect 2100 1020 2220 1080
rect 7980 1020 8100 1080
rect 2100 1000 8100 1020
rect 2100 980 2200 1000
rect 2100 -780 2120 980
rect 2180 -780 2200 980
rect 8000 980 8100 1000
rect 2340 180 2620 880
rect 2340 120 2440 180
rect 2500 120 2620 180
rect 2340 80 2620 120
rect 2340 20 2440 80
rect 2500 20 2620 80
rect 2340 -20 2620 20
rect 2340 -80 2440 -20
rect 2500 -80 2620 -20
rect 2340 -700 2620 -80
rect 2100 -800 2200 -780
rect 2880 -800 3000 800
rect 3500 -800 3620 800
rect 4120 -800 4240 800
rect 4720 -800 4840 800
rect 5340 -800 5460 800
rect 5960 -800 6080 800
rect 6580 -800 6700 800
rect 7200 -800 7320 800
rect 7580 180 7860 880
rect 7580 120 7680 180
rect 7740 120 7860 180
rect 7580 80 7860 120
rect 7580 20 7680 80
rect 7740 20 7860 80
rect 7580 -20 7860 20
rect 7580 -80 7680 -20
rect 7740 -80 7860 -20
rect 7580 -700 7860 -80
rect 8000 -780 8020 980
rect 8080 -780 8100 980
rect 8000 -800 8100 -780
rect 2100 -820 8100 -800
rect 2100 -880 2120 -820
rect 2180 -880 2220 -820
rect 7980 -880 8100 -820
rect 2100 -900 8100 -880
<< viali >>
rect 2440 120 2500 180
rect 2440 20 2500 80
rect 2440 -80 2500 -20
rect 7680 120 7740 180
rect 7680 20 7740 80
rect 7680 -80 7740 -20
rect 2120 -880 2180 -820
<< metal1 >>
rect 2660 860 7540 940
rect 1800 180 2100 200
rect 1800 120 1820 180
rect 1880 120 1920 180
rect 1980 120 2020 180
rect 2080 120 2100 180
rect 1800 80 2100 120
rect 1800 20 1820 80
rect 1880 20 1920 80
rect 1980 20 2020 80
rect 2080 20 2100 80
rect 1800 -20 2100 20
rect 1800 -80 1820 -20
rect 1880 -80 1920 -20
rect 1980 -80 2020 -20
rect 2080 -80 2100 -20
rect 1800 -100 2100 -80
rect 2420 180 2520 200
rect 2420 120 2440 180
rect 2500 120 2520 180
rect 2420 80 2520 120
rect 2420 20 2440 80
rect 2500 20 2520 80
rect 2420 -20 2520 20
rect 2420 -80 2440 -20
rect 2500 -80 2520 -20
rect 2420 -100 2520 -80
rect 3180 -320 3320 860
rect 3820 180 3920 200
rect 3820 120 3840 180
rect 3900 120 3920 180
rect 3820 80 3920 120
rect 3820 20 3840 80
rect 3900 20 3920 80
rect 3820 -20 3920 20
rect 3820 -80 3840 -20
rect 3900 -80 3920 -20
rect 3820 -100 3920 -80
rect 3180 -380 3220 -320
rect 3280 -380 3320 -320
rect 3180 -420 3320 -380
rect 3180 -480 3220 -420
rect 3280 -480 3320 -420
rect 3180 -520 3320 -480
rect 3180 -580 3220 -520
rect 3280 -580 3320 -520
rect 3180 -700 3320 -580
rect 4420 -320 4560 860
rect 5060 180 5160 200
rect 5060 120 5080 180
rect 5140 120 5160 180
rect 5060 80 5160 120
rect 5060 20 5080 80
rect 5140 20 5160 80
rect 5060 -20 5160 20
rect 5060 -80 5080 -20
rect 5140 -80 5160 -20
rect 5060 -100 5160 -80
rect 4420 -380 4460 -320
rect 4520 -380 4560 -320
rect 4420 -420 4560 -380
rect 4420 -480 4460 -420
rect 4520 -480 4560 -420
rect 4420 -520 4560 -480
rect 4420 -580 4460 -520
rect 4520 -580 4560 -520
rect 4420 -700 4560 -580
rect 5640 -320 5780 860
rect 6280 180 6380 200
rect 6280 120 6300 180
rect 6360 120 6380 180
rect 6280 80 6380 120
rect 6280 20 6300 80
rect 6360 20 6380 80
rect 6280 -20 6380 20
rect 6280 -80 6300 -20
rect 6360 -80 6380 -20
rect 6280 -100 6380 -80
rect 5640 -380 5680 -320
rect 5740 -380 5780 -320
rect 5640 -420 5780 -380
rect 5640 -480 5680 -420
rect 5740 -480 5780 -420
rect 5640 -520 5780 -480
rect 5640 -580 5680 -520
rect 5740 -580 5780 -520
rect 5640 -700 5780 -580
rect 6860 -320 7000 860
rect 7660 180 7760 200
rect 7660 120 7680 180
rect 7740 120 7760 180
rect 7660 80 7760 120
rect 7660 20 7680 80
rect 7740 20 7760 80
rect 7660 -20 7760 20
rect 7660 -80 7680 -20
rect 7740 -80 7760 -20
rect 7660 -100 7760 -80
rect 8100 180 8400 200
rect 8100 120 8120 180
rect 8180 120 8220 180
rect 8280 120 8320 180
rect 8380 120 8400 180
rect 8100 80 8400 120
rect 8100 20 8120 80
rect 8180 20 8220 80
rect 8280 20 8320 80
rect 8380 20 8400 80
rect 8100 -20 8400 20
rect 8100 -80 8120 -20
rect 8180 -80 8220 -20
rect 8280 -80 8320 -20
rect 8380 -80 8400 -20
rect 8100 -100 8400 -80
rect 6860 -380 6900 -320
rect 6960 -380 7000 -320
rect 6860 -420 7000 -380
rect 6860 -480 6900 -420
rect 6960 -480 7000 -420
rect 6860 -520 7000 -480
rect 6860 -580 6900 -520
rect 6960 -580 7000 -520
rect 6860 -700 7000 -580
rect 2100 -820 2200 -800
rect 2100 -880 2120 -820
rect 2180 -880 2200 -820
rect 2100 -900 2200 -880
rect 5000 -1620 5200 -1600
rect 5000 -1680 5020 -1620
rect 5080 -1680 5120 -1620
rect 5180 -1680 5200 -1620
rect 5000 -1720 5200 -1680
rect 5000 -1780 5020 -1720
rect 5080 -1780 5120 -1720
rect 5180 -1780 5200 -1720
rect 5000 -1800 5200 -1780
<< via1 >>
rect 1820 120 1880 180
rect 1920 120 1980 180
rect 2020 120 2080 180
rect 1820 20 1880 80
rect 1920 20 1980 80
rect 2020 20 2080 80
rect 1820 -80 1880 -20
rect 1920 -80 1980 -20
rect 2020 -80 2080 -20
rect 2440 120 2500 180
rect 2440 20 2500 80
rect 2440 -80 2500 -20
rect 3840 120 3900 180
rect 3840 20 3900 80
rect 3840 -80 3900 -20
rect 3220 -380 3280 -320
rect 3220 -480 3280 -420
rect 3220 -580 3280 -520
rect 5080 120 5140 180
rect 5080 20 5140 80
rect 5080 -80 5140 -20
rect 4460 -380 4520 -320
rect 4460 -480 4520 -420
rect 4460 -580 4520 -520
rect 6300 120 6360 180
rect 6300 20 6360 80
rect 6300 -80 6360 -20
rect 5680 -380 5740 -320
rect 5680 -480 5740 -420
rect 5680 -580 5740 -520
rect 7680 120 7740 180
rect 7680 20 7740 80
rect 7680 -80 7740 -20
rect 8120 120 8180 180
rect 8220 120 8280 180
rect 8320 120 8380 180
rect 8120 20 8180 80
rect 8220 20 8280 80
rect 8320 20 8380 80
rect 8120 -80 8180 -20
rect 8220 -80 8280 -20
rect 8320 -80 8380 -20
rect 6900 -380 6960 -320
rect 6900 -480 6960 -420
rect 6900 -580 6960 -520
rect 5020 -1680 5080 -1620
rect 5120 -1680 5180 -1620
rect 5020 -1780 5080 -1720
rect 5120 -1780 5180 -1720
<< metal2 >>
rect 1800 180 8400 200
rect 1800 120 1820 180
rect 1880 120 1920 180
rect 1980 120 2020 180
rect 2080 120 2440 180
rect 2500 120 3840 180
rect 3900 120 5080 180
rect 5140 120 6300 180
rect 6360 120 7680 180
rect 7740 120 8120 180
rect 8180 120 8220 180
rect 8280 120 8320 180
rect 8380 120 8400 180
rect 1800 80 8400 120
rect 1800 20 1820 80
rect 1880 20 1920 80
rect 1980 20 2020 80
rect 2080 20 2440 80
rect 2500 20 3840 80
rect 3900 20 5080 80
rect 5140 20 6300 80
rect 6360 20 7680 80
rect 7740 20 8120 80
rect 8180 20 8220 80
rect 8280 20 8320 80
rect 8380 20 8400 80
rect 1800 -20 8400 20
rect 1800 -80 1820 -20
rect 1880 -80 1920 -20
rect 1980 -80 2020 -20
rect 2080 -80 2440 -20
rect 2500 -80 3840 -20
rect 3900 -80 5080 -20
rect 5140 -80 6300 -20
rect 6360 -80 7680 -20
rect 7740 -80 8120 -20
rect 8180 -80 8220 -20
rect 8280 -80 8320 -20
rect 8380 -80 8400 -20
rect 1800 -100 8400 -80
rect 3100 -320 7100 -300
rect 3100 -380 3220 -320
rect 3280 -380 4460 -320
rect 4520 -380 5680 -320
rect 5740 -380 6900 -320
rect 6960 -380 7100 -320
rect 3100 -420 7100 -380
rect 3100 -480 3220 -420
rect 3280 -480 4460 -420
rect 4520 -480 5680 -420
rect 5740 -480 6900 -420
rect 6960 -480 7100 -420
rect 3100 -520 7100 -480
rect 3100 -580 3220 -520
rect 3280 -580 4460 -520
rect 4520 -580 5680 -520
rect 5740 -580 6900 -520
rect 6960 -580 7100 -520
rect 3100 -600 7100 -580
rect 5000 -1620 5200 -600
rect 5000 -1680 5020 -1620
rect 5080 -1680 5120 -1620
rect 5180 -1680 5200 -1620
rect 5000 -1720 5200 -1680
rect 5000 -1780 5020 -1720
rect 5080 -1780 5120 -1720
rect 5180 -1780 5200 -1720
rect 5000 -1800 5200 -1780
use sky130_fd_pr__nfet_g5v0d10v5_7GKDBD  XM6 /foss/designs/icdec-biomedical-pmic/xschem/error-amplifier/schematics/sub-blocks
timestamp 1770003475
transform 1 0 5101 0 1 107
box -2801 -807 2801 807
<< labels >>
flabel metal1 5000 -1800 5200 -1600 0 FreeSans 256 0 0 0 IBIAS
port 0 nsew
flabel metal1 2100 -900 2200 -800 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 1860 -40 2060 160 0 FreeSans 256 0 0 0 S
port 1 nsew
<< end >>
