magic
tech sky130A
magscale 1 2
timestamp 1770105080
<< mvnmos >>
rect -129 -444 -29 506
rect 29 -444 129 506
<< mvndiff >>
rect -187 494 -129 506
rect -187 -432 -175 494
rect -141 -432 -129 494
rect -187 -444 -129 -432
rect -29 494 29 506
rect -29 -432 -17 494
rect 17 -432 29 494
rect -29 -444 29 -432
rect 129 494 187 506
rect 129 -432 141 494
rect 175 -432 187 494
rect 129 -444 187 -432
<< mvndiffc >>
rect -175 -432 -141 494
rect -17 -432 17 494
rect 141 -432 175 494
<< poly >>
rect -129 506 -29 532
rect 29 506 129 532
rect -129 -482 -29 -444
rect -129 -516 -113 -482
rect -45 -516 -29 -482
rect -129 -532 -29 -516
rect 29 -482 129 -444
rect 29 -516 45 -482
rect 113 -516 129 -482
rect 29 -532 129 -516
<< polycont >>
rect -113 -516 -45 -482
rect 45 -516 113 -482
<< locali >>
rect -175 494 -141 510
rect -175 -448 -141 -432
rect -17 494 17 510
rect -17 -448 17 -432
rect 141 494 175 510
rect 141 -448 175 -432
rect -129 -516 -113 -482
rect -45 -516 -29 -482
rect 29 -516 45 -482
rect 113 -516 129 -482
<< viali >>
rect -175 -432 -141 494
rect -17 -432 17 494
rect 141 -432 175 494
rect -113 -516 -45 -482
rect 45 -516 113 -482
<< metal1 >>
rect -181 494 -135 506
rect -181 -432 -175 494
rect -141 -432 -135 494
rect -181 -444 -135 -432
rect -23 494 23 506
rect -23 -432 -17 494
rect 17 -432 23 494
rect -23 -444 23 -432
rect 135 494 181 506
rect 135 -432 141 494
rect 175 -432 181 494
rect 135 -444 181 -432
rect -125 -482 -33 -476
rect -125 -516 -113 -482
rect -45 -516 -33 -482
rect -125 -522 -33 -516
rect 33 -482 125 -476
rect 33 -516 45 -482
rect 113 -516 125 -482
rect 33 -522 125 -516
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.75 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
