magic
tech sky130A
magscale 1 2
timestamp 1769172933
<< nwell >>
rect 400 3800 13000 11200
<< pwell >>
rect 400 -1200 13000 3800
<< psubdiff >>
rect 3000 3400 10400 3600
rect 3000 2000 3200 3400
rect 4600 2000 4800 3400
rect 6600 2000 6800 3400
rect 8600 2000 8800 3400
rect 10200 2000 10400 3400
rect 600 1800 12800 2000
rect 4600 -600 4800 1800
rect 8600 -600 8800 1800
rect 12600 -600 12800 1800
rect 600 -800 12800 -600
<< nsubdiff >>
rect 2800 10800 10400 11000
rect 2800 7800 3000 10800
rect 10200 7800 10400 10800
rect 2200 7600 11200 7800
rect 2200 6000 2400 7600
rect 6600 6000 6800 7600
rect 11000 6000 11200 7600
rect 800 5800 12600 6000
rect 800 4200 1000 5800
rect 2200 4200 2400 5800
rect 6600 4200 6800 5800
rect 11000 4200 11200 5800
rect 12400 4200 12600 5800
rect 800 4000 12600 4200
<< locali >>
rect -11400 10800 24600 12400
rect 2800 7800 3000 10800
rect 10200 7800 10400 10800
rect 2200 7600 11200 7800
rect 2200 6000 2400 7600
rect 6600 6000 6800 7600
rect 11000 6000 11200 7600
rect 800 5800 12600 6000
rect 800 4200 1000 5800
rect 2200 4200 2400 5800
rect 6600 4200 6800 5800
rect 11000 4200 11200 5800
rect 12400 4200 12600 5800
rect 800 4000 12600 4200
rect 3000 3400 10400 3600
rect 3000 2000 3200 3400
rect 4600 2000 4800 3400
rect 6600 2000 6800 3400
rect 8600 2000 8800 3400
rect 10200 2000 10400 3400
rect 600 1800 12800 2000
rect 600 -600 800 1800
rect 4600 -600 4800 1800
rect 8600 -600 8800 1800
rect 12600 -600 12800 1800
rect -11200 -2200 24800 -600
<< metal1 >>
rect -11400 10800 24600 12400
rect -11200 -2200 24800 -600
rect 6000 -3400 6200 -3200
rect 6000 -3800 6200 -3600
rect 6600 -4000 6800 -3800
rect 6000 -4200 6200 -4000
<< metal2 >>
rect 0 -3800 800 3200
rect 1000 -400 12400 0
rect 6200 -4400 7200 -400
rect 12600 -3800 13400 3200
use sky130_fd_pr__cap_mim_m3_1_RK594X  sky130_fd_pr__cap_mim_m3_1_RK594X_0
timestamp 1769170640
transform 1 0 19092 0 1 4920
box -5492 -5320 5492 5320
use sky130_fd_pr__nfet_g5v0d10v5_686LLZ  sky130_fd_pr__nfet_g5v0d10v5_686LLZ_0
timestamp 1769172933
transform 1 0 6681 0 1 807
box -1681 -807 1681 807
use sky130_fd_pr__nfet_g5v0d10v5_686LLZ  sky130_fd_pr__nfet_g5v0d10v5_686LLZ_1
timestamp 1769172933
transform 1 0 10681 0 1 807
box -1681 -807 1681 807
use sky130_fd_pr__nfet_g5v0d10v5_B9VV4Y  sky130_fd_pr__nfet_g5v0d10v5_B9VV4Y_0
timestamp 1769172933
transform 1 0 9525 0 1 2728
box -525 -528 525 528
use sky130_fd_pr__nfet_g5v0d10v5_B9VV4Y  sky130_fd_pr__nfet_g5v0d10v5_B9VV4Y_3
timestamp 1769172933
transform 1 0 3925 0 1 2728
box -525 -528 525 528
use sky130_fd_pr__nfet_g5v0d10v5_TJAW4Y  sky130_fd_pr__nfet_g5v0d10v5_TJAW4Y_0
timestamp 1769172933
transform 1 0 5725 0 1 2728
box -525 -528 525 528
use sky130_fd_pr__nfet_g5v0d10v5_TJAW4Y  sky130_fd_pr__nfet_g5v0d10v5_TJAW4Y_1
timestamp 1769172933
transform 1 0 7725 0 1 2728
box -525 -528 525 528
use sky130_fd_pr__pfet_g5v0d10v5_AXLSKB  sky130_fd_pr__pfet_g5v0d10v5_AXLSKB_0
timestamp 1769172933
transform 1 0 1593 0 1 4964
box -393 -564 393 602
use sky130_fd_pr__pfet_g5v0d10v5_HENH7L  sky130_fd_pr__pfet_g5v0d10v5_HENH7L_0
timestamp 1769170640
transform 1 0 6659 0 1 9464
box -3459 -1064 3459 1102
use sky130_fd_pr__pfet_g5v0d10v5_UABD3S  sky130_fd_pr__pfet_g5v0d10v5_UABD3S_0
timestamp 1769172933
transform 1 0 4347 0 1 6772
box -1747 -572 1747 534
use sky130_fd_pr__pfet_g5v0d10v5_UABD3S  sky130_fd_pr__pfet_g5v0d10v5_UABD3S_1
timestamp 1769172933
transform 1 0 9147 0 1 6772
box -1747 -572 1747 534
use sky130_fd_pr__pfet_g5v0d10v5_UABDA8  sky130_fd_pr__pfet_g5v0d10v5_UABDA8_0
timestamp 1769172933
transform 1 0 4347 0 1 4934
box -1747 -534 1747 572
use sky130_fd_pr__pfet_g5v0d10v5_UABDA8  sky130_fd_pr__pfet_g5v0d10v5_UABDA8_1
timestamp 1769172933
transform 1 0 9147 0 1 4934
box -1747 -534 1747 572
use sky130_fd_pr__cap_mim_m3_1_RK594X  XC1
timestamp 1769170640
transform 1 0 -5908 0 1 5120
box -5492 -5320 5492 5320
use sky130_fd_pr__nfet_g5v0d10v5_686LLZ  XM5
timestamp 1769172933
transform 1 0 2681 0 1 807
box -1681 -807 1681 807
use sky130_fd_pr__pfet_g5v0d10v5_AXLSKB  XM9
timestamp 1769172933
transform 1 0 11793 0 1 4964
box -393 -564 393 602
<< labels >>
flabel metal1 -10600 -2000 -10400 -1800 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 -10800 11400 -10600 11600 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 6000 -3400 6200 -3200 0 FreeSans 256 0 0 0 VP
port 2 nsew
flabel metal1 6000 -3800 6200 -3600 0 FreeSans 256 0 0 0 VN
port 3 nsew
flabel metal1 6000 -4200 6200 -4000 0 FreeSans 256 0 0 0 IBIAS
port 4 nsew
flabel metal1 6600 -4000 6800 -3800 0 FreeSans 256 0 0 0 OUT
port 1 nsew
<< end >>
