** sch_path: /foss/designs/icdec-biomedical-pmic/xschem/error-amplifier2/schematics/1st-stage.sch
.subckt 1st-stage VDD VP VN IBIAS VSS OUT
*.PININFO VDD:B VP:I VN:I IBIAS:I VSS:B OUT:O
XM1 net2 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.25 W=75.2 nf=8 m=1
XM2 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.25 W=75.2 nf=8 m=1
XM3 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=18.8 nf=2 m=1
XM4 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=18.8 nf=2 m=1
XM5 net2 VN net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=38 nf=2 m=1
XM6 net1 VP net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=38 nf=2 m=1
XM7 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM8 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM9 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM10 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM11 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM12 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM13 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM14 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM15 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM16 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM17 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM18 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM19 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM20 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM21 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM22 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=9.5 nf=2 m=1
XM23 net3 IBIAS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1.25 W=60 nf=4 m=1
XM24 IBIAS IBIAS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1.25 W=60 nf=4 m=1
XM25 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=15 nf=2 m=1
XM26 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=15 nf=2 m=1
XM27 OUT net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.25 W=160 nf=16 m=1
XM28 OUT IBIAS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1.25 W=60 nf=8 m=1
XC1 net4 net2 sky130_fd_pr__cap_mim_m3_1 W=25 L=25 m=8
XM29 OUT VSS net4 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.9 W=20 nf=4 m=1
.ends
