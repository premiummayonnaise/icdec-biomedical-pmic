magic
tech sky130A
magscale 1 2
timestamp 1770035380
<< error_p >>
rect -2344 791 -2276 797
rect -2036 791 -1968 797
rect -1728 791 -1660 797
rect -1420 791 -1352 797
rect -1112 791 -1044 797
rect -804 791 -736 797
rect -496 791 -428 797
rect -188 791 -120 797
rect 120 791 188 797
rect 428 791 496 797
rect 736 791 804 797
rect 1044 791 1112 797
rect 1352 791 1420 797
rect 1660 791 1728 797
rect 1968 791 2036 797
rect 2276 791 2344 797
rect -2344 757 -2332 791
rect -2036 757 -2024 791
rect -1728 757 -1716 791
rect -1420 757 -1408 791
rect -1112 757 -1100 791
rect -804 757 -792 791
rect -496 757 -484 791
rect -188 757 -176 791
rect 120 757 132 791
rect 428 757 440 791
rect 736 757 748 791
rect 1044 757 1056 791
rect 1352 757 1364 791
rect 1660 757 1672 791
rect 1968 757 1980 791
rect 2276 757 2288 791
rect -2344 751 -2276 757
rect -2036 751 -1968 757
rect -1728 751 -1660 757
rect -1420 751 -1352 757
rect -1112 751 -1044 757
rect -804 751 -736 757
rect -496 751 -428 757
rect -188 751 -120 757
rect 120 751 188 757
rect 428 751 496 757
rect 736 751 804 757
rect 1044 751 1112 757
rect 1352 751 1420 757
rect 1660 751 1728 757
rect 1968 751 2036 757
rect 2276 751 2344 757
<< mvnmos >>
rect -2435 -781 -2185 719
rect -2127 -781 -1877 719
rect -1819 -781 -1569 719
rect -1511 -781 -1261 719
rect -1203 -781 -953 719
rect -895 -781 -645 719
rect -587 -781 -337 719
rect -279 -781 -29 719
rect 29 -781 279 719
rect 337 -781 587 719
rect 645 -781 895 719
rect 953 -781 1203 719
rect 1261 -781 1511 719
rect 1569 -781 1819 719
rect 1877 -781 2127 719
rect 2185 -781 2435 719
<< mvndiff >>
rect -2493 707 -2435 719
rect -2493 -769 -2481 707
rect -2447 -769 -2435 707
rect -2493 -781 -2435 -769
rect -2185 707 -2127 719
rect -2185 -769 -2173 707
rect -2139 -769 -2127 707
rect -2185 -781 -2127 -769
rect -1877 707 -1819 719
rect -1877 -769 -1865 707
rect -1831 -769 -1819 707
rect -1877 -781 -1819 -769
rect -1569 707 -1511 719
rect -1569 -769 -1557 707
rect -1523 -769 -1511 707
rect -1569 -781 -1511 -769
rect -1261 707 -1203 719
rect -1261 -769 -1249 707
rect -1215 -769 -1203 707
rect -1261 -781 -1203 -769
rect -953 707 -895 719
rect -953 -769 -941 707
rect -907 -769 -895 707
rect -953 -781 -895 -769
rect -645 707 -587 719
rect -645 -769 -633 707
rect -599 -769 -587 707
rect -645 -781 -587 -769
rect -337 707 -279 719
rect -337 -769 -325 707
rect -291 -769 -279 707
rect -337 -781 -279 -769
rect -29 707 29 719
rect -29 -769 -17 707
rect 17 -769 29 707
rect -29 -781 29 -769
rect 279 707 337 719
rect 279 -769 291 707
rect 325 -769 337 707
rect 279 -781 337 -769
rect 587 707 645 719
rect 587 -769 599 707
rect 633 -769 645 707
rect 587 -781 645 -769
rect 895 707 953 719
rect 895 -769 907 707
rect 941 -769 953 707
rect 895 -781 953 -769
rect 1203 707 1261 719
rect 1203 -769 1215 707
rect 1249 -769 1261 707
rect 1203 -781 1261 -769
rect 1511 707 1569 719
rect 1511 -769 1523 707
rect 1557 -769 1569 707
rect 1511 -781 1569 -769
rect 1819 707 1877 719
rect 1819 -769 1831 707
rect 1865 -769 1877 707
rect 1819 -781 1877 -769
rect 2127 707 2185 719
rect 2127 -769 2139 707
rect 2173 -769 2185 707
rect 2127 -781 2185 -769
rect 2435 707 2493 719
rect 2435 -769 2447 707
rect 2481 -769 2493 707
rect 2435 -781 2493 -769
<< mvndiffc >>
rect -2481 -769 -2447 707
rect -2173 -769 -2139 707
rect -1865 -769 -1831 707
rect -1557 -769 -1523 707
rect -1249 -769 -1215 707
rect -941 -769 -907 707
rect -633 -769 -599 707
rect -325 -769 -291 707
rect -17 -769 17 707
rect 291 -769 325 707
rect 599 -769 633 707
rect 907 -769 941 707
rect 1215 -769 1249 707
rect 1523 -769 1557 707
rect 1831 -769 1865 707
rect 2139 -769 2173 707
rect 2447 -769 2481 707
<< poly >>
rect -2348 791 -2272 807
rect -2348 774 -2332 791
rect -2435 757 -2332 774
rect -2288 774 -2272 791
rect -2040 791 -1964 807
rect -2040 774 -2024 791
rect -2288 757 -2185 774
rect -2435 719 -2185 757
rect -2127 757 -2024 774
rect -1980 774 -1964 791
rect -1732 791 -1656 807
rect -1732 774 -1716 791
rect -1980 757 -1877 774
rect -2127 719 -1877 757
rect -1819 757 -1716 774
rect -1672 774 -1656 791
rect -1424 791 -1348 807
rect -1424 774 -1408 791
rect -1672 757 -1569 774
rect -1819 719 -1569 757
rect -1511 757 -1408 774
rect -1364 774 -1348 791
rect -1116 791 -1040 807
rect -1116 774 -1100 791
rect -1364 757 -1261 774
rect -1511 719 -1261 757
rect -1203 757 -1100 774
rect -1056 774 -1040 791
rect -808 791 -732 807
rect -808 774 -792 791
rect -1056 757 -953 774
rect -1203 719 -953 757
rect -895 757 -792 774
rect -748 774 -732 791
rect -500 791 -424 807
rect -500 774 -484 791
rect -748 757 -645 774
rect -895 719 -645 757
rect -587 757 -484 774
rect -440 774 -424 791
rect -192 791 -116 807
rect -192 774 -176 791
rect -440 757 -337 774
rect -587 719 -337 757
rect -279 757 -176 774
rect -132 774 -116 791
rect 116 791 192 807
rect 116 774 132 791
rect -132 757 -29 774
rect -279 719 -29 757
rect 29 757 132 774
rect 176 774 192 791
rect 424 791 500 807
rect 424 774 440 791
rect 176 757 279 774
rect 29 719 279 757
rect 337 757 440 774
rect 484 774 500 791
rect 732 791 808 807
rect 732 774 748 791
rect 484 757 587 774
rect 337 719 587 757
rect 645 757 748 774
rect 792 774 808 791
rect 1040 791 1116 807
rect 1040 774 1056 791
rect 792 757 895 774
rect 645 719 895 757
rect 953 757 1056 774
rect 1100 774 1116 791
rect 1348 791 1424 807
rect 1348 774 1364 791
rect 1100 757 1203 774
rect 953 719 1203 757
rect 1261 757 1364 774
rect 1408 774 1424 791
rect 1656 791 1732 807
rect 1656 774 1672 791
rect 1408 757 1511 774
rect 1261 719 1511 757
rect 1569 757 1672 774
rect 1716 774 1732 791
rect 1964 791 2040 807
rect 1964 774 1980 791
rect 1716 757 1819 774
rect 1569 719 1819 757
rect 1877 757 1980 774
rect 2024 774 2040 791
rect 2272 791 2348 807
rect 2272 774 2288 791
rect 2024 757 2127 774
rect 1877 719 2127 757
rect 2185 757 2288 774
rect 2332 774 2348 791
rect 2332 757 2435 774
rect 2185 719 2435 757
rect -2435 -807 -2185 -781
rect -2127 -807 -1877 -781
rect -1819 -807 -1569 -781
rect -1511 -807 -1261 -781
rect -1203 -807 -953 -781
rect -895 -807 -645 -781
rect -587 -807 -337 -781
rect -279 -807 -29 -781
rect 29 -807 279 -781
rect 337 -807 587 -781
rect 645 -807 895 -781
rect 953 -807 1203 -781
rect 1261 -807 1511 -781
rect 1569 -807 1819 -781
rect 1877 -807 2127 -781
rect 2185 -807 2435 -781
<< polycont >>
rect -2332 757 -2288 791
rect -2024 757 -1980 791
rect -1716 757 -1672 791
rect -1408 757 -1364 791
rect -1100 757 -1056 791
rect -792 757 -748 791
rect -484 757 -440 791
rect -176 757 -132 791
rect 132 757 176 791
rect 440 757 484 791
rect 748 757 792 791
rect 1056 757 1100 791
rect 1364 757 1408 791
rect 1672 757 1716 791
rect 1980 757 2024 791
rect 2288 757 2332 791
<< locali >>
rect -2348 757 -2332 791
rect -2288 757 -2272 791
rect -2040 757 -2024 791
rect -1980 757 -1964 791
rect -1732 757 -1716 791
rect -1672 757 -1656 791
rect -1424 757 -1408 791
rect -1364 757 -1348 791
rect -1116 757 -1100 791
rect -1056 757 -1040 791
rect -808 757 -792 791
rect -748 757 -732 791
rect -500 757 -484 791
rect -440 757 -424 791
rect -192 757 -176 791
rect -132 757 -116 791
rect 116 757 132 791
rect 176 757 192 791
rect 424 757 440 791
rect 484 757 500 791
rect 732 757 748 791
rect 792 757 808 791
rect 1040 757 1056 791
rect 1100 757 1116 791
rect 1348 757 1364 791
rect 1408 757 1424 791
rect 1656 757 1672 791
rect 1716 757 1732 791
rect 1964 757 1980 791
rect 2024 757 2040 791
rect 2272 757 2288 791
rect 2332 757 2348 791
rect -2481 707 -2447 723
rect -2481 -785 -2447 -769
rect -2173 707 -2139 723
rect -2173 -785 -2139 -769
rect -1865 707 -1831 723
rect -1865 -785 -1831 -769
rect -1557 707 -1523 723
rect -1557 -785 -1523 -769
rect -1249 707 -1215 723
rect -1249 -785 -1215 -769
rect -941 707 -907 723
rect -941 -785 -907 -769
rect -633 707 -599 723
rect -633 -785 -599 -769
rect -325 707 -291 723
rect -325 -785 -291 -769
rect -17 707 17 723
rect -17 -785 17 -769
rect 291 707 325 723
rect 291 -785 325 -769
rect 599 707 633 723
rect 599 -785 633 -769
rect 907 707 941 723
rect 907 -785 941 -769
rect 1215 707 1249 723
rect 1215 -785 1249 -769
rect 1523 707 1557 723
rect 1523 -785 1557 -769
rect 1831 707 1865 723
rect 1831 -785 1865 -769
rect 2139 707 2173 723
rect 2139 -785 2173 -769
rect 2447 707 2481 723
rect 2447 -785 2481 -769
<< viali >>
rect -2332 757 -2288 791
rect -2024 757 -1980 791
rect -1716 757 -1672 791
rect -1408 757 -1364 791
rect -1100 757 -1056 791
rect -792 757 -748 791
rect -484 757 -440 791
rect -176 757 -132 791
rect 132 757 176 791
rect 440 757 484 791
rect 748 757 792 791
rect 1056 757 1100 791
rect 1364 757 1408 791
rect 1672 757 1716 791
rect 1980 757 2024 791
rect 2288 757 2332 791
rect -2481 -769 -2447 707
rect -2173 -769 -2139 707
rect -1865 -769 -1831 707
rect -1557 -769 -1523 707
rect -1249 -769 -1215 707
rect -941 -769 -907 707
rect -633 -769 -599 707
rect -325 -769 -291 707
rect -17 -769 17 707
rect 291 -769 325 707
rect 599 -769 633 707
rect 907 -769 941 707
rect 1215 -769 1249 707
rect 1523 -769 1557 707
rect 1831 -769 1865 707
rect 2139 -769 2173 707
rect 2447 -769 2481 707
<< metal1 >>
rect -2344 791 -2276 797
rect -2344 757 -2332 791
rect -2288 757 -2276 791
rect -2344 751 -2276 757
rect -2036 791 -1968 797
rect -2036 757 -2024 791
rect -1980 757 -1968 791
rect -2036 751 -1968 757
rect -1728 791 -1660 797
rect -1728 757 -1716 791
rect -1672 757 -1660 791
rect -1728 751 -1660 757
rect -1420 791 -1352 797
rect -1420 757 -1408 791
rect -1364 757 -1352 791
rect -1420 751 -1352 757
rect -1112 791 -1044 797
rect -1112 757 -1100 791
rect -1056 757 -1044 791
rect -1112 751 -1044 757
rect -804 791 -736 797
rect -804 757 -792 791
rect -748 757 -736 791
rect -804 751 -736 757
rect -496 791 -428 797
rect -496 757 -484 791
rect -440 757 -428 791
rect -496 751 -428 757
rect -188 791 -120 797
rect -188 757 -176 791
rect -132 757 -120 791
rect -188 751 -120 757
rect 120 791 188 797
rect 120 757 132 791
rect 176 757 188 791
rect 120 751 188 757
rect 428 791 496 797
rect 428 757 440 791
rect 484 757 496 791
rect 428 751 496 757
rect 736 791 804 797
rect 736 757 748 791
rect 792 757 804 791
rect 736 751 804 757
rect 1044 791 1112 797
rect 1044 757 1056 791
rect 1100 757 1112 791
rect 1044 751 1112 757
rect 1352 791 1420 797
rect 1352 757 1364 791
rect 1408 757 1420 791
rect 1352 751 1420 757
rect 1660 791 1728 797
rect 1660 757 1672 791
rect 1716 757 1728 791
rect 1660 751 1728 757
rect 1968 791 2036 797
rect 1968 757 1980 791
rect 2024 757 2036 791
rect 1968 751 2036 757
rect 2276 791 2344 797
rect 2276 757 2288 791
rect 2332 757 2344 791
rect 2276 751 2344 757
rect -2487 707 -2441 719
rect -2487 -769 -2481 707
rect -2447 -769 -2441 707
rect -2487 -781 -2441 -769
rect -2179 707 -2133 719
rect -2179 -769 -2173 707
rect -2139 -769 -2133 707
rect -2179 -781 -2133 -769
rect -1871 707 -1825 719
rect -1871 -769 -1865 707
rect -1831 -769 -1825 707
rect -1871 -781 -1825 -769
rect -1563 707 -1517 719
rect -1563 -769 -1557 707
rect -1523 -769 -1517 707
rect -1563 -781 -1517 -769
rect -1255 707 -1209 719
rect -1255 -769 -1249 707
rect -1215 -769 -1209 707
rect -1255 -781 -1209 -769
rect -947 707 -901 719
rect -947 -769 -941 707
rect -907 -769 -901 707
rect -947 -781 -901 -769
rect -639 707 -593 719
rect -639 -769 -633 707
rect -599 -769 -593 707
rect -639 -781 -593 -769
rect -331 707 -285 719
rect -331 -769 -325 707
rect -291 -769 -285 707
rect -331 -781 -285 -769
rect -23 707 23 719
rect -23 -769 -17 707
rect 17 200 23 707
rect 285 707 331 719
rect 17 0 200 200
rect 17 -200 23 0
rect 17 -400 200 -200
rect 17 -600 23 -400
rect 17 -769 200 -600
rect -23 -781 200 -769
rect 285 -769 291 707
rect 325 -769 331 707
rect 285 -781 331 -769
rect 593 707 639 719
rect 593 -769 599 707
rect 633 -769 639 707
rect 593 -781 639 -769
rect 901 707 947 719
rect 901 -769 907 707
rect 941 -769 947 707
rect 901 -781 947 -769
rect 1209 707 1255 719
rect 1209 -769 1215 707
rect 1249 -769 1255 707
rect 1209 -781 1255 -769
rect 1517 707 1563 719
rect 1517 -769 1523 707
rect 1557 -769 1563 707
rect 1517 -781 1563 -769
rect 1825 707 1871 719
rect 1825 -769 1831 707
rect 1865 -769 1871 707
rect 1825 -781 1871 -769
rect 2133 707 2179 719
rect 2133 -769 2139 707
rect 2173 -769 2179 707
rect 2133 -781 2179 -769
rect 2441 707 2487 719
rect 2441 -769 2447 707
rect 2481 -769 2487 707
rect 2441 -781 2487 -769
rect 0 -800 200 -781
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
rect 0 -8800 200 -8600
rect 0 -9200 200 -9000
rect 0 -9600 200 -9400
rect 0 -10000 200 -9800
rect 0 -10400 200 -10200
rect 0 -10800 200 -10600
rect 0 -11200 200 -11000
rect 0 -11600 200 -11400
rect 0 -12000 200 -11800
rect 0 -12400 200 -12200
rect 0 -12800 200 -12600
rect 0 -13200 200 -13000
rect 0 -13600 200 -13400
rect 0 -14000 200 -13800
rect 0 -14400 200 -14200
rect 0 -14800 200 -14600
rect 0 -15200 200 -15000
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X0
timestamp 0
transform 1 0 -2205 0 1 -14257
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X1
timestamp 0
transform 1 0 -1564 0 1 -14322
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X2
timestamp 0
transform 1 0 -923 0 1 -14387
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X3
timestamp 0
transform 1 0 -282 0 1 -14452
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X4
timestamp 0
transform 1 0 359 0 1 -14517
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X5
timestamp 0
transform 1 0 1000 0 1 -14582
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X6
timestamp 0
transform 1 0 1641 0 1 -14647
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X7
timestamp 0
transform 1 0 2282 0 1 -14712
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X8
timestamp 0
transform 1 0 2923 0 1 -14777
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_XZ8YPJ  X9
timestamp 0
transform 1 0 3564 0 1 -14842
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_X6YUYU  X10
timestamp 0
transform 1 0 4205 0 1 -14907
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X11
timestamp 0
transform 1 0 4846 0 1 -14972
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X12
timestamp 0
transform 1 0 5487 0 1 -15037
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X13
timestamp 0
transform 1 0 6128 0 1 -15102
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X14
timestamp 0
transform 1 0 6769 0 1 -15167
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X15
timestamp 0
transform 1 0 7410 0 1 -15232
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 a_n953_n781#
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 a_2185_n807#
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 a_n587_n807#
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 {}
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 a_645_n807#
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 a_29_n807#
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 a_2435_n781#
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 a_n2185_n781#
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 a_1261_n807#
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 a_1569_n807#
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 a_279_n781#
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 a_895_n781#
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 a_n2435_n807#
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 a_n1261_n781#
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 a_1511_n781#
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 a_1819_n781#
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 a_n1569_n781#
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 {}
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 a_n29_n781#
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 a_n645_n781#
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 256 0 0 0 a_n1511_n807#
port 21 nsew
flabel metal1 0 -8800 200 -8600 0 FreeSans 256 0 0 0 a_n279_n807#
port 22 nsew
flabel metal1 0 -9200 200 -9000 0 FreeSans 256 0 0 0 a_n1819_n807#
port 23 nsew
flabel metal1 0 -9600 200 -9400 0 FreeSans 256 0 0 0 a_n895_n807#
port 24 nsew
flabel metal1 0 -10000 200 -9800 0 FreeSans 256 0 0 0 a_337_n807#
port 25 nsew
flabel metal1 0 -10400 200 -10200 0 FreeSans 256 0 0 0 {}
port 26 nsew
flabel metal1 0 -10800 200 -10600 0 FreeSans 256 0 0 0 a_953_n807#
port 27 nsew
flabel metal1 0 -11200 200 -11000 0 FreeSans 256 0 0 0 a_2127_n781#
port 28 nsew
flabel metal1 0 -11600 200 -11400 0 FreeSans 256 0 0 0 a_n2493_n781#
port 29 nsew
flabel metal1 0 -12000 200 -11800 0 FreeSans 256 0 0 0 a_587_n781#
port 30 nsew
flabel metal1 0 -12400 200 -12200 0 FreeSans 256 0 0 0 a_1877_n807#
port 31 nsew
flabel metal1 0 -12800 200 -12600 0 FreeSans 256 0 0 0 a_n2127_n807#
port 32 nsew
flabel metal1 0 -13200 200 -13000 0 FreeSans 256 0 0 0 a_1203_n781#
port 33 nsew
flabel metal1 0 -13600 200 -13400 0 FreeSans 256 0 0 0 {}
port 34 nsew
flabel metal1 0 -14000 200 -13800 0 FreeSans 256 0 0 0 a_n1877_n781#
port 35 nsew
flabel metal1 0 -14400 200 -14200 0 FreeSans 256 0 0 0 a_n337_n781#
port 36 nsew
flabel metal1 0 -14800 200 -14600 0 FreeSans 256 0 0 0 a_n1203_n807#
port 37 nsew
flabel metal1 0 -15200 200 -15000 0 FreeSans 256 0 0 0 VSUBS
port 38 nsew
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 16 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
