magic
tech sky130A
magscale 1 2
timestamp 1770023980
<< metal4 >>
rect -5898 10639 -200 10680
rect -5898 5561 -456 10639
rect -220 5561 -200 10639
rect -5898 5520 -200 5561
rect 200 10639 5898 10680
rect 200 5561 5642 10639
rect 5878 5561 5898 10639
rect 200 5520 5898 5561
rect -5898 5239 -200 5280
rect -5898 161 -456 5239
rect -220 161 -200 5239
rect -5898 120 -200 161
rect 200 5239 5898 5280
rect 200 161 5642 5239
rect 5878 161 5898 5239
rect 200 120 5898 161
rect -5898 -161 -200 -120
rect -5898 -5239 -456 -161
rect -220 -5239 -200 -161
rect -5898 -5280 -200 -5239
rect 200 -161 5898 -120
rect 200 -5239 5642 -161
rect 5878 -5239 5898 -161
rect 200 -5280 5898 -5239
rect -5898 -5561 -200 -5520
rect -5898 -10639 -456 -5561
rect -220 -10639 -200 -5561
rect -5898 -10680 -200 -10639
rect 200 -5561 5898 -5520
rect 200 -10639 5642 -5561
rect 5878 -10639 5898 -5561
rect 200 -10680 5898 -10639
<< via4 >>
rect -456 5561 -220 10639
rect 5642 5561 5878 10639
rect -456 161 -220 5239
rect 5642 161 5878 5239
rect -456 -5239 -220 -161
rect 5642 -5239 5878 -161
rect -456 -10639 -220 -5561
rect 5642 -10639 5878 -5561
<< mimcap2 >>
rect -5818 10560 -818 10600
rect -5818 5640 -5778 10560
rect -858 5640 -818 10560
rect -5818 5600 -818 5640
rect 280 10560 5280 10600
rect 280 5640 320 10560
rect 5240 5640 5280 10560
rect 280 5600 5280 5640
rect -5818 5160 -818 5200
rect -5818 240 -5778 5160
rect -858 240 -818 5160
rect -5818 200 -818 240
rect 280 5160 5280 5200
rect 280 240 320 5160
rect 5240 240 5280 5160
rect 280 200 5280 240
rect -5818 -240 -818 -200
rect -5818 -5160 -5778 -240
rect -858 -5160 -818 -240
rect -5818 -5200 -818 -5160
rect 280 -240 5280 -200
rect 280 -5160 320 -240
rect 5240 -5160 5280 -240
rect 280 -5200 5280 -5160
rect -5818 -5640 -818 -5600
rect -5818 -10560 -5778 -5640
rect -858 -10560 -818 -5640
rect -5818 -10600 -818 -10560
rect 280 -5640 5280 -5600
rect 280 -10560 320 -5640
rect 5240 -10560 5280 -5640
rect 280 -10600 5280 -10560
<< mimcap2contact >>
rect -5778 5640 -858 10560
rect 320 5640 5240 10560
rect -5778 240 -858 5160
rect 320 240 5240 5160
rect -5778 -5160 -858 -240
rect 320 -5160 5240 -240
rect -5778 -10560 -858 -5640
rect 320 -10560 5240 -5640
<< metal5 >>
rect -3478 10584 -3158 10800
rect -498 10639 -178 10800
rect -5802 10560 -834 10584
rect -5802 5640 -5778 10560
rect -858 5640 -834 10560
rect -5802 5616 -834 5640
rect -3478 5184 -3158 5616
rect -498 5561 -456 10639
rect -220 5561 -178 10639
rect 2620 10584 2940 10800
rect 5600 10639 5920 10800
rect 296 10560 5264 10584
rect 296 5640 320 10560
rect 5240 5640 5264 10560
rect 296 5616 5264 5640
rect -498 5239 -178 5561
rect -5802 5160 -834 5184
rect -5802 240 -5778 5160
rect -858 240 -834 5160
rect -5802 216 -834 240
rect -3478 -216 -3158 216
rect -498 161 -456 5239
rect -220 161 -178 5239
rect 2620 5184 2940 5616
rect 5600 5561 5642 10639
rect 5878 5561 5920 10639
rect 5600 5239 5920 5561
rect 296 5160 5264 5184
rect 296 240 320 5160
rect 5240 240 5264 5160
rect 296 216 5264 240
rect -498 -161 -178 161
rect -5802 -240 -834 -216
rect -5802 -5160 -5778 -240
rect -858 -5160 -834 -240
rect -5802 -5184 -834 -5160
rect -3478 -5616 -3158 -5184
rect -498 -5239 -456 -161
rect -220 -5239 -178 -161
rect 2620 -216 2940 216
rect 5600 161 5642 5239
rect 5878 161 5920 5239
rect 5600 -161 5920 161
rect 296 -240 5264 -216
rect 296 -5160 320 -240
rect 5240 -5160 5264 -240
rect 296 -5184 5264 -5160
rect -498 -5561 -178 -5239
rect -5802 -5640 -834 -5616
rect -5802 -10560 -5778 -5640
rect -858 -10560 -834 -5640
rect -5802 -10584 -834 -10560
rect -3478 -10800 -3158 -10584
rect -498 -10639 -456 -5561
rect -220 -10639 -178 -5561
rect 2620 -5616 2940 -5184
rect 5600 -5239 5642 -161
rect 5878 -5239 5920 -161
rect 5600 -5561 5920 -5239
rect 296 -5640 5264 -5616
rect 296 -10560 320 -5640
rect 5240 -10560 5264 -5640
rect 296 -10584 5264 -10560
rect -498 -10800 -178 -10639
rect 2620 -10800 2940 -10584
rect 5600 -10639 5642 -5561
rect 5878 -10639 5920 -5561
rect 5600 -10800 5920 -10639
<< properties >>
string FIXED_BBOX 200 5520 5360 10680
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25 l 25 val 1.269k carea 2.00 cperi 0.19 class capacitor nx 2 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
