magic
tech sky130A
magscale 1 2
timestamp 1770083657
<< pwell >>
rect -2827 -807 2827 745
<< mvnmos >>
rect -2743 -781 -2493 719
rect -2435 -781 -2185 719
rect -2127 -781 -1877 719
rect -1819 -781 -1569 719
rect -1511 -781 -1261 719
rect -1203 -781 -953 719
rect -895 -781 -645 719
rect -587 -781 -337 719
rect -279 -781 -29 719
rect 29 -781 279 719
rect 337 -781 587 719
rect 645 -781 895 719
rect 953 -781 1203 719
rect 1261 -781 1511 719
rect 1569 -781 1819 719
rect 1877 -781 2127 719
rect 2185 -781 2435 719
rect 2493 -781 2743 719
<< mvndiff >>
rect -2801 700 -2743 719
rect -2801 666 -2789 700
rect -2755 666 -2743 700
rect -2801 632 -2743 666
rect -2801 598 -2789 632
rect -2755 598 -2743 632
rect -2801 564 -2743 598
rect -2801 530 -2789 564
rect -2755 530 -2743 564
rect -2801 496 -2743 530
rect -2801 462 -2789 496
rect -2755 462 -2743 496
rect -2801 428 -2743 462
rect -2801 394 -2789 428
rect -2755 394 -2743 428
rect -2801 360 -2743 394
rect -2801 326 -2789 360
rect -2755 326 -2743 360
rect -2801 292 -2743 326
rect -2801 258 -2789 292
rect -2755 258 -2743 292
rect -2801 224 -2743 258
rect -2801 190 -2789 224
rect -2755 190 -2743 224
rect -2801 156 -2743 190
rect -2801 122 -2789 156
rect -2755 122 -2743 156
rect -2801 88 -2743 122
rect -2801 54 -2789 88
rect -2755 54 -2743 88
rect -2801 20 -2743 54
rect -2801 -14 -2789 20
rect -2755 -14 -2743 20
rect -2801 -48 -2743 -14
rect -2801 -82 -2789 -48
rect -2755 -82 -2743 -48
rect -2801 -116 -2743 -82
rect -2801 -150 -2789 -116
rect -2755 -150 -2743 -116
rect -2801 -184 -2743 -150
rect -2801 -218 -2789 -184
rect -2755 -218 -2743 -184
rect -2801 -252 -2743 -218
rect -2801 -286 -2789 -252
rect -2755 -286 -2743 -252
rect -2801 -320 -2743 -286
rect -2801 -354 -2789 -320
rect -2755 -354 -2743 -320
rect -2801 -388 -2743 -354
rect -2801 -422 -2789 -388
rect -2755 -422 -2743 -388
rect -2801 -456 -2743 -422
rect -2801 -490 -2789 -456
rect -2755 -490 -2743 -456
rect -2801 -524 -2743 -490
rect -2801 -558 -2789 -524
rect -2755 -558 -2743 -524
rect -2801 -592 -2743 -558
rect -2801 -626 -2789 -592
rect -2755 -626 -2743 -592
rect -2801 -660 -2743 -626
rect -2801 -694 -2789 -660
rect -2755 -694 -2743 -660
rect -2801 -728 -2743 -694
rect -2801 -762 -2789 -728
rect -2755 -762 -2743 -728
rect -2801 -781 -2743 -762
rect -2493 700 -2435 719
rect -2493 666 -2481 700
rect -2447 666 -2435 700
rect -2493 632 -2435 666
rect -2493 598 -2481 632
rect -2447 598 -2435 632
rect -2493 564 -2435 598
rect -2493 530 -2481 564
rect -2447 530 -2435 564
rect -2493 496 -2435 530
rect -2493 462 -2481 496
rect -2447 462 -2435 496
rect -2493 428 -2435 462
rect -2493 394 -2481 428
rect -2447 394 -2435 428
rect -2493 360 -2435 394
rect -2493 326 -2481 360
rect -2447 326 -2435 360
rect -2493 292 -2435 326
rect -2493 258 -2481 292
rect -2447 258 -2435 292
rect -2493 224 -2435 258
rect -2493 190 -2481 224
rect -2447 190 -2435 224
rect -2493 156 -2435 190
rect -2493 122 -2481 156
rect -2447 122 -2435 156
rect -2493 88 -2435 122
rect -2493 54 -2481 88
rect -2447 54 -2435 88
rect -2493 20 -2435 54
rect -2493 -14 -2481 20
rect -2447 -14 -2435 20
rect -2493 -48 -2435 -14
rect -2493 -82 -2481 -48
rect -2447 -82 -2435 -48
rect -2493 -116 -2435 -82
rect -2493 -150 -2481 -116
rect -2447 -150 -2435 -116
rect -2493 -184 -2435 -150
rect -2493 -218 -2481 -184
rect -2447 -218 -2435 -184
rect -2493 -252 -2435 -218
rect -2493 -286 -2481 -252
rect -2447 -286 -2435 -252
rect -2493 -320 -2435 -286
rect -2493 -354 -2481 -320
rect -2447 -354 -2435 -320
rect -2493 -388 -2435 -354
rect -2493 -422 -2481 -388
rect -2447 -422 -2435 -388
rect -2493 -456 -2435 -422
rect -2493 -490 -2481 -456
rect -2447 -490 -2435 -456
rect -2493 -524 -2435 -490
rect -2493 -558 -2481 -524
rect -2447 -558 -2435 -524
rect -2493 -592 -2435 -558
rect -2493 -626 -2481 -592
rect -2447 -626 -2435 -592
rect -2493 -660 -2435 -626
rect -2493 -694 -2481 -660
rect -2447 -694 -2435 -660
rect -2493 -728 -2435 -694
rect -2493 -762 -2481 -728
rect -2447 -762 -2435 -728
rect -2493 -781 -2435 -762
rect -2185 700 -2127 719
rect -2185 666 -2173 700
rect -2139 666 -2127 700
rect -2185 632 -2127 666
rect -2185 598 -2173 632
rect -2139 598 -2127 632
rect -2185 564 -2127 598
rect -2185 530 -2173 564
rect -2139 530 -2127 564
rect -2185 496 -2127 530
rect -2185 462 -2173 496
rect -2139 462 -2127 496
rect -2185 428 -2127 462
rect -2185 394 -2173 428
rect -2139 394 -2127 428
rect -2185 360 -2127 394
rect -2185 326 -2173 360
rect -2139 326 -2127 360
rect -2185 292 -2127 326
rect -2185 258 -2173 292
rect -2139 258 -2127 292
rect -2185 224 -2127 258
rect -2185 190 -2173 224
rect -2139 190 -2127 224
rect -2185 156 -2127 190
rect -2185 122 -2173 156
rect -2139 122 -2127 156
rect -2185 88 -2127 122
rect -2185 54 -2173 88
rect -2139 54 -2127 88
rect -2185 20 -2127 54
rect -2185 -14 -2173 20
rect -2139 -14 -2127 20
rect -2185 -48 -2127 -14
rect -2185 -82 -2173 -48
rect -2139 -82 -2127 -48
rect -2185 -116 -2127 -82
rect -2185 -150 -2173 -116
rect -2139 -150 -2127 -116
rect -2185 -184 -2127 -150
rect -2185 -218 -2173 -184
rect -2139 -218 -2127 -184
rect -2185 -252 -2127 -218
rect -2185 -286 -2173 -252
rect -2139 -286 -2127 -252
rect -2185 -320 -2127 -286
rect -2185 -354 -2173 -320
rect -2139 -354 -2127 -320
rect -2185 -388 -2127 -354
rect -2185 -422 -2173 -388
rect -2139 -422 -2127 -388
rect -2185 -456 -2127 -422
rect -2185 -490 -2173 -456
rect -2139 -490 -2127 -456
rect -2185 -524 -2127 -490
rect -2185 -558 -2173 -524
rect -2139 -558 -2127 -524
rect -2185 -592 -2127 -558
rect -2185 -626 -2173 -592
rect -2139 -626 -2127 -592
rect -2185 -660 -2127 -626
rect -2185 -694 -2173 -660
rect -2139 -694 -2127 -660
rect -2185 -728 -2127 -694
rect -2185 -762 -2173 -728
rect -2139 -762 -2127 -728
rect -2185 -781 -2127 -762
rect -1877 700 -1819 719
rect -1877 666 -1865 700
rect -1831 666 -1819 700
rect -1877 632 -1819 666
rect -1877 598 -1865 632
rect -1831 598 -1819 632
rect -1877 564 -1819 598
rect -1877 530 -1865 564
rect -1831 530 -1819 564
rect -1877 496 -1819 530
rect -1877 462 -1865 496
rect -1831 462 -1819 496
rect -1877 428 -1819 462
rect -1877 394 -1865 428
rect -1831 394 -1819 428
rect -1877 360 -1819 394
rect -1877 326 -1865 360
rect -1831 326 -1819 360
rect -1877 292 -1819 326
rect -1877 258 -1865 292
rect -1831 258 -1819 292
rect -1877 224 -1819 258
rect -1877 190 -1865 224
rect -1831 190 -1819 224
rect -1877 156 -1819 190
rect -1877 122 -1865 156
rect -1831 122 -1819 156
rect -1877 88 -1819 122
rect -1877 54 -1865 88
rect -1831 54 -1819 88
rect -1877 20 -1819 54
rect -1877 -14 -1865 20
rect -1831 -14 -1819 20
rect -1877 -48 -1819 -14
rect -1877 -82 -1865 -48
rect -1831 -82 -1819 -48
rect -1877 -116 -1819 -82
rect -1877 -150 -1865 -116
rect -1831 -150 -1819 -116
rect -1877 -184 -1819 -150
rect -1877 -218 -1865 -184
rect -1831 -218 -1819 -184
rect -1877 -252 -1819 -218
rect -1877 -286 -1865 -252
rect -1831 -286 -1819 -252
rect -1877 -320 -1819 -286
rect -1877 -354 -1865 -320
rect -1831 -354 -1819 -320
rect -1877 -388 -1819 -354
rect -1877 -422 -1865 -388
rect -1831 -422 -1819 -388
rect -1877 -456 -1819 -422
rect -1877 -490 -1865 -456
rect -1831 -490 -1819 -456
rect -1877 -524 -1819 -490
rect -1877 -558 -1865 -524
rect -1831 -558 -1819 -524
rect -1877 -592 -1819 -558
rect -1877 -626 -1865 -592
rect -1831 -626 -1819 -592
rect -1877 -660 -1819 -626
rect -1877 -694 -1865 -660
rect -1831 -694 -1819 -660
rect -1877 -728 -1819 -694
rect -1877 -762 -1865 -728
rect -1831 -762 -1819 -728
rect -1877 -781 -1819 -762
rect -1569 700 -1511 719
rect -1569 666 -1557 700
rect -1523 666 -1511 700
rect -1569 632 -1511 666
rect -1569 598 -1557 632
rect -1523 598 -1511 632
rect -1569 564 -1511 598
rect -1569 530 -1557 564
rect -1523 530 -1511 564
rect -1569 496 -1511 530
rect -1569 462 -1557 496
rect -1523 462 -1511 496
rect -1569 428 -1511 462
rect -1569 394 -1557 428
rect -1523 394 -1511 428
rect -1569 360 -1511 394
rect -1569 326 -1557 360
rect -1523 326 -1511 360
rect -1569 292 -1511 326
rect -1569 258 -1557 292
rect -1523 258 -1511 292
rect -1569 224 -1511 258
rect -1569 190 -1557 224
rect -1523 190 -1511 224
rect -1569 156 -1511 190
rect -1569 122 -1557 156
rect -1523 122 -1511 156
rect -1569 88 -1511 122
rect -1569 54 -1557 88
rect -1523 54 -1511 88
rect -1569 20 -1511 54
rect -1569 -14 -1557 20
rect -1523 -14 -1511 20
rect -1569 -48 -1511 -14
rect -1569 -82 -1557 -48
rect -1523 -82 -1511 -48
rect -1569 -116 -1511 -82
rect -1569 -150 -1557 -116
rect -1523 -150 -1511 -116
rect -1569 -184 -1511 -150
rect -1569 -218 -1557 -184
rect -1523 -218 -1511 -184
rect -1569 -252 -1511 -218
rect -1569 -286 -1557 -252
rect -1523 -286 -1511 -252
rect -1569 -320 -1511 -286
rect -1569 -354 -1557 -320
rect -1523 -354 -1511 -320
rect -1569 -388 -1511 -354
rect -1569 -422 -1557 -388
rect -1523 -422 -1511 -388
rect -1569 -456 -1511 -422
rect -1569 -490 -1557 -456
rect -1523 -490 -1511 -456
rect -1569 -524 -1511 -490
rect -1569 -558 -1557 -524
rect -1523 -558 -1511 -524
rect -1569 -592 -1511 -558
rect -1569 -626 -1557 -592
rect -1523 -626 -1511 -592
rect -1569 -660 -1511 -626
rect -1569 -694 -1557 -660
rect -1523 -694 -1511 -660
rect -1569 -728 -1511 -694
rect -1569 -762 -1557 -728
rect -1523 -762 -1511 -728
rect -1569 -781 -1511 -762
rect -1261 700 -1203 719
rect -1261 666 -1249 700
rect -1215 666 -1203 700
rect -1261 632 -1203 666
rect -1261 598 -1249 632
rect -1215 598 -1203 632
rect -1261 564 -1203 598
rect -1261 530 -1249 564
rect -1215 530 -1203 564
rect -1261 496 -1203 530
rect -1261 462 -1249 496
rect -1215 462 -1203 496
rect -1261 428 -1203 462
rect -1261 394 -1249 428
rect -1215 394 -1203 428
rect -1261 360 -1203 394
rect -1261 326 -1249 360
rect -1215 326 -1203 360
rect -1261 292 -1203 326
rect -1261 258 -1249 292
rect -1215 258 -1203 292
rect -1261 224 -1203 258
rect -1261 190 -1249 224
rect -1215 190 -1203 224
rect -1261 156 -1203 190
rect -1261 122 -1249 156
rect -1215 122 -1203 156
rect -1261 88 -1203 122
rect -1261 54 -1249 88
rect -1215 54 -1203 88
rect -1261 20 -1203 54
rect -1261 -14 -1249 20
rect -1215 -14 -1203 20
rect -1261 -48 -1203 -14
rect -1261 -82 -1249 -48
rect -1215 -82 -1203 -48
rect -1261 -116 -1203 -82
rect -1261 -150 -1249 -116
rect -1215 -150 -1203 -116
rect -1261 -184 -1203 -150
rect -1261 -218 -1249 -184
rect -1215 -218 -1203 -184
rect -1261 -252 -1203 -218
rect -1261 -286 -1249 -252
rect -1215 -286 -1203 -252
rect -1261 -320 -1203 -286
rect -1261 -354 -1249 -320
rect -1215 -354 -1203 -320
rect -1261 -388 -1203 -354
rect -1261 -422 -1249 -388
rect -1215 -422 -1203 -388
rect -1261 -456 -1203 -422
rect -1261 -490 -1249 -456
rect -1215 -490 -1203 -456
rect -1261 -524 -1203 -490
rect -1261 -558 -1249 -524
rect -1215 -558 -1203 -524
rect -1261 -592 -1203 -558
rect -1261 -626 -1249 -592
rect -1215 -626 -1203 -592
rect -1261 -660 -1203 -626
rect -1261 -694 -1249 -660
rect -1215 -694 -1203 -660
rect -1261 -728 -1203 -694
rect -1261 -762 -1249 -728
rect -1215 -762 -1203 -728
rect -1261 -781 -1203 -762
rect -953 700 -895 719
rect -953 666 -941 700
rect -907 666 -895 700
rect -953 632 -895 666
rect -953 598 -941 632
rect -907 598 -895 632
rect -953 564 -895 598
rect -953 530 -941 564
rect -907 530 -895 564
rect -953 496 -895 530
rect -953 462 -941 496
rect -907 462 -895 496
rect -953 428 -895 462
rect -953 394 -941 428
rect -907 394 -895 428
rect -953 360 -895 394
rect -953 326 -941 360
rect -907 326 -895 360
rect -953 292 -895 326
rect -953 258 -941 292
rect -907 258 -895 292
rect -953 224 -895 258
rect -953 190 -941 224
rect -907 190 -895 224
rect -953 156 -895 190
rect -953 122 -941 156
rect -907 122 -895 156
rect -953 88 -895 122
rect -953 54 -941 88
rect -907 54 -895 88
rect -953 20 -895 54
rect -953 -14 -941 20
rect -907 -14 -895 20
rect -953 -48 -895 -14
rect -953 -82 -941 -48
rect -907 -82 -895 -48
rect -953 -116 -895 -82
rect -953 -150 -941 -116
rect -907 -150 -895 -116
rect -953 -184 -895 -150
rect -953 -218 -941 -184
rect -907 -218 -895 -184
rect -953 -252 -895 -218
rect -953 -286 -941 -252
rect -907 -286 -895 -252
rect -953 -320 -895 -286
rect -953 -354 -941 -320
rect -907 -354 -895 -320
rect -953 -388 -895 -354
rect -953 -422 -941 -388
rect -907 -422 -895 -388
rect -953 -456 -895 -422
rect -953 -490 -941 -456
rect -907 -490 -895 -456
rect -953 -524 -895 -490
rect -953 -558 -941 -524
rect -907 -558 -895 -524
rect -953 -592 -895 -558
rect -953 -626 -941 -592
rect -907 -626 -895 -592
rect -953 -660 -895 -626
rect -953 -694 -941 -660
rect -907 -694 -895 -660
rect -953 -728 -895 -694
rect -953 -762 -941 -728
rect -907 -762 -895 -728
rect -953 -781 -895 -762
rect -645 700 -587 719
rect -645 666 -633 700
rect -599 666 -587 700
rect -645 632 -587 666
rect -645 598 -633 632
rect -599 598 -587 632
rect -645 564 -587 598
rect -645 530 -633 564
rect -599 530 -587 564
rect -645 496 -587 530
rect -645 462 -633 496
rect -599 462 -587 496
rect -645 428 -587 462
rect -645 394 -633 428
rect -599 394 -587 428
rect -645 360 -587 394
rect -645 326 -633 360
rect -599 326 -587 360
rect -645 292 -587 326
rect -645 258 -633 292
rect -599 258 -587 292
rect -645 224 -587 258
rect -645 190 -633 224
rect -599 190 -587 224
rect -645 156 -587 190
rect -645 122 -633 156
rect -599 122 -587 156
rect -645 88 -587 122
rect -645 54 -633 88
rect -599 54 -587 88
rect -645 20 -587 54
rect -645 -14 -633 20
rect -599 -14 -587 20
rect -645 -48 -587 -14
rect -645 -82 -633 -48
rect -599 -82 -587 -48
rect -645 -116 -587 -82
rect -645 -150 -633 -116
rect -599 -150 -587 -116
rect -645 -184 -587 -150
rect -645 -218 -633 -184
rect -599 -218 -587 -184
rect -645 -252 -587 -218
rect -645 -286 -633 -252
rect -599 -286 -587 -252
rect -645 -320 -587 -286
rect -645 -354 -633 -320
rect -599 -354 -587 -320
rect -645 -388 -587 -354
rect -645 -422 -633 -388
rect -599 -422 -587 -388
rect -645 -456 -587 -422
rect -645 -490 -633 -456
rect -599 -490 -587 -456
rect -645 -524 -587 -490
rect -645 -558 -633 -524
rect -599 -558 -587 -524
rect -645 -592 -587 -558
rect -645 -626 -633 -592
rect -599 -626 -587 -592
rect -645 -660 -587 -626
rect -645 -694 -633 -660
rect -599 -694 -587 -660
rect -645 -728 -587 -694
rect -645 -762 -633 -728
rect -599 -762 -587 -728
rect -645 -781 -587 -762
rect -337 700 -279 719
rect -337 666 -325 700
rect -291 666 -279 700
rect -337 632 -279 666
rect -337 598 -325 632
rect -291 598 -279 632
rect -337 564 -279 598
rect -337 530 -325 564
rect -291 530 -279 564
rect -337 496 -279 530
rect -337 462 -325 496
rect -291 462 -279 496
rect -337 428 -279 462
rect -337 394 -325 428
rect -291 394 -279 428
rect -337 360 -279 394
rect -337 326 -325 360
rect -291 326 -279 360
rect -337 292 -279 326
rect -337 258 -325 292
rect -291 258 -279 292
rect -337 224 -279 258
rect -337 190 -325 224
rect -291 190 -279 224
rect -337 156 -279 190
rect -337 122 -325 156
rect -291 122 -279 156
rect -337 88 -279 122
rect -337 54 -325 88
rect -291 54 -279 88
rect -337 20 -279 54
rect -337 -14 -325 20
rect -291 -14 -279 20
rect -337 -48 -279 -14
rect -337 -82 -325 -48
rect -291 -82 -279 -48
rect -337 -116 -279 -82
rect -337 -150 -325 -116
rect -291 -150 -279 -116
rect -337 -184 -279 -150
rect -337 -218 -325 -184
rect -291 -218 -279 -184
rect -337 -252 -279 -218
rect -337 -286 -325 -252
rect -291 -286 -279 -252
rect -337 -320 -279 -286
rect -337 -354 -325 -320
rect -291 -354 -279 -320
rect -337 -388 -279 -354
rect -337 -422 -325 -388
rect -291 -422 -279 -388
rect -337 -456 -279 -422
rect -337 -490 -325 -456
rect -291 -490 -279 -456
rect -337 -524 -279 -490
rect -337 -558 -325 -524
rect -291 -558 -279 -524
rect -337 -592 -279 -558
rect -337 -626 -325 -592
rect -291 -626 -279 -592
rect -337 -660 -279 -626
rect -337 -694 -325 -660
rect -291 -694 -279 -660
rect -337 -728 -279 -694
rect -337 -762 -325 -728
rect -291 -762 -279 -728
rect -337 -781 -279 -762
rect -29 700 29 719
rect -29 666 -17 700
rect 17 666 29 700
rect -29 632 29 666
rect -29 598 -17 632
rect 17 598 29 632
rect -29 564 29 598
rect -29 530 -17 564
rect 17 530 29 564
rect -29 496 29 530
rect -29 462 -17 496
rect 17 462 29 496
rect -29 428 29 462
rect -29 394 -17 428
rect 17 394 29 428
rect -29 360 29 394
rect -29 326 -17 360
rect 17 326 29 360
rect -29 292 29 326
rect -29 258 -17 292
rect 17 258 29 292
rect -29 224 29 258
rect -29 190 -17 224
rect 17 190 29 224
rect -29 156 29 190
rect -29 122 -17 156
rect 17 122 29 156
rect -29 88 29 122
rect -29 54 -17 88
rect 17 54 29 88
rect -29 20 29 54
rect -29 -14 -17 20
rect 17 -14 29 20
rect -29 -48 29 -14
rect -29 -82 -17 -48
rect 17 -82 29 -48
rect -29 -116 29 -82
rect -29 -150 -17 -116
rect 17 -150 29 -116
rect -29 -184 29 -150
rect -29 -218 -17 -184
rect 17 -218 29 -184
rect -29 -252 29 -218
rect -29 -286 -17 -252
rect 17 -286 29 -252
rect -29 -320 29 -286
rect -29 -354 -17 -320
rect 17 -354 29 -320
rect -29 -388 29 -354
rect -29 -422 -17 -388
rect 17 -422 29 -388
rect -29 -456 29 -422
rect -29 -490 -17 -456
rect 17 -490 29 -456
rect -29 -524 29 -490
rect -29 -558 -17 -524
rect 17 -558 29 -524
rect -29 -592 29 -558
rect -29 -626 -17 -592
rect 17 -626 29 -592
rect -29 -660 29 -626
rect -29 -694 -17 -660
rect 17 -694 29 -660
rect -29 -728 29 -694
rect -29 -762 -17 -728
rect 17 -762 29 -728
rect -29 -781 29 -762
rect 279 700 337 719
rect 279 666 291 700
rect 325 666 337 700
rect 279 632 337 666
rect 279 598 291 632
rect 325 598 337 632
rect 279 564 337 598
rect 279 530 291 564
rect 325 530 337 564
rect 279 496 337 530
rect 279 462 291 496
rect 325 462 337 496
rect 279 428 337 462
rect 279 394 291 428
rect 325 394 337 428
rect 279 360 337 394
rect 279 326 291 360
rect 325 326 337 360
rect 279 292 337 326
rect 279 258 291 292
rect 325 258 337 292
rect 279 224 337 258
rect 279 190 291 224
rect 325 190 337 224
rect 279 156 337 190
rect 279 122 291 156
rect 325 122 337 156
rect 279 88 337 122
rect 279 54 291 88
rect 325 54 337 88
rect 279 20 337 54
rect 279 -14 291 20
rect 325 -14 337 20
rect 279 -48 337 -14
rect 279 -82 291 -48
rect 325 -82 337 -48
rect 279 -116 337 -82
rect 279 -150 291 -116
rect 325 -150 337 -116
rect 279 -184 337 -150
rect 279 -218 291 -184
rect 325 -218 337 -184
rect 279 -252 337 -218
rect 279 -286 291 -252
rect 325 -286 337 -252
rect 279 -320 337 -286
rect 279 -354 291 -320
rect 325 -354 337 -320
rect 279 -388 337 -354
rect 279 -422 291 -388
rect 325 -422 337 -388
rect 279 -456 337 -422
rect 279 -490 291 -456
rect 325 -490 337 -456
rect 279 -524 337 -490
rect 279 -558 291 -524
rect 325 -558 337 -524
rect 279 -592 337 -558
rect 279 -626 291 -592
rect 325 -626 337 -592
rect 279 -660 337 -626
rect 279 -694 291 -660
rect 325 -694 337 -660
rect 279 -728 337 -694
rect 279 -762 291 -728
rect 325 -762 337 -728
rect 279 -781 337 -762
rect 587 700 645 719
rect 587 666 599 700
rect 633 666 645 700
rect 587 632 645 666
rect 587 598 599 632
rect 633 598 645 632
rect 587 564 645 598
rect 587 530 599 564
rect 633 530 645 564
rect 587 496 645 530
rect 587 462 599 496
rect 633 462 645 496
rect 587 428 645 462
rect 587 394 599 428
rect 633 394 645 428
rect 587 360 645 394
rect 587 326 599 360
rect 633 326 645 360
rect 587 292 645 326
rect 587 258 599 292
rect 633 258 645 292
rect 587 224 645 258
rect 587 190 599 224
rect 633 190 645 224
rect 587 156 645 190
rect 587 122 599 156
rect 633 122 645 156
rect 587 88 645 122
rect 587 54 599 88
rect 633 54 645 88
rect 587 20 645 54
rect 587 -14 599 20
rect 633 -14 645 20
rect 587 -48 645 -14
rect 587 -82 599 -48
rect 633 -82 645 -48
rect 587 -116 645 -82
rect 587 -150 599 -116
rect 633 -150 645 -116
rect 587 -184 645 -150
rect 587 -218 599 -184
rect 633 -218 645 -184
rect 587 -252 645 -218
rect 587 -286 599 -252
rect 633 -286 645 -252
rect 587 -320 645 -286
rect 587 -354 599 -320
rect 633 -354 645 -320
rect 587 -388 645 -354
rect 587 -422 599 -388
rect 633 -422 645 -388
rect 587 -456 645 -422
rect 587 -490 599 -456
rect 633 -490 645 -456
rect 587 -524 645 -490
rect 587 -558 599 -524
rect 633 -558 645 -524
rect 587 -592 645 -558
rect 587 -626 599 -592
rect 633 -626 645 -592
rect 587 -660 645 -626
rect 587 -694 599 -660
rect 633 -694 645 -660
rect 587 -728 645 -694
rect 587 -762 599 -728
rect 633 -762 645 -728
rect 587 -781 645 -762
rect 895 700 953 719
rect 895 666 907 700
rect 941 666 953 700
rect 895 632 953 666
rect 895 598 907 632
rect 941 598 953 632
rect 895 564 953 598
rect 895 530 907 564
rect 941 530 953 564
rect 895 496 953 530
rect 895 462 907 496
rect 941 462 953 496
rect 895 428 953 462
rect 895 394 907 428
rect 941 394 953 428
rect 895 360 953 394
rect 895 326 907 360
rect 941 326 953 360
rect 895 292 953 326
rect 895 258 907 292
rect 941 258 953 292
rect 895 224 953 258
rect 895 190 907 224
rect 941 190 953 224
rect 895 156 953 190
rect 895 122 907 156
rect 941 122 953 156
rect 895 88 953 122
rect 895 54 907 88
rect 941 54 953 88
rect 895 20 953 54
rect 895 -14 907 20
rect 941 -14 953 20
rect 895 -48 953 -14
rect 895 -82 907 -48
rect 941 -82 953 -48
rect 895 -116 953 -82
rect 895 -150 907 -116
rect 941 -150 953 -116
rect 895 -184 953 -150
rect 895 -218 907 -184
rect 941 -218 953 -184
rect 895 -252 953 -218
rect 895 -286 907 -252
rect 941 -286 953 -252
rect 895 -320 953 -286
rect 895 -354 907 -320
rect 941 -354 953 -320
rect 895 -388 953 -354
rect 895 -422 907 -388
rect 941 -422 953 -388
rect 895 -456 953 -422
rect 895 -490 907 -456
rect 941 -490 953 -456
rect 895 -524 953 -490
rect 895 -558 907 -524
rect 941 -558 953 -524
rect 895 -592 953 -558
rect 895 -626 907 -592
rect 941 -626 953 -592
rect 895 -660 953 -626
rect 895 -694 907 -660
rect 941 -694 953 -660
rect 895 -728 953 -694
rect 895 -762 907 -728
rect 941 -762 953 -728
rect 895 -781 953 -762
rect 1203 700 1261 719
rect 1203 666 1215 700
rect 1249 666 1261 700
rect 1203 632 1261 666
rect 1203 598 1215 632
rect 1249 598 1261 632
rect 1203 564 1261 598
rect 1203 530 1215 564
rect 1249 530 1261 564
rect 1203 496 1261 530
rect 1203 462 1215 496
rect 1249 462 1261 496
rect 1203 428 1261 462
rect 1203 394 1215 428
rect 1249 394 1261 428
rect 1203 360 1261 394
rect 1203 326 1215 360
rect 1249 326 1261 360
rect 1203 292 1261 326
rect 1203 258 1215 292
rect 1249 258 1261 292
rect 1203 224 1261 258
rect 1203 190 1215 224
rect 1249 190 1261 224
rect 1203 156 1261 190
rect 1203 122 1215 156
rect 1249 122 1261 156
rect 1203 88 1261 122
rect 1203 54 1215 88
rect 1249 54 1261 88
rect 1203 20 1261 54
rect 1203 -14 1215 20
rect 1249 -14 1261 20
rect 1203 -48 1261 -14
rect 1203 -82 1215 -48
rect 1249 -82 1261 -48
rect 1203 -116 1261 -82
rect 1203 -150 1215 -116
rect 1249 -150 1261 -116
rect 1203 -184 1261 -150
rect 1203 -218 1215 -184
rect 1249 -218 1261 -184
rect 1203 -252 1261 -218
rect 1203 -286 1215 -252
rect 1249 -286 1261 -252
rect 1203 -320 1261 -286
rect 1203 -354 1215 -320
rect 1249 -354 1261 -320
rect 1203 -388 1261 -354
rect 1203 -422 1215 -388
rect 1249 -422 1261 -388
rect 1203 -456 1261 -422
rect 1203 -490 1215 -456
rect 1249 -490 1261 -456
rect 1203 -524 1261 -490
rect 1203 -558 1215 -524
rect 1249 -558 1261 -524
rect 1203 -592 1261 -558
rect 1203 -626 1215 -592
rect 1249 -626 1261 -592
rect 1203 -660 1261 -626
rect 1203 -694 1215 -660
rect 1249 -694 1261 -660
rect 1203 -728 1261 -694
rect 1203 -762 1215 -728
rect 1249 -762 1261 -728
rect 1203 -781 1261 -762
rect 1511 700 1569 719
rect 1511 666 1523 700
rect 1557 666 1569 700
rect 1511 632 1569 666
rect 1511 598 1523 632
rect 1557 598 1569 632
rect 1511 564 1569 598
rect 1511 530 1523 564
rect 1557 530 1569 564
rect 1511 496 1569 530
rect 1511 462 1523 496
rect 1557 462 1569 496
rect 1511 428 1569 462
rect 1511 394 1523 428
rect 1557 394 1569 428
rect 1511 360 1569 394
rect 1511 326 1523 360
rect 1557 326 1569 360
rect 1511 292 1569 326
rect 1511 258 1523 292
rect 1557 258 1569 292
rect 1511 224 1569 258
rect 1511 190 1523 224
rect 1557 190 1569 224
rect 1511 156 1569 190
rect 1511 122 1523 156
rect 1557 122 1569 156
rect 1511 88 1569 122
rect 1511 54 1523 88
rect 1557 54 1569 88
rect 1511 20 1569 54
rect 1511 -14 1523 20
rect 1557 -14 1569 20
rect 1511 -48 1569 -14
rect 1511 -82 1523 -48
rect 1557 -82 1569 -48
rect 1511 -116 1569 -82
rect 1511 -150 1523 -116
rect 1557 -150 1569 -116
rect 1511 -184 1569 -150
rect 1511 -218 1523 -184
rect 1557 -218 1569 -184
rect 1511 -252 1569 -218
rect 1511 -286 1523 -252
rect 1557 -286 1569 -252
rect 1511 -320 1569 -286
rect 1511 -354 1523 -320
rect 1557 -354 1569 -320
rect 1511 -388 1569 -354
rect 1511 -422 1523 -388
rect 1557 -422 1569 -388
rect 1511 -456 1569 -422
rect 1511 -490 1523 -456
rect 1557 -490 1569 -456
rect 1511 -524 1569 -490
rect 1511 -558 1523 -524
rect 1557 -558 1569 -524
rect 1511 -592 1569 -558
rect 1511 -626 1523 -592
rect 1557 -626 1569 -592
rect 1511 -660 1569 -626
rect 1511 -694 1523 -660
rect 1557 -694 1569 -660
rect 1511 -728 1569 -694
rect 1511 -762 1523 -728
rect 1557 -762 1569 -728
rect 1511 -781 1569 -762
rect 1819 700 1877 719
rect 1819 666 1831 700
rect 1865 666 1877 700
rect 1819 632 1877 666
rect 1819 598 1831 632
rect 1865 598 1877 632
rect 1819 564 1877 598
rect 1819 530 1831 564
rect 1865 530 1877 564
rect 1819 496 1877 530
rect 1819 462 1831 496
rect 1865 462 1877 496
rect 1819 428 1877 462
rect 1819 394 1831 428
rect 1865 394 1877 428
rect 1819 360 1877 394
rect 1819 326 1831 360
rect 1865 326 1877 360
rect 1819 292 1877 326
rect 1819 258 1831 292
rect 1865 258 1877 292
rect 1819 224 1877 258
rect 1819 190 1831 224
rect 1865 190 1877 224
rect 1819 156 1877 190
rect 1819 122 1831 156
rect 1865 122 1877 156
rect 1819 88 1877 122
rect 1819 54 1831 88
rect 1865 54 1877 88
rect 1819 20 1877 54
rect 1819 -14 1831 20
rect 1865 -14 1877 20
rect 1819 -48 1877 -14
rect 1819 -82 1831 -48
rect 1865 -82 1877 -48
rect 1819 -116 1877 -82
rect 1819 -150 1831 -116
rect 1865 -150 1877 -116
rect 1819 -184 1877 -150
rect 1819 -218 1831 -184
rect 1865 -218 1877 -184
rect 1819 -252 1877 -218
rect 1819 -286 1831 -252
rect 1865 -286 1877 -252
rect 1819 -320 1877 -286
rect 1819 -354 1831 -320
rect 1865 -354 1877 -320
rect 1819 -388 1877 -354
rect 1819 -422 1831 -388
rect 1865 -422 1877 -388
rect 1819 -456 1877 -422
rect 1819 -490 1831 -456
rect 1865 -490 1877 -456
rect 1819 -524 1877 -490
rect 1819 -558 1831 -524
rect 1865 -558 1877 -524
rect 1819 -592 1877 -558
rect 1819 -626 1831 -592
rect 1865 -626 1877 -592
rect 1819 -660 1877 -626
rect 1819 -694 1831 -660
rect 1865 -694 1877 -660
rect 1819 -728 1877 -694
rect 1819 -762 1831 -728
rect 1865 -762 1877 -728
rect 1819 -781 1877 -762
rect 2127 700 2185 719
rect 2127 666 2139 700
rect 2173 666 2185 700
rect 2127 632 2185 666
rect 2127 598 2139 632
rect 2173 598 2185 632
rect 2127 564 2185 598
rect 2127 530 2139 564
rect 2173 530 2185 564
rect 2127 496 2185 530
rect 2127 462 2139 496
rect 2173 462 2185 496
rect 2127 428 2185 462
rect 2127 394 2139 428
rect 2173 394 2185 428
rect 2127 360 2185 394
rect 2127 326 2139 360
rect 2173 326 2185 360
rect 2127 292 2185 326
rect 2127 258 2139 292
rect 2173 258 2185 292
rect 2127 224 2185 258
rect 2127 190 2139 224
rect 2173 190 2185 224
rect 2127 156 2185 190
rect 2127 122 2139 156
rect 2173 122 2185 156
rect 2127 88 2185 122
rect 2127 54 2139 88
rect 2173 54 2185 88
rect 2127 20 2185 54
rect 2127 -14 2139 20
rect 2173 -14 2185 20
rect 2127 -48 2185 -14
rect 2127 -82 2139 -48
rect 2173 -82 2185 -48
rect 2127 -116 2185 -82
rect 2127 -150 2139 -116
rect 2173 -150 2185 -116
rect 2127 -184 2185 -150
rect 2127 -218 2139 -184
rect 2173 -218 2185 -184
rect 2127 -252 2185 -218
rect 2127 -286 2139 -252
rect 2173 -286 2185 -252
rect 2127 -320 2185 -286
rect 2127 -354 2139 -320
rect 2173 -354 2185 -320
rect 2127 -388 2185 -354
rect 2127 -422 2139 -388
rect 2173 -422 2185 -388
rect 2127 -456 2185 -422
rect 2127 -490 2139 -456
rect 2173 -490 2185 -456
rect 2127 -524 2185 -490
rect 2127 -558 2139 -524
rect 2173 -558 2185 -524
rect 2127 -592 2185 -558
rect 2127 -626 2139 -592
rect 2173 -626 2185 -592
rect 2127 -660 2185 -626
rect 2127 -694 2139 -660
rect 2173 -694 2185 -660
rect 2127 -728 2185 -694
rect 2127 -762 2139 -728
rect 2173 -762 2185 -728
rect 2127 -781 2185 -762
rect 2435 700 2493 719
rect 2435 666 2447 700
rect 2481 666 2493 700
rect 2435 632 2493 666
rect 2435 598 2447 632
rect 2481 598 2493 632
rect 2435 564 2493 598
rect 2435 530 2447 564
rect 2481 530 2493 564
rect 2435 496 2493 530
rect 2435 462 2447 496
rect 2481 462 2493 496
rect 2435 428 2493 462
rect 2435 394 2447 428
rect 2481 394 2493 428
rect 2435 360 2493 394
rect 2435 326 2447 360
rect 2481 326 2493 360
rect 2435 292 2493 326
rect 2435 258 2447 292
rect 2481 258 2493 292
rect 2435 224 2493 258
rect 2435 190 2447 224
rect 2481 190 2493 224
rect 2435 156 2493 190
rect 2435 122 2447 156
rect 2481 122 2493 156
rect 2435 88 2493 122
rect 2435 54 2447 88
rect 2481 54 2493 88
rect 2435 20 2493 54
rect 2435 -14 2447 20
rect 2481 -14 2493 20
rect 2435 -48 2493 -14
rect 2435 -82 2447 -48
rect 2481 -82 2493 -48
rect 2435 -116 2493 -82
rect 2435 -150 2447 -116
rect 2481 -150 2493 -116
rect 2435 -184 2493 -150
rect 2435 -218 2447 -184
rect 2481 -218 2493 -184
rect 2435 -252 2493 -218
rect 2435 -286 2447 -252
rect 2481 -286 2493 -252
rect 2435 -320 2493 -286
rect 2435 -354 2447 -320
rect 2481 -354 2493 -320
rect 2435 -388 2493 -354
rect 2435 -422 2447 -388
rect 2481 -422 2493 -388
rect 2435 -456 2493 -422
rect 2435 -490 2447 -456
rect 2481 -490 2493 -456
rect 2435 -524 2493 -490
rect 2435 -558 2447 -524
rect 2481 -558 2493 -524
rect 2435 -592 2493 -558
rect 2435 -626 2447 -592
rect 2481 -626 2493 -592
rect 2435 -660 2493 -626
rect 2435 -694 2447 -660
rect 2481 -694 2493 -660
rect 2435 -728 2493 -694
rect 2435 -762 2447 -728
rect 2481 -762 2493 -728
rect 2435 -781 2493 -762
rect 2743 700 2801 719
rect 2743 666 2755 700
rect 2789 666 2801 700
rect 2743 632 2801 666
rect 2743 598 2755 632
rect 2789 598 2801 632
rect 2743 564 2801 598
rect 2743 530 2755 564
rect 2789 530 2801 564
rect 2743 496 2801 530
rect 2743 462 2755 496
rect 2789 462 2801 496
rect 2743 428 2801 462
rect 2743 394 2755 428
rect 2789 394 2801 428
rect 2743 360 2801 394
rect 2743 326 2755 360
rect 2789 326 2801 360
rect 2743 292 2801 326
rect 2743 258 2755 292
rect 2789 258 2801 292
rect 2743 224 2801 258
rect 2743 190 2755 224
rect 2789 190 2801 224
rect 2743 156 2801 190
rect 2743 122 2755 156
rect 2789 122 2801 156
rect 2743 88 2801 122
rect 2743 54 2755 88
rect 2789 54 2801 88
rect 2743 20 2801 54
rect 2743 -14 2755 20
rect 2789 -14 2801 20
rect 2743 -48 2801 -14
rect 2743 -82 2755 -48
rect 2789 -82 2801 -48
rect 2743 -116 2801 -82
rect 2743 -150 2755 -116
rect 2789 -150 2801 -116
rect 2743 -184 2801 -150
rect 2743 -218 2755 -184
rect 2789 -218 2801 -184
rect 2743 -252 2801 -218
rect 2743 -286 2755 -252
rect 2789 -286 2801 -252
rect 2743 -320 2801 -286
rect 2743 -354 2755 -320
rect 2789 -354 2801 -320
rect 2743 -388 2801 -354
rect 2743 -422 2755 -388
rect 2789 -422 2801 -388
rect 2743 -456 2801 -422
rect 2743 -490 2755 -456
rect 2789 -490 2801 -456
rect 2743 -524 2801 -490
rect 2743 -558 2755 -524
rect 2789 -558 2801 -524
rect 2743 -592 2801 -558
rect 2743 -626 2755 -592
rect 2789 -626 2801 -592
rect 2743 -660 2801 -626
rect 2743 -694 2755 -660
rect 2789 -694 2801 -660
rect 2743 -728 2801 -694
rect 2743 -762 2755 -728
rect 2789 -762 2801 -728
rect 2743 -781 2801 -762
<< mvndiffc >>
rect -2789 666 -2755 700
rect -2789 598 -2755 632
rect -2789 530 -2755 564
rect -2789 462 -2755 496
rect -2789 394 -2755 428
rect -2789 326 -2755 360
rect -2789 258 -2755 292
rect -2789 190 -2755 224
rect -2789 122 -2755 156
rect -2789 54 -2755 88
rect -2789 -14 -2755 20
rect -2789 -82 -2755 -48
rect -2789 -150 -2755 -116
rect -2789 -218 -2755 -184
rect -2789 -286 -2755 -252
rect -2789 -354 -2755 -320
rect -2789 -422 -2755 -388
rect -2789 -490 -2755 -456
rect -2789 -558 -2755 -524
rect -2789 -626 -2755 -592
rect -2789 -694 -2755 -660
rect -2789 -762 -2755 -728
rect -2481 666 -2447 700
rect -2481 598 -2447 632
rect -2481 530 -2447 564
rect -2481 462 -2447 496
rect -2481 394 -2447 428
rect -2481 326 -2447 360
rect -2481 258 -2447 292
rect -2481 190 -2447 224
rect -2481 122 -2447 156
rect -2481 54 -2447 88
rect -2481 -14 -2447 20
rect -2481 -82 -2447 -48
rect -2481 -150 -2447 -116
rect -2481 -218 -2447 -184
rect -2481 -286 -2447 -252
rect -2481 -354 -2447 -320
rect -2481 -422 -2447 -388
rect -2481 -490 -2447 -456
rect -2481 -558 -2447 -524
rect -2481 -626 -2447 -592
rect -2481 -694 -2447 -660
rect -2481 -762 -2447 -728
rect -2173 666 -2139 700
rect -2173 598 -2139 632
rect -2173 530 -2139 564
rect -2173 462 -2139 496
rect -2173 394 -2139 428
rect -2173 326 -2139 360
rect -2173 258 -2139 292
rect -2173 190 -2139 224
rect -2173 122 -2139 156
rect -2173 54 -2139 88
rect -2173 -14 -2139 20
rect -2173 -82 -2139 -48
rect -2173 -150 -2139 -116
rect -2173 -218 -2139 -184
rect -2173 -286 -2139 -252
rect -2173 -354 -2139 -320
rect -2173 -422 -2139 -388
rect -2173 -490 -2139 -456
rect -2173 -558 -2139 -524
rect -2173 -626 -2139 -592
rect -2173 -694 -2139 -660
rect -2173 -762 -2139 -728
rect -1865 666 -1831 700
rect -1865 598 -1831 632
rect -1865 530 -1831 564
rect -1865 462 -1831 496
rect -1865 394 -1831 428
rect -1865 326 -1831 360
rect -1865 258 -1831 292
rect -1865 190 -1831 224
rect -1865 122 -1831 156
rect -1865 54 -1831 88
rect -1865 -14 -1831 20
rect -1865 -82 -1831 -48
rect -1865 -150 -1831 -116
rect -1865 -218 -1831 -184
rect -1865 -286 -1831 -252
rect -1865 -354 -1831 -320
rect -1865 -422 -1831 -388
rect -1865 -490 -1831 -456
rect -1865 -558 -1831 -524
rect -1865 -626 -1831 -592
rect -1865 -694 -1831 -660
rect -1865 -762 -1831 -728
rect -1557 666 -1523 700
rect -1557 598 -1523 632
rect -1557 530 -1523 564
rect -1557 462 -1523 496
rect -1557 394 -1523 428
rect -1557 326 -1523 360
rect -1557 258 -1523 292
rect -1557 190 -1523 224
rect -1557 122 -1523 156
rect -1557 54 -1523 88
rect -1557 -14 -1523 20
rect -1557 -82 -1523 -48
rect -1557 -150 -1523 -116
rect -1557 -218 -1523 -184
rect -1557 -286 -1523 -252
rect -1557 -354 -1523 -320
rect -1557 -422 -1523 -388
rect -1557 -490 -1523 -456
rect -1557 -558 -1523 -524
rect -1557 -626 -1523 -592
rect -1557 -694 -1523 -660
rect -1557 -762 -1523 -728
rect -1249 666 -1215 700
rect -1249 598 -1215 632
rect -1249 530 -1215 564
rect -1249 462 -1215 496
rect -1249 394 -1215 428
rect -1249 326 -1215 360
rect -1249 258 -1215 292
rect -1249 190 -1215 224
rect -1249 122 -1215 156
rect -1249 54 -1215 88
rect -1249 -14 -1215 20
rect -1249 -82 -1215 -48
rect -1249 -150 -1215 -116
rect -1249 -218 -1215 -184
rect -1249 -286 -1215 -252
rect -1249 -354 -1215 -320
rect -1249 -422 -1215 -388
rect -1249 -490 -1215 -456
rect -1249 -558 -1215 -524
rect -1249 -626 -1215 -592
rect -1249 -694 -1215 -660
rect -1249 -762 -1215 -728
rect -941 666 -907 700
rect -941 598 -907 632
rect -941 530 -907 564
rect -941 462 -907 496
rect -941 394 -907 428
rect -941 326 -907 360
rect -941 258 -907 292
rect -941 190 -907 224
rect -941 122 -907 156
rect -941 54 -907 88
rect -941 -14 -907 20
rect -941 -82 -907 -48
rect -941 -150 -907 -116
rect -941 -218 -907 -184
rect -941 -286 -907 -252
rect -941 -354 -907 -320
rect -941 -422 -907 -388
rect -941 -490 -907 -456
rect -941 -558 -907 -524
rect -941 -626 -907 -592
rect -941 -694 -907 -660
rect -941 -762 -907 -728
rect -633 666 -599 700
rect -633 598 -599 632
rect -633 530 -599 564
rect -633 462 -599 496
rect -633 394 -599 428
rect -633 326 -599 360
rect -633 258 -599 292
rect -633 190 -599 224
rect -633 122 -599 156
rect -633 54 -599 88
rect -633 -14 -599 20
rect -633 -82 -599 -48
rect -633 -150 -599 -116
rect -633 -218 -599 -184
rect -633 -286 -599 -252
rect -633 -354 -599 -320
rect -633 -422 -599 -388
rect -633 -490 -599 -456
rect -633 -558 -599 -524
rect -633 -626 -599 -592
rect -633 -694 -599 -660
rect -633 -762 -599 -728
rect -325 666 -291 700
rect -325 598 -291 632
rect -325 530 -291 564
rect -325 462 -291 496
rect -325 394 -291 428
rect -325 326 -291 360
rect -325 258 -291 292
rect -325 190 -291 224
rect -325 122 -291 156
rect -325 54 -291 88
rect -325 -14 -291 20
rect -325 -82 -291 -48
rect -325 -150 -291 -116
rect -325 -218 -291 -184
rect -325 -286 -291 -252
rect -325 -354 -291 -320
rect -325 -422 -291 -388
rect -325 -490 -291 -456
rect -325 -558 -291 -524
rect -325 -626 -291 -592
rect -325 -694 -291 -660
rect -325 -762 -291 -728
rect -17 666 17 700
rect -17 598 17 632
rect -17 530 17 564
rect -17 462 17 496
rect -17 394 17 428
rect -17 326 17 360
rect -17 258 17 292
rect -17 190 17 224
rect -17 122 17 156
rect -17 54 17 88
rect -17 -14 17 20
rect -17 -82 17 -48
rect -17 -150 17 -116
rect -17 -218 17 -184
rect -17 -286 17 -252
rect -17 -354 17 -320
rect -17 -422 17 -388
rect -17 -490 17 -456
rect -17 -558 17 -524
rect -17 -626 17 -592
rect -17 -694 17 -660
rect -17 -762 17 -728
rect 291 666 325 700
rect 291 598 325 632
rect 291 530 325 564
rect 291 462 325 496
rect 291 394 325 428
rect 291 326 325 360
rect 291 258 325 292
rect 291 190 325 224
rect 291 122 325 156
rect 291 54 325 88
rect 291 -14 325 20
rect 291 -82 325 -48
rect 291 -150 325 -116
rect 291 -218 325 -184
rect 291 -286 325 -252
rect 291 -354 325 -320
rect 291 -422 325 -388
rect 291 -490 325 -456
rect 291 -558 325 -524
rect 291 -626 325 -592
rect 291 -694 325 -660
rect 291 -762 325 -728
rect 599 666 633 700
rect 599 598 633 632
rect 599 530 633 564
rect 599 462 633 496
rect 599 394 633 428
rect 599 326 633 360
rect 599 258 633 292
rect 599 190 633 224
rect 599 122 633 156
rect 599 54 633 88
rect 599 -14 633 20
rect 599 -82 633 -48
rect 599 -150 633 -116
rect 599 -218 633 -184
rect 599 -286 633 -252
rect 599 -354 633 -320
rect 599 -422 633 -388
rect 599 -490 633 -456
rect 599 -558 633 -524
rect 599 -626 633 -592
rect 599 -694 633 -660
rect 599 -762 633 -728
rect 907 666 941 700
rect 907 598 941 632
rect 907 530 941 564
rect 907 462 941 496
rect 907 394 941 428
rect 907 326 941 360
rect 907 258 941 292
rect 907 190 941 224
rect 907 122 941 156
rect 907 54 941 88
rect 907 -14 941 20
rect 907 -82 941 -48
rect 907 -150 941 -116
rect 907 -218 941 -184
rect 907 -286 941 -252
rect 907 -354 941 -320
rect 907 -422 941 -388
rect 907 -490 941 -456
rect 907 -558 941 -524
rect 907 -626 941 -592
rect 907 -694 941 -660
rect 907 -762 941 -728
rect 1215 666 1249 700
rect 1215 598 1249 632
rect 1215 530 1249 564
rect 1215 462 1249 496
rect 1215 394 1249 428
rect 1215 326 1249 360
rect 1215 258 1249 292
rect 1215 190 1249 224
rect 1215 122 1249 156
rect 1215 54 1249 88
rect 1215 -14 1249 20
rect 1215 -82 1249 -48
rect 1215 -150 1249 -116
rect 1215 -218 1249 -184
rect 1215 -286 1249 -252
rect 1215 -354 1249 -320
rect 1215 -422 1249 -388
rect 1215 -490 1249 -456
rect 1215 -558 1249 -524
rect 1215 -626 1249 -592
rect 1215 -694 1249 -660
rect 1215 -762 1249 -728
rect 1523 666 1557 700
rect 1523 598 1557 632
rect 1523 530 1557 564
rect 1523 462 1557 496
rect 1523 394 1557 428
rect 1523 326 1557 360
rect 1523 258 1557 292
rect 1523 190 1557 224
rect 1523 122 1557 156
rect 1523 54 1557 88
rect 1523 -14 1557 20
rect 1523 -82 1557 -48
rect 1523 -150 1557 -116
rect 1523 -218 1557 -184
rect 1523 -286 1557 -252
rect 1523 -354 1557 -320
rect 1523 -422 1557 -388
rect 1523 -490 1557 -456
rect 1523 -558 1557 -524
rect 1523 -626 1557 -592
rect 1523 -694 1557 -660
rect 1523 -762 1557 -728
rect 1831 666 1865 700
rect 1831 598 1865 632
rect 1831 530 1865 564
rect 1831 462 1865 496
rect 1831 394 1865 428
rect 1831 326 1865 360
rect 1831 258 1865 292
rect 1831 190 1865 224
rect 1831 122 1865 156
rect 1831 54 1865 88
rect 1831 -14 1865 20
rect 1831 -82 1865 -48
rect 1831 -150 1865 -116
rect 1831 -218 1865 -184
rect 1831 -286 1865 -252
rect 1831 -354 1865 -320
rect 1831 -422 1865 -388
rect 1831 -490 1865 -456
rect 1831 -558 1865 -524
rect 1831 -626 1865 -592
rect 1831 -694 1865 -660
rect 1831 -762 1865 -728
rect 2139 666 2173 700
rect 2139 598 2173 632
rect 2139 530 2173 564
rect 2139 462 2173 496
rect 2139 394 2173 428
rect 2139 326 2173 360
rect 2139 258 2173 292
rect 2139 190 2173 224
rect 2139 122 2173 156
rect 2139 54 2173 88
rect 2139 -14 2173 20
rect 2139 -82 2173 -48
rect 2139 -150 2173 -116
rect 2139 -218 2173 -184
rect 2139 -286 2173 -252
rect 2139 -354 2173 -320
rect 2139 -422 2173 -388
rect 2139 -490 2173 -456
rect 2139 -558 2173 -524
rect 2139 -626 2173 -592
rect 2139 -694 2173 -660
rect 2139 -762 2173 -728
rect 2447 666 2481 700
rect 2447 598 2481 632
rect 2447 530 2481 564
rect 2447 462 2481 496
rect 2447 394 2481 428
rect 2447 326 2481 360
rect 2447 258 2481 292
rect 2447 190 2481 224
rect 2447 122 2481 156
rect 2447 54 2481 88
rect 2447 -14 2481 20
rect 2447 -82 2481 -48
rect 2447 -150 2481 -116
rect 2447 -218 2481 -184
rect 2447 -286 2481 -252
rect 2447 -354 2481 -320
rect 2447 -422 2481 -388
rect 2447 -490 2481 -456
rect 2447 -558 2481 -524
rect 2447 -626 2481 -592
rect 2447 -694 2481 -660
rect 2447 -762 2481 -728
rect 2755 666 2789 700
rect 2755 598 2789 632
rect 2755 530 2789 564
rect 2755 462 2789 496
rect 2755 394 2789 428
rect 2755 326 2789 360
rect 2755 258 2789 292
rect 2755 190 2789 224
rect 2755 122 2789 156
rect 2755 54 2789 88
rect 2755 -14 2789 20
rect 2755 -82 2789 -48
rect 2755 -150 2789 -116
rect 2755 -218 2789 -184
rect 2755 -286 2789 -252
rect 2755 -354 2789 -320
rect 2755 -422 2789 -388
rect 2755 -490 2789 -456
rect 2755 -558 2789 -524
rect 2755 -626 2789 -592
rect 2755 -694 2789 -660
rect 2755 -762 2789 -728
<< poly >>
rect -2743 791 -2493 807
rect -2743 757 -2703 791
rect -2669 757 -2635 791
rect -2601 757 -2567 791
rect -2533 757 -2493 791
rect -2743 719 -2493 757
rect -2435 791 -2185 807
rect -2435 757 -2395 791
rect -2361 757 -2327 791
rect -2293 757 -2259 791
rect -2225 757 -2185 791
rect -2435 719 -2185 757
rect -2127 791 -1877 807
rect -2127 757 -2087 791
rect -2053 757 -2019 791
rect -1985 757 -1951 791
rect -1917 757 -1877 791
rect -2127 719 -1877 757
rect -1819 791 -1569 807
rect -1819 757 -1779 791
rect -1745 757 -1711 791
rect -1677 757 -1643 791
rect -1609 757 -1569 791
rect -1819 719 -1569 757
rect -1511 791 -1261 807
rect -1511 757 -1471 791
rect -1437 757 -1403 791
rect -1369 757 -1335 791
rect -1301 757 -1261 791
rect -1511 719 -1261 757
rect -1203 791 -953 807
rect -1203 757 -1163 791
rect -1129 757 -1095 791
rect -1061 757 -1027 791
rect -993 757 -953 791
rect -1203 719 -953 757
rect -895 791 -645 807
rect -895 757 -855 791
rect -821 757 -787 791
rect -753 757 -719 791
rect -685 757 -645 791
rect -895 719 -645 757
rect -587 791 -337 807
rect -587 757 -547 791
rect -513 757 -479 791
rect -445 757 -411 791
rect -377 757 -337 791
rect -587 719 -337 757
rect -279 791 -29 807
rect -279 757 -239 791
rect -205 757 -171 791
rect -137 757 -103 791
rect -69 757 -29 791
rect -279 719 -29 757
rect 29 791 279 807
rect 29 757 69 791
rect 103 757 137 791
rect 171 757 205 791
rect 239 757 279 791
rect 29 719 279 757
rect 337 791 587 807
rect 337 757 377 791
rect 411 757 445 791
rect 479 757 513 791
rect 547 757 587 791
rect 337 719 587 757
rect 645 791 895 807
rect 645 757 685 791
rect 719 757 753 791
rect 787 757 821 791
rect 855 757 895 791
rect 645 719 895 757
rect 953 791 1203 807
rect 953 757 993 791
rect 1027 757 1061 791
rect 1095 757 1129 791
rect 1163 757 1203 791
rect 953 719 1203 757
rect 1261 791 1511 807
rect 1261 757 1301 791
rect 1335 757 1369 791
rect 1403 757 1437 791
rect 1471 757 1511 791
rect 1261 719 1511 757
rect 1569 791 1819 807
rect 1569 757 1609 791
rect 1643 757 1677 791
rect 1711 757 1745 791
rect 1779 757 1819 791
rect 1569 719 1819 757
rect 1877 791 2127 807
rect 1877 757 1917 791
rect 1951 757 1985 791
rect 2019 757 2053 791
rect 2087 757 2127 791
rect 1877 719 2127 757
rect 2185 791 2435 807
rect 2185 757 2225 791
rect 2259 757 2293 791
rect 2327 757 2361 791
rect 2395 757 2435 791
rect 2185 719 2435 757
rect 2493 791 2743 807
rect 2493 757 2533 791
rect 2567 757 2601 791
rect 2635 757 2669 791
rect 2703 757 2743 791
rect 2493 719 2743 757
rect -2743 -807 -2493 -781
rect -2435 -807 -2185 -781
rect -2127 -807 -1877 -781
rect -1819 -807 -1569 -781
rect -1511 -807 -1261 -781
rect -1203 -807 -953 -781
rect -895 -807 -645 -781
rect -587 -807 -337 -781
rect -279 -807 -29 -781
rect 29 -807 279 -781
rect 337 -807 587 -781
rect 645 -807 895 -781
rect 953 -807 1203 -781
rect 1261 -807 1511 -781
rect 1569 -807 1819 -781
rect 1877 -807 2127 -781
rect 2185 -807 2435 -781
rect 2493 -807 2743 -781
<< polycont >>
rect -2703 757 -2669 791
rect -2635 757 -2601 791
rect -2567 757 -2533 791
rect -2395 757 -2361 791
rect -2327 757 -2293 791
rect -2259 757 -2225 791
rect -2087 757 -2053 791
rect -2019 757 -1985 791
rect -1951 757 -1917 791
rect -1779 757 -1745 791
rect -1711 757 -1677 791
rect -1643 757 -1609 791
rect -1471 757 -1437 791
rect -1403 757 -1369 791
rect -1335 757 -1301 791
rect -1163 757 -1129 791
rect -1095 757 -1061 791
rect -1027 757 -993 791
rect -855 757 -821 791
rect -787 757 -753 791
rect -719 757 -685 791
rect -547 757 -513 791
rect -479 757 -445 791
rect -411 757 -377 791
rect -239 757 -205 791
rect -171 757 -137 791
rect -103 757 -69 791
rect 69 757 103 791
rect 137 757 171 791
rect 205 757 239 791
rect 377 757 411 791
rect 445 757 479 791
rect 513 757 547 791
rect 685 757 719 791
rect 753 757 787 791
rect 821 757 855 791
rect 993 757 1027 791
rect 1061 757 1095 791
rect 1129 757 1163 791
rect 1301 757 1335 791
rect 1369 757 1403 791
rect 1437 757 1471 791
rect 1609 757 1643 791
rect 1677 757 1711 791
rect 1745 757 1779 791
rect 1917 757 1951 791
rect 1985 757 2019 791
rect 2053 757 2087 791
rect 2225 757 2259 791
rect 2293 757 2327 791
rect 2361 757 2395 791
rect 2533 757 2567 791
rect 2601 757 2635 791
rect 2669 757 2703 791
<< locali >>
rect -2743 757 -2707 791
rect -2669 757 -2635 791
rect -2601 757 -2567 791
rect -2529 757 -2493 791
rect -2435 757 -2399 791
rect -2361 757 -2327 791
rect -2293 757 -2259 791
rect -2221 757 -2185 791
rect -2127 757 -2091 791
rect -2053 757 -2019 791
rect -1985 757 -1951 791
rect -1913 757 -1877 791
rect -1819 757 -1783 791
rect -1745 757 -1711 791
rect -1677 757 -1643 791
rect -1605 757 -1569 791
rect -1511 757 -1475 791
rect -1437 757 -1403 791
rect -1369 757 -1335 791
rect -1297 757 -1261 791
rect -1203 757 -1167 791
rect -1129 757 -1095 791
rect -1061 757 -1027 791
rect -989 757 -953 791
rect -895 757 -859 791
rect -821 757 -787 791
rect -753 757 -719 791
rect -681 757 -645 791
rect -587 757 -551 791
rect -513 757 -479 791
rect -445 757 -411 791
rect -373 757 -337 791
rect -279 757 -243 791
rect -205 757 -171 791
rect -137 757 -103 791
rect -65 757 -29 791
rect 29 757 65 791
rect 103 757 137 791
rect 171 757 205 791
rect 243 757 279 791
rect 337 757 373 791
rect 411 757 445 791
rect 479 757 513 791
rect 551 757 587 791
rect 645 757 681 791
rect 719 757 753 791
rect 787 757 821 791
rect 859 757 895 791
rect 953 757 989 791
rect 1027 757 1061 791
rect 1095 757 1129 791
rect 1167 757 1203 791
rect 1261 757 1297 791
rect 1335 757 1369 791
rect 1403 757 1437 791
rect 1475 757 1511 791
rect 1569 757 1605 791
rect 1643 757 1677 791
rect 1711 757 1745 791
rect 1783 757 1819 791
rect 1877 757 1913 791
rect 1951 757 1985 791
rect 2019 757 2053 791
rect 2091 757 2127 791
rect 2185 757 2221 791
rect 2259 757 2293 791
rect 2327 757 2361 791
rect 2399 757 2435 791
rect 2493 757 2529 791
rect 2567 757 2601 791
rect 2635 757 2669 791
rect 2707 757 2743 791
rect -2789 706 -2755 723
rect -2789 634 -2755 666
rect -2789 564 -2755 598
rect -2789 496 -2755 528
rect -2789 428 -2755 456
rect -2789 360 -2755 384
rect -2789 292 -2755 312
rect -2789 224 -2755 240
rect -2789 156 -2755 168
rect -2789 88 -2755 96
rect -2789 20 -2755 24
rect -2789 -86 -2755 -82
rect -2789 -158 -2755 -150
rect -2789 -230 -2755 -218
rect -2789 -302 -2755 -286
rect -2789 -374 -2755 -354
rect -2789 -446 -2755 -422
rect -2789 -518 -2755 -490
rect -2789 -590 -2755 -558
rect -2789 -660 -2755 -626
rect -2789 -728 -2755 -696
rect -2789 -785 -2755 -768
rect -2481 706 -2447 723
rect -2481 634 -2447 666
rect -2481 564 -2447 598
rect -2481 496 -2447 528
rect -2481 428 -2447 456
rect -2481 360 -2447 384
rect -2481 292 -2447 312
rect -2481 224 -2447 240
rect -2481 156 -2447 168
rect -2481 88 -2447 96
rect -2481 20 -2447 24
rect -2481 -86 -2447 -82
rect -2481 -158 -2447 -150
rect -2481 -230 -2447 -218
rect -2481 -302 -2447 -286
rect -2481 -374 -2447 -354
rect -2481 -446 -2447 -422
rect -2481 -518 -2447 -490
rect -2481 -590 -2447 -558
rect -2481 -660 -2447 -626
rect -2481 -728 -2447 -696
rect -2481 -785 -2447 -768
rect -2173 706 -2139 723
rect -2173 634 -2139 666
rect -2173 564 -2139 598
rect -2173 496 -2139 528
rect -2173 428 -2139 456
rect -2173 360 -2139 384
rect -2173 292 -2139 312
rect -2173 224 -2139 240
rect -2173 156 -2139 168
rect -2173 88 -2139 96
rect -2173 20 -2139 24
rect -2173 -86 -2139 -82
rect -2173 -158 -2139 -150
rect -2173 -230 -2139 -218
rect -2173 -302 -2139 -286
rect -2173 -374 -2139 -354
rect -2173 -446 -2139 -422
rect -2173 -518 -2139 -490
rect -2173 -590 -2139 -558
rect -2173 -660 -2139 -626
rect -2173 -728 -2139 -696
rect -2173 -785 -2139 -768
rect -1865 706 -1831 723
rect -1865 634 -1831 666
rect -1865 564 -1831 598
rect -1865 496 -1831 528
rect -1865 428 -1831 456
rect -1865 360 -1831 384
rect -1865 292 -1831 312
rect -1865 224 -1831 240
rect -1865 156 -1831 168
rect -1865 88 -1831 96
rect -1865 20 -1831 24
rect -1865 -86 -1831 -82
rect -1865 -158 -1831 -150
rect -1865 -230 -1831 -218
rect -1865 -302 -1831 -286
rect -1865 -374 -1831 -354
rect -1865 -446 -1831 -422
rect -1865 -518 -1831 -490
rect -1865 -590 -1831 -558
rect -1865 -660 -1831 -626
rect -1865 -728 -1831 -696
rect -1865 -785 -1831 -768
rect -1557 706 -1523 723
rect -1557 634 -1523 666
rect -1557 564 -1523 598
rect -1557 496 -1523 528
rect -1557 428 -1523 456
rect -1557 360 -1523 384
rect -1557 292 -1523 312
rect -1557 224 -1523 240
rect -1557 156 -1523 168
rect -1557 88 -1523 96
rect -1557 20 -1523 24
rect -1557 -86 -1523 -82
rect -1557 -158 -1523 -150
rect -1557 -230 -1523 -218
rect -1557 -302 -1523 -286
rect -1557 -374 -1523 -354
rect -1557 -446 -1523 -422
rect -1557 -518 -1523 -490
rect -1557 -590 -1523 -558
rect -1557 -660 -1523 -626
rect -1557 -728 -1523 -696
rect -1557 -785 -1523 -768
rect -1249 706 -1215 723
rect -1249 634 -1215 666
rect -1249 564 -1215 598
rect -1249 496 -1215 528
rect -1249 428 -1215 456
rect -1249 360 -1215 384
rect -1249 292 -1215 312
rect -1249 224 -1215 240
rect -1249 156 -1215 168
rect -1249 88 -1215 96
rect -1249 20 -1215 24
rect -1249 -86 -1215 -82
rect -1249 -158 -1215 -150
rect -1249 -230 -1215 -218
rect -1249 -302 -1215 -286
rect -1249 -374 -1215 -354
rect -1249 -446 -1215 -422
rect -1249 -518 -1215 -490
rect -1249 -590 -1215 -558
rect -1249 -660 -1215 -626
rect -1249 -728 -1215 -696
rect -1249 -785 -1215 -768
rect -941 706 -907 723
rect -941 634 -907 666
rect -941 564 -907 598
rect -941 496 -907 528
rect -941 428 -907 456
rect -941 360 -907 384
rect -941 292 -907 312
rect -941 224 -907 240
rect -941 156 -907 168
rect -941 88 -907 96
rect -941 20 -907 24
rect -941 -86 -907 -82
rect -941 -158 -907 -150
rect -941 -230 -907 -218
rect -941 -302 -907 -286
rect -941 -374 -907 -354
rect -941 -446 -907 -422
rect -941 -518 -907 -490
rect -941 -590 -907 -558
rect -941 -660 -907 -626
rect -941 -728 -907 -696
rect -941 -785 -907 -768
rect -633 706 -599 723
rect -633 634 -599 666
rect -633 564 -599 598
rect -633 496 -599 528
rect -633 428 -599 456
rect -633 360 -599 384
rect -633 292 -599 312
rect -633 224 -599 240
rect -633 156 -599 168
rect -633 88 -599 96
rect -633 20 -599 24
rect -633 -86 -599 -82
rect -633 -158 -599 -150
rect -633 -230 -599 -218
rect -633 -302 -599 -286
rect -633 -374 -599 -354
rect -633 -446 -599 -422
rect -633 -518 -599 -490
rect -633 -590 -599 -558
rect -633 -660 -599 -626
rect -633 -728 -599 -696
rect -633 -785 -599 -768
rect -325 706 -291 723
rect -325 634 -291 666
rect -325 564 -291 598
rect -325 496 -291 528
rect -325 428 -291 456
rect -325 360 -291 384
rect -325 292 -291 312
rect -325 224 -291 240
rect -325 156 -291 168
rect -325 88 -291 96
rect -325 20 -291 24
rect -325 -86 -291 -82
rect -325 -158 -291 -150
rect -325 -230 -291 -218
rect -325 -302 -291 -286
rect -325 -374 -291 -354
rect -325 -446 -291 -422
rect -325 -518 -291 -490
rect -325 -590 -291 -558
rect -325 -660 -291 -626
rect -325 -728 -291 -696
rect -325 -785 -291 -768
rect -17 706 17 723
rect -17 634 17 666
rect -17 564 17 598
rect -17 496 17 528
rect -17 428 17 456
rect -17 360 17 384
rect -17 292 17 312
rect -17 224 17 240
rect -17 156 17 168
rect -17 88 17 96
rect -17 20 17 24
rect -17 -86 17 -82
rect -17 -158 17 -150
rect -17 -230 17 -218
rect -17 -302 17 -286
rect -17 -374 17 -354
rect -17 -446 17 -422
rect -17 -518 17 -490
rect -17 -590 17 -558
rect -17 -660 17 -626
rect -17 -728 17 -696
rect -17 -785 17 -768
rect 291 706 325 723
rect 291 634 325 666
rect 291 564 325 598
rect 291 496 325 528
rect 291 428 325 456
rect 291 360 325 384
rect 291 292 325 312
rect 291 224 325 240
rect 291 156 325 168
rect 291 88 325 96
rect 291 20 325 24
rect 291 -86 325 -82
rect 291 -158 325 -150
rect 291 -230 325 -218
rect 291 -302 325 -286
rect 291 -374 325 -354
rect 291 -446 325 -422
rect 291 -518 325 -490
rect 291 -590 325 -558
rect 291 -660 325 -626
rect 291 -728 325 -696
rect 291 -785 325 -768
rect 599 706 633 723
rect 599 634 633 666
rect 599 564 633 598
rect 599 496 633 528
rect 599 428 633 456
rect 599 360 633 384
rect 599 292 633 312
rect 599 224 633 240
rect 599 156 633 168
rect 599 88 633 96
rect 599 20 633 24
rect 599 -86 633 -82
rect 599 -158 633 -150
rect 599 -230 633 -218
rect 599 -302 633 -286
rect 599 -374 633 -354
rect 599 -446 633 -422
rect 599 -518 633 -490
rect 599 -590 633 -558
rect 599 -660 633 -626
rect 599 -728 633 -696
rect 599 -785 633 -768
rect 907 706 941 723
rect 907 634 941 666
rect 907 564 941 598
rect 907 496 941 528
rect 907 428 941 456
rect 907 360 941 384
rect 907 292 941 312
rect 907 224 941 240
rect 907 156 941 168
rect 907 88 941 96
rect 907 20 941 24
rect 907 -86 941 -82
rect 907 -158 941 -150
rect 907 -230 941 -218
rect 907 -302 941 -286
rect 907 -374 941 -354
rect 907 -446 941 -422
rect 907 -518 941 -490
rect 907 -590 941 -558
rect 907 -660 941 -626
rect 907 -728 941 -696
rect 907 -785 941 -768
rect 1215 706 1249 723
rect 1215 634 1249 666
rect 1215 564 1249 598
rect 1215 496 1249 528
rect 1215 428 1249 456
rect 1215 360 1249 384
rect 1215 292 1249 312
rect 1215 224 1249 240
rect 1215 156 1249 168
rect 1215 88 1249 96
rect 1215 20 1249 24
rect 1215 -86 1249 -82
rect 1215 -158 1249 -150
rect 1215 -230 1249 -218
rect 1215 -302 1249 -286
rect 1215 -374 1249 -354
rect 1215 -446 1249 -422
rect 1215 -518 1249 -490
rect 1215 -590 1249 -558
rect 1215 -660 1249 -626
rect 1215 -728 1249 -696
rect 1215 -785 1249 -768
rect 1523 706 1557 723
rect 1523 634 1557 666
rect 1523 564 1557 598
rect 1523 496 1557 528
rect 1523 428 1557 456
rect 1523 360 1557 384
rect 1523 292 1557 312
rect 1523 224 1557 240
rect 1523 156 1557 168
rect 1523 88 1557 96
rect 1523 20 1557 24
rect 1523 -86 1557 -82
rect 1523 -158 1557 -150
rect 1523 -230 1557 -218
rect 1523 -302 1557 -286
rect 1523 -374 1557 -354
rect 1523 -446 1557 -422
rect 1523 -518 1557 -490
rect 1523 -590 1557 -558
rect 1523 -660 1557 -626
rect 1523 -728 1557 -696
rect 1523 -785 1557 -768
rect 1831 706 1865 723
rect 1831 634 1865 666
rect 1831 564 1865 598
rect 1831 496 1865 528
rect 1831 428 1865 456
rect 1831 360 1865 384
rect 1831 292 1865 312
rect 1831 224 1865 240
rect 1831 156 1865 168
rect 1831 88 1865 96
rect 1831 20 1865 24
rect 1831 -86 1865 -82
rect 1831 -158 1865 -150
rect 1831 -230 1865 -218
rect 1831 -302 1865 -286
rect 1831 -374 1865 -354
rect 1831 -446 1865 -422
rect 1831 -518 1865 -490
rect 1831 -590 1865 -558
rect 1831 -660 1865 -626
rect 1831 -728 1865 -696
rect 1831 -785 1865 -768
rect 2139 706 2173 723
rect 2139 634 2173 666
rect 2139 564 2173 598
rect 2139 496 2173 528
rect 2139 428 2173 456
rect 2139 360 2173 384
rect 2139 292 2173 312
rect 2139 224 2173 240
rect 2139 156 2173 168
rect 2139 88 2173 96
rect 2139 20 2173 24
rect 2139 -86 2173 -82
rect 2139 -158 2173 -150
rect 2139 -230 2173 -218
rect 2139 -302 2173 -286
rect 2139 -374 2173 -354
rect 2139 -446 2173 -422
rect 2139 -518 2173 -490
rect 2139 -590 2173 -558
rect 2139 -660 2173 -626
rect 2139 -728 2173 -696
rect 2139 -785 2173 -768
rect 2447 706 2481 723
rect 2447 634 2481 666
rect 2447 564 2481 598
rect 2447 496 2481 528
rect 2447 428 2481 456
rect 2447 360 2481 384
rect 2447 292 2481 312
rect 2447 224 2481 240
rect 2447 156 2481 168
rect 2447 88 2481 96
rect 2447 20 2481 24
rect 2447 -86 2481 -82
rect 2447 -158 2481 -150
rect 2447 -230 2481 -218
rect 2447 -302 2481 -286
rect 2447 -374 2481 -354
rect 2447 -446 2481 -422
rect 2447 -518 2481 -490
rect 2447 -590 2481 -558
rect 2447 -660 2481 -626
rect 2447 -728 2481 -696
rect 2447 -785 2481 -768
rect 2755 706 2789 723
rect 2755 634 2789 666
rect 2755 564 2789 598
rect 2755 496 2789 528
rect 2755 428 2789 456
rect 2755 360 2789 384
rect 2755 292 2789 312
rect 2755 224 2789 240
rect 2755 156 2789 168
rect 2755 88 2789 96
rect 2755 20 2789 24
rect 2755 -86 2789 -82
rect 2755 -158 2789 -150
rect 2755 -230 2789 -218
rect 2755 -302 2789 -286
rect 2755 -374 2789 -354
rect 2755 -446 2789 -422
rect 2755 -518 2789 -490
rect 2755 -590 2789 -558
rect 2755 -660 2789 -626
rect 2755 -728 2789 -696
rect 2755 -785 2789 -768
<< viali >>
rect -2707 757 -2703 791
rect -2703 757 -2673 791
rect -2635 757 -2601 791
rect -2563 757 -2533 791
rect -2533 757 -2529 791
rect -2399 757 -2395 791
rect -2395 757 -2365 791
rect -2327 757 -2293 791
rect -2255 757 -2225 791
rect -2225 757 -2221 791
rect -2091 757 -2087 791
rect -2087 757 -2057 791
rect -2019 757 -1985 791
rect -1947 757 -1917 791
rect -1917 757 -1913 791
rect -1783 757 -1779 791
rect -1779 757 -1749 791
rect -1711 757 -1677 791
rect -1639 757 -1609 791
rect -1609 757 -1605 791
rect -1475 757 -1471 791
rect -1471 757 -1441 791
rect -1403 757 -1369 791
rect -1331 757 -1301 791
rect -1301 757 -1297 791
rect -1167 757 -1163 791
rect -1163 757 -1133 791
rect -1095 757 -1061 791
rect -1023 757 -993 791
rect -993 757 -989 791
rect -859 757 -855 791
rect -855 757 -825 791
rect -787 757 -753 791
rect -715 757 -685 791
rect -685 757 -681 791
rect -551 757 -547 791
rect -547 757 -517 791
rect -479 757 -445 791
rect -407 757 -377 791
rect -377 757 -373 791
rect -243 757 -239 791
rect -239 757 -209 791
rect -171 757 -137 791
rect -99 757 -69 791
rect -69 757 -65 791
rect 65 757 69 791
rect 69 757 99 791
rect 137 757 171 791
rect 209 757 239 791
rect 239 757 243 791
rect 373 757 377 791
rect 377 757 407 791
rect 445 757 479 791
rect 517 757 547 791
rect 547 757 551 791
rect 681 757 685 791
rect 685 757 715 791
rect 753 757 787 791
rect 825 757 855 791
rect 855 757 859 791
rect 989 757 993 791
rect 993 757 1023 791
rect 1061 757 1095 791
rect 1133 757 1163 791
rect 1163 757 1167 791
rect 1297 757 1301 791
rect 1301 757 1331 791
rect 1369 757 1403 791
rect 1441 757 1471 791
rect 1471 757 1475 791
rect 1605 757 1609 791
rect 1609 757 1639 791
rect 1677 757 1711 791
rect 1749 757 1779 791
rect 1779 757 1783 791
rect 1913 757 1917 791
rect 1917 757 1947 791
rect 1985 757 2019 791
rect 2057 757 2087 791
rect 2087 757 2091 791
rect 2221 757 2225 791
rect 2225 757 2255 791
rect 2293 757 2327 791
rect 2365 757 2395 791
rect 2395 757 2399 791
rect 2529 757 2533 791
rect 2533 757 2563 791
rect 2601 757 2635 791
rect 2673 757 2703 791
rect 2703 757 2707 791
rect -2789 700 -2755 706
rect -2789 672 -2755 700
rect -2789 632 -2755 634
rect -2789 600 -2755 632
rect -2789 530 -2755 562
rect -2789 528 -2755 530
rect -2789 462 -2755 490
rect -2789 456 -2755 462
rect -2789 394 -2755 418
rect -2789 384 -2755 394
rect -2789 326 -2755 346
rect -2789 312 -2755 326
rect -2789 258 -2755 274
rect -2789 240 -2755 258
rect -2789 190 -2755 202
rect -2789 168 -2755 190
rect -2789 122 -2755 130
rect -2789 96 -2755 122
rect -2789 54 -2755 58
rect -2789 24 -2755 54
rect -2789 -48 -2755 -14
rect -2789 -116 -2755 -86
rect -2789 -120 -2755 -116
rect -2789 -184 -2755 -158
rect -2789 -192 -2755 -184
rect -2789 -252 -2755 -230
rect -2789 -264 -2755 -252
rect -2789 -320 -2755 -302
rect -2789 -336 -2755 -320
rect -2789 -388 -2755 -374
rect -2789 -408 -2755 -388
rect -2789 -456 -2755 -446
rect -2789 -480 -2755 -456
rect -2789 -524 -2755 -518
rect -2789 -552 -2755 -524
rect -2789 -592 -2755 -590
rect -2789 -624 -2755 -592
rect -2789 -694 -2755 -662
rect -2789 -696 -2755 -694
rect -2789 -762 -2755 -734
rect -2789 -768 -2755 -762
rect -2481 700 -2447 706
rect -2481 672 -2447 700
rect -2481 632 -2447 634
rect -2481 600 -2447 632
rect -2481 530 -2447 562
rect -2481 528 -2447 530
rect -2481 462 -2447 490
rect -2481 456 -2447 462
rect -2481 394 -2447 418
rect -2481 384 -2447 394
rect -2481 326 -2447 346
rect -2481 312 -2447 326
rect -2481 258 -2447 274
rect -2481 240 -2447 258
rect -2481 190 -2447 202
rect -2481 168 -2447 190
rect -2481 122 -2447 130
rect -2481 96 -2447 122
rect -2481 54 -2447 58
rect -2481 24 -2447 54
rect -2481 -48 -2447 -14
rect -2481 -116 -2447 -86
rect -2481 -120 -2447 -116
rect -2481 -184 -2447 -158
rect -2481 -192 -2447 -184
rect -2481 -252 -2447 -230
rect -2481 -264 -2447 -252
rect -2481 -320 -2447 -302
rect -2481 -336 -2447 -320
rect -2481 -388 -2447 -374
rect -2481 -408 -2447 -388
rect -2481 -456 -2447 -446
rect -2481 -480 -2447 -456
rect -2481 -524 -2447 -518
rect -2481 -552 -2447 -524
rect -2481 -592 -2447 -590
rect -2481 -624 -2447 -592
rect -2481 -694 -2447 -662
rect -2481 -696 -2447 -694
rect -2481 -762 -2447 -734
rect -2481 -768 -2447 -762
rect -2173 700 -2139 706
rect -2173 672 -2139 700
rect -2173 632 -2139 634
rect -2173 600 -2139 632
rect -2173 530 -2139 562
rect -2173 528 -2139 530
rect -2173 462 -2139 490
rect -2173 456 -2139 462
rect -2173 394 -2139 418
rect -2173 384 -2139 394
rect -2173 326 -2139 346
rect -2173 312 -2139 326
rect -2173 258 -2139 274
rect -2173 240 -2139 258
rect -2173 190 -2139 202
rect -2173 168 -2139 190
rect -2173 122 -2139 130
rect -2173 96 -2139 122
rect -2173 54 -2139 58
rect -2173 24 -2139 54
rect -2173 -48 -2139 -14
rect -2173 -116 -2139 -86
rect -2173 -120 -2139 -116
rect -2173 -184 -2139 -158
rect -2173 -192 -2139 -184
rect -2173 -252 -2139 -230
rect -2173 -264 -2139 -252
rect -2173 -320 -2139 -302
rect -2173 -336 -2139 -320
rect -2173 -388 -2139 -374
rect -2173 -408 -2139 -388
rect -2173 -456 -2139 -446
rect -2173 -480 -2139 -456
rect -2173 -524 -2139 -518
rect -2173 -552 -2139 -524
rect -2173 -592 -2139 -590
rect -2173 -624 -2139 -592
rect -2173 -694 -2139 -662
rect -2173 -696 -2139 -694
rect -2173 -762 -2139 -734
rect -2173 -768 -2139 -762
rect -1865 700 -1831 706
rect -1865 672 -1831 700
rect -1865 632 -1831 634
rect -1865 600 -1831 632
rect -1865 530 -1831 562
rect -1865 528 -1831 530
rect -1865 462 -1831 490
rect -1865 456 -1831 462
rect -1865 394 -1831 418
rect -1865 384 -1831 394
rect -1865 326 -1831 346
rect -1865 312 -1831 326
rect -1865 258 -1831 274
rect -1865 240 -1831 258
rect -1865 190 -1831 202
rect -1865 168 -1831 190
rect -1865 122 -1831 130
rect -1865 96 -1831 122
rect -1865 54 -1831 58
rect -1865 24 -1831 54
rect -1865 -48 -1831 -14
rect -1865 -116 -1831 -86
rect -1865 -120 -1831 -116
rect -1865 -184 -1831 -158
rect -1865 -192 -1831 -184
rect -1865 -252 -1831 -230
rect -1865 -264 -1831 -252
rect -1865 -320 -1831 -302
rect -1865 -336 -1831 -320
rect -1865 -388 -1831 -374
rect -1865 -408 -1831 -388
rect -1865 -456 -1831 -446
rect -1865 -480 -1831 -456
rect -1865 -524 -1831 -518
rect -1865 -552 -1831 -524
rect -1865 -592 -1831 -590
rect -1865 -624 -1831 -592
rect -1865 -694 -1831 -662
rect -1865 -696 -1831 -694
rect -1865 -762 -1831 -734
rect -1865 -768 -1831 -762
rect -1557 700 -1523 706
rect -1557 672 -1523 700
rect -1557 632 -1523 634
rect -1557 600 -1523 632
rect -1557 530 -1523 562
rect -1557 528 -1523 530
rect -1557 462 -1523 490
rect -1557 456 -1523 462
rect -1557 394 -1523 418
rect -1557 384 -1523 394
rect -1557 326 -1523 346
rect -1557 312 -1523 326
rect -1557 258 -1523 274
rect -1557 240 -1523 258
rect -1557 190 -1523 202
rect -1557 168 -1523 190
rect -1557 122 -1523 130
rect -1557 96 -1523 122
rect -1557 54 -1523 58
rect -1557 24 -1523 54
rect -1557 -48 -1523 -14
rect -1557 -116 -1523 -86
rect -1557 -120 -1523 -116
rect -1557 -184 -1523 -158
rect -1557 -192 -1523 -184
rect -1557 -252 -1523 -230
rect -1557 -264 -1523 -252
rect -1557 -320 -1523 -302
rect -1557 -336 -1523 -320
rect -1557 -388 -1523 -374
rect -1557 -408 -1523 -388
rect -1557 -456 -1523 -446
rect -1557 -480 -1523 -456
rect -1557 -524 -1523 -518
rect -1557 -552 -1523 -524
rect -1557 -592 -1523 -590
rect -1557 -624 -1523 -592
rect -1557 -694 -1523 -662
rect -1557 -696 -1523 -694
rect -1557 -762 -1523 -734
rect -1557 -768 -1523 -762
rect -1249 700 -1215 706
rect -1249 672 -1215 700
rect -1249 632 -1215 634
rect -1249 600 -1215 632
rect -1249 530 -1215 562
rect -1249 528 -1215 530
rect -1249 462 -1215 490
rect -1249 456 -1215 462
rect -1249 394 -1215 418
rect -1249 384 -1215 394
rect -1249 326 -1215 346
rect -1249 312 -1215 326
rect -1249 258 -1215 274
rect -1249 240 -1215 258
rect -1249 190 -1215 202
rect -1249 168 -1215 190
rect -1249 122 -1215 130
rect -1249 96 -1215 122
rect -1249 54 -1215 58
rect -1249 24 -1215 54
rect -1249 -48 -1215 -14
rect -1249 -116 -1215 -86
rect -1249 -120 -1215 -116
rect -1249 -184 -1215 -158
rect -1249 -192 -1215 -184
rect -1249 -252 -1215 -230
rect -1249 -264 -1215 -252
rect -1249 -320 -1215 -302
rect -1249 -336 -1215 -320
rect -1249 -388 -1215 -374
rect -1249 -408 -1215 -388
rect -1249 -456 -1215 -446
rect -1249 -480 -1215 -456
rect -1249 -524 -1215 -518
rect -1249 -552 -1215 -524
rect -1249 -592 -1215 -590
rect -1249 -624 -1215 -592
rect -1249 -694 -1215 -662
rect -1249 -696 -1215 -694
rect -1249 -762 -1215 -734
rect -1249 -768 -1215 -762
rect -941 700 -907 706
rect -941 672 -907 700
rect -941 632 -907 634
rect -941 600 -907 632
rect -941 530 -907 562
rect -941 528 -907 530
rect -941 462 -907 490
rect -941 456 -907 462
rect -941 394 -907 418
rect -941 384 -907 394
rect -941 326 -907 346
rect -941 312 -907 326
rect -941 258 -907 274
rect -941 240 -907 258
rect -941 190 -907 202
rect -941 168 -907 190
rect -941 122 -907 130
rect -941 96 -907 122
rect -941 54 -907 58
rect -941 24 -907 54
rect -941 -48 -907 -14
rect -941 -116 -907 -86
rect -941 -120 -907 -116
rect -941 -184 -907 -158
rect -941 -192 -907 -184
rect -941 -252 -907 -230
rect -941 -264 -907 -252
rect -941 -320 -907 -302
rect -941 -336 -907 -320
rect -941 -388 -907 -374
rect -941 -408 -907 -388
rect -941 -456 -907 -446
rect -941 -480 -907 -456
rect -941 -524 -907 -518
rect -941 -552 -907 -524
rect -941 -592 -907 -590
rect -941 -624 -907 -592
rect -941 -694 -907 -662
rect -941 -696 -907 -694
rect -941 -762 -907 -734
rect -941 -768 -907 -762
rect -633 700 -599 706
rect -633 672 -599 700
rect -633 632 -599 634
rect -633 600 -599 632
rect -633 530 -599 562
rect -633 528 -599 530
rect -633 462 -599 490
rect -633 456 -599 462
rect -633 394 -599 418
rect -633 384 -599 394
rect -633 326 -599 346
rect -633 312 -599 326
rect -633 258 -599 274
rect -633 240 -599 258
rect -633 190 -599 202
rect -633 168 -599 190
rect -633 122 -599 130
rect -633 96 -599 122
rect -633 54 -599 58
rect -633 24 -599 54
rect -633 -48 -599 -14
rect -633 -116 -599 -86
rect -633 -120 -599 -116
rect -633 -184 -599 -158
rect -633 -192 -599 -184
rect -633 -252 -599 -230
rect -633 -264 -599 -252
rect -633 -320 -599 -302
rect -633 -336 -599 -320
rect -633 -388 -599 -374
rect -633 -408 -599 -388
rect -633 -456 -599 -446
rect -633 -480 -599 -456
rect -633 -524 -599 -518
rect -633 -552 -599 -524
rect -633 -592 -599 -590
rect -633 -624 -599 -592
rect -633 -694 -599 -662
rect -633 -696 -599 -694
rect -633 -762 -599 -734
rect -633 -768 -599 -762
rect -325 700 -291 706
rect -325 672 -291 700
rect -325 632 -291 634
rect -325 600 -291 632
rect -325 530 -291 562
rect -325 528 -291 530
rect -325 462 -291 490
rect -325 456 -291 462
rect -325 394 -291 418
rect -325 384 -291 394
rect -325 326 -291 346
rect -325 312 -291 326
rect -325 258 -291 274
rect -325 240 -291 258
rect -325 190 -291 202
rect -325 168 -291 190
rect -325 122 -291 130
rect -325 96 -291 122
rect -325 54 -291 58
rect -325 24 -291 54
rect -325 -48 -291 -14
rect -325 -116 -291 -86
rect -325 -120 -291 -116
rect -325 -184 -291 -158
rect -325 -192 -291 -184
rect -325 -252 -291 -230
rect -325 -264 -291 -252
rect -325 -320 -291 -302
rect -325 -336 -291 -320
rect -325 -388 -291 -374
rect -325 -408 -291 -388
rect -325 -456 -291 -446
rect -325 -480 -291 -456
rect -325 -524 -291 -518
rect -325 -552 -291 -524
rect -325 -592 -291 -590
rect -325 -624 -291 -592
rect -325 -694 -291 -662
rect -325 -696 -291 -694
rect -325 -762 -291 -734
rect -325 -768 -291 -762
rect -17 700 17 706
rect -17 672 17 700
rect -17 632 17 634
rect -17 600 17 632
rect -17 530 17 562
rect -17 528 17 530
rect -17 462 17 490
rect -17 456 17 462
rect -17 394 17 418
rect -17 384 17 394
rect -17 326 17 346
rect -17 312 17 326
rect -17 258 17 274
rect -17 240 17 258
rect -17 190 17 202
rect -17 168 17 190
rect -17 122 17 130
rect -17 96 17 122
rect -17 54 17 58
rect -17 24 17 54
rect -17 -48 17 -14
rect -17 -116 17 -86
rect -17 -120 17 -116
rect -17 -184 17 -158
rect -17 -192 17 -184
rect -17 -252 17 -230
rect -17 -264 17 -252
rect -17 -320 17 -302
rect -17 -336 17 -320
rect -17 -388 17 -374
rect -17 -408 17 -388
rect -17 -456 17 -446
rect -17 -480 17 -456
rect -17 -524 17 -518
rect -17 -552 17 -524
rect -17 -592 17 -590
rect -17 -624 17 -592
rect -17 -694 17 -662
rect -17 -696 17 -694
rect -17 -762 17 -734
rect -17 -768 17 -762
rect 291 700 325 706
rect 291 672 325 700
rect 291 632 325 634
rect 291 600 325 632
rect 291 530 325 562
rect 291 528 325 530
rect 291 462 325 490
rect 291 456 325 462
rect 291 394 325 418
rect 291 384 325 394
rect 291 326 325 346
rect 291 312 325 326
rect 291 258 325 274
rect 291 240 325 258
rect 291 190 325 202
rect 291 168 325 190
rect 291 122 325 130
rect 291 96 325 122
rect 291 54 325 58
rect 291 24 325 54
rect 291 -48 325 -14
rect 291 -116 325 -86
rect 291 -120 325 -116
rect 291 -184 325 -158
rect 291 -192 325 -184
rect 291 -252 325 -230
rect 291 -264 325 -252
rect 291 -320 325 -302
rect 291 -336 325 -320
rect 291 -388 325 -374
rect 291 -408 325 -388
rect 291 -456 325 -446
rect 291 -480 325 -456
rect 291 -524 325 -518
rect 291 -552 325 -524
rect 291 -592 325 -590
rect 291 -624 325 -592
rect 291 -694 325 -662
rect 291 -696 325 -694
rect 291 -762 325 -734
rect 291 -768 325 -762
rect 599 700 633 706
rect 599 672 633 700
rect 599 632 633 634
rect 599 600 633 632
rect 599 530 633 562
rect 599 528 633 530
rect 599 462 633 490
rect 599 456 633 462
rect 599 394 633 418
rect 599 384 633 394
rect 599 326 633 346
rect 599 312 633 326
rect 599 258 633 274
rect 599 240 633 258
rect 599 190 633 202
rect 599 168 633 190
rect 599 122 633 130
rect 599 96 633 122
rect 599 54 633 58
rect 599 24 633 54
rect 599 -48 633 -14
rect 599 -116 633 -86
rect 599 -120 633 -116
rect 599 -184 633 -158
rect 599 -192 633 -184
rect 599 -252 633 -230
rect 599 -264 633 -252
rect 599 -320 633 -302
rect 599 -336 633 -320
rect 599 -388 633 -374
rect 599 -408 633 -388
rect 599 -456 633 -446
rect 599 -480 633 -456
rect 599 -524 633 -518
rect 599 -552 633 -524
rect 599 -592 633 -590
rect 599 -624 633 -592
rect 599 -694 633 -662
rect 599 -696 633 -694
rect 599 -762 633 -734
rect 599 -768 633 -762
rect 907 700 941 706
rect 907 672 941 700
rect 907 632 941 634
rect 907 600 941 632
rect 907 530 941 562
rect 907 528 941 530
rect 907 462 941 490
rect 907 456 941 462
rect 907 394 941 418
rect 907 384 941 394
rect 907 326 941 346
rect 907 312 941 326
rect 907 258 941 274
rect 907 240 941 258
rect 907 190 941 202
rect 907 168 941 190
rect 907 122 941 130
rect 907 96 941 122
rect 907 54 941 58
rect 907 24 941 54
rect 907 -48 941 -14
rect 907 -116 941 -86
rect 907 -120 941 -116
rect 907 -184 941 -158
rect 907 -192 941 -184
rect 907 -252 941 -230
rect 907 -264 941 -252
rect 907 -320 941 -302
rect 907 -336 941 -320
rect 907 -388 941 -374
rect 907 -408 941 -388
rect 907 -456 941 -446
rect 907 -480 941 -456
rect 907 -524 941 -518
rect 907 -552 941 -524
rect 907 -592 941 -590
rect 907 -624 941 -592
rect 907 -694 941 -662
rect 907 -696 941 -694
rect 907 -762 941 -734
rect 907 -768 941 -762
rect 1215 700 1249 706
rect 1215 672 1249 700
rect 1215 632 1249 634
rect 1215 600 1249 632
rect 1215 530 1249 562
rect 1215 528 1249 530
rect 1215 462 1249 490
rect 1215 456 1249 462
rect 1215 394 1249 418
rect 1215 384 1249 394
rect 1215 326 1249 346
rect 1215 312 1249 326
rect 1215 258 1249 274
rect 1215 240 1249 258
rect 1215 190 1249 202
rect 1215 168 1249 190
rect 1215 122 1249 130
rect 1215 96 1249 122
rect 1215 54 1249 58
rect 1215 24 1249 54
rect 1215 -48 1249 -14
rect 1215 -116 1249 -86
rect 1215 -120 1249 -116
rect 1215 -184 1249 -158
rect 1215 -192 1249 -184
rect 1215 -252 1249 -230
rect 1215 -264 1249 -252
rect 1215 -320 1249 -302
rect 1215 -336 1249 -320
rect 1215 -388 1249 -374
rect 1215 -408 1249 -388
rect 1215 -456 1249 -446
rect 1215 -480 1249 -456
rect 1215 -524 1249 -518
rect 1215 -552 1249 -524
rect 1215 -592 1249 -590
rect 1215 -624 1249 -592
rect 1215 -694 1249 -662
rect 1215 -696 1249 -694
rect 1215 -762 1249 -734
rect 1215 -768 1249 -762
rect 1523 700 1557 706
rect 1523 672 1557 700
rect 1523 632 1557 634
rect 1523 600 1557 632
rect 1523 530 1557 562
rect 1523 528 1557 530
rect 1523 462 1557 490
rect 1523 456 1557 462
rect 1523 394 1557 418
rect 1523 384 1557 394
rect 1523 326 1557 346
rect 1523 312 1557 326
rect 1523 258 1557 274
rect 1523 240 1557 258
rect 1523 190 1557 202
rect 1523 168 1557 190
rect 1523 122 1557 130
rect 1523 96 1557 122
rect 1523 54 1557 58
rect 1523 24 1557 54
rect 1523 -48 1557 -14
rect 1523 -116 1557 -86
rect 1523 -120 1557 -116
rect 1523 -184 1557 -158
rect 1523 -192 1557 -184
rect 1523 -252 1557 -230
rect 1523 -264 1557 -252
rect 1523 -320 1557 -302
rect 1523 -336 1557 -320
rect 1523 -388 1557 -374
rect 1523 -408 1557 -388
rect 1523 -456 1557 -446
rect 1523 -480 1557 -456
rect 1523 -524 1557 -518
rect 1523 -552 1557 -524
rect 1523 -592 1557 -590
rect 1523 -624 1557 -592
rect 1523 -694 1557 -662
rect 1523 -696 1557 -694
rect 1523 -762 1557 -734
rect 1523 -768 1557 -762
rect 1831 700 1865 706
rect 1831 672 1865 700
rect 1831 632 1865 634
rect 1831 600 1865 632
rect 1831 530 1865 562
rect 1831 528 1865 530
rect 1831 462 1865 490
rect 1831 456 1865 462
rect 1831 394 1865 418
rect 1831 384 1865 394
rect 1831 326 1865 346
rect 1831 312 1865 326
rect 1831 258 1865 274
rect 1831 240 1865 258
rect 1831 190 1865 202
rect 1831 168 1865 190
rect 1831 122 1865 130
rect 1831 96 1865 122
rect 1831 54 1865 58
rect 1831 24 1865 54
rect 1831 -48 1865 -14
rect 1831 -116 1865 -86
rect 1831 -120 1865 -116
rect 1831 -184 1865 -158
rect 1831 -192 1865 -184
rect 1831 -252 1865 -230
rect 1831 -264 1865 -252
rect 1831 -320 1865 -302
rect 1831 -336 1865 -320
rect 1831 -388 1865 -374
rect 1831 -408 1865 -388
rect 1831 -456 1865 -446
rect 1831 -480 1865 -456
rect 1831 -524 1865 -518
rect 1831 -552 1865 -524
rect 1831 -592 1865 -590
rect 1831 -624 1865 -592
rect 1831 -694 1865 -662
rect 1831 -696 1865 -694
rect 1831 -762 1865 -734
rect 1831 -768 1865 -762
rect 2139 700 2173 706
rect 2139 672 2173 700
rect 2139 632 2173 634
rect 2139 600 2173 632
rect 2139 530 2173 562
rect 2139 528 2173 530
rect 2139 462 2173 490
rect 2139 456 2173 462
rect 2139 394 2173 418
rect 2139 384 2173 394
rect 2139 326 2173 346
rect 2139 312 2173 326
rect 2139 258 2173 274
rect 2139 240 2173 258
rect 2139 190 2173 202
rect 2139 168 2173 190
rect 2139 122 2173 130
rect 2139 96 2173 122
rect 2139 54 2173 58
rect 2139 24 2173 54
rect 2139 -48 2173 -14
rect 2139 -116 2173 -86
rect 2139 -120 2173 -116
rect 2139 -184 2173 -158
rect 2139 -192 2173 -184
rect 2139 -252 2173 -230
rect 2139 -264 2173 -252
rect 2139 -320 2173 -302
rect 2139 -336 2173 -320
rect 2139 -388 2173 -374
rect 2139 -408 2173 -388
rect 2139 -456 2173 -446
rect 2139 -480 2173 -456
rect 2139 -524 2173 -518
rect 2139 -552 2173 -524
rect 2139 -592 2173 -590
rect 2139 -624 2173 -592
rect 2139 -694 2173 -662
rect 2139 -696 2173 -694
rect 2139 -762 2173 -734
rect 2139 -768 2173 -762
rect 2447 700 2481 706
rect 2447 672 2481 700
rect 2447 632 2481 634
rect 2447 600 2481 632
rect 2447 530 2481 562
rect 2447 528 2481 530
rect 2447 462 2481 490
rect 2447 456 2481 462
rect 2447 394 2481 418
rect 2447 384 2481 394
rect 2447 326 2481 346
rect 2447 312 2481 326
rect 2447 258 2481 274
rect 2447 240 2481 258
rect 2447 190 2481 202
rect 2447 168 2481 190
rect 2447 122 2481 130
rect 2447 96 2481 122
rect 2447 54 2481 58
rect 2447 24 2481 54
rect 2447 -48 2481 -14
rect 2447 -116 2481 -86
rect 2447 -120 2481 -116
rect 2447 -184 2481 -158
rect 2447 -192 2481 -184
rect 2447 -252 2481 -230
rect 2447 -264 2481 -252
rect 2447 -320 2481 -302
rect 2447 -336 2481 -320
rect 2447 -388 2481 -374
rect 2447 -408 2481 -388
rect 2447 -456 2481 -446
rect 2447 -480 2481 -456
rect 2447 -524 2481 -518
rect 2447 -552 2481 -524
rect 2447 -592 2481 -590
rect 2447 -624 2481 -592
rect 2447 -694 2481 -662
rect 2447 -696 2481 -694
rect 2447 -762 2481 -734
rect 2447 -768 2481 -762
rect 2755 700 2789 706
rect 2755 672 2789 700
rect 2755 632 2789 634
rect 2755 600 2789 632
rect 2755 530 2789 562
rect 2755 528 2789 530
rect 2755 462 2789 490
rect 2755 456 2789 462
rect 2755 394 2789 418
rect 2755 384 2789 394
rect 2755 326 2789 346
rect 2755 312 2789 326
rect 2755 258 2789 274
rect 2755 240 2789 258
rect 2755 190 2789 202
rect 2755 168 2789 190
rect 2755 122 2789 130
rect 2755 96 2789 122
rect 2755 54 2789 58
rect 2755 24 2789 54
rect 2755 -48 2789 -14
rect 2755 -116 2789 -86
rect 2755 -120 2789 -116
rect 2755 -184 2789 -158
rect 2755 -192 2789 -184
rect 2755 -252 2789 -230
rect 2755 -264 2789 -252
rect 2755 -320 2789 -302
rect 2755 -336 2789 -320
rect 2755 -388 2789 -374
rect 2755 -408 2789 -388
rect 2755 -456 2789 -446
rect 2755 -480 2789 -456
rect 2755 -524 2789 -518
rect 2755 -552 2789 -524
rect 2755 -592 2789 -590
rect 2755 -624 2789 -592
rect 2755 -694 2789 -662
rect 2755 -696 2789 -694
rect 2755 -762 2789 -734
rect 2755 -768 2789 -762
<< metal1 >>
rect -2739 791 -2497 797
rect -2739 757 -2707 791
rect -2673 757 -2635 791
rect -2601 757 -2563 791
rect -2529 757 -2497 791
rect -2739 751 -2497 757
rect -2431 791 -2189 797
rect -2431 757 -2399 791
rect -2365 757 -2327 791
rect -2293 757 -2255 791
rect -2221 757 -2189 791
rect -2431 751 -2189 757
rect -2123 791 -1881 797
rect -2123 757 -2091 791
rect -2057 757 -2019 791
rect -1985 757 -1947 791
rect -1913 757 -1881 791
rect -2123 751 -1881 757
rect -1815 791 -1573 797
rect -1815 757 -1783 791
rect -1749 757 -1711 791
rect -1677 757 -1639 791
rect -1605 757 -1573 791
rect -1815 751 -1573 757
rect -1507 791 -1265 797
rect -1507 757 -1475 791
rect -1441 757 -1403 791
rect -1369 757 -1331 791
rect -1297 757 -1265 791
rect -1507 751 -1265 757
rect -1199 791 -957 797
rect -1199 757 -1167 791
rect -1133 757 -1095 791
rect -1061 757 -1023 791
rect -989 757 -957 791
rect -1199 751 -957 757
rect -891 791 -649 797
rect -891 757 -859 791
rect -825 757 -787 791
rect -753 757 -715 791
rect -681 757 -649 791
rect -891 751 -649 757
rect -583 791 -341 797
rect -583 757 -551 791
rect -517 757 -479 791
rect -445 757 -407 791
rect -373 757 -341 791
rect -583 751 -341 757
rect -275 791 -33 797
rect -275 757 -243 791
rect -209 757 -171 791
rect -137 757 -99 791
rect -65 757 -33 791
rect -275 751 -33 757
rect 33 791 275 797
rect 33 757 65 791
rect 99 757 137 791
rect 171 757 209 791
rect 243 757 275 791
rect 33 751 275 757
rect 341 791 583 797
rect 341 757 373 791
rect 407 757 445 791
rect 479 757 517 791
rect 551 757 583 791
rect 341 751 583 757
rect 649 791 891 797
rect 649 757 681 791
rect 715 757 753 791
rect 787 757 825 791
rect 859 757 891 791
rect 649 751 891 757
rect 957 791 1199 797
rect 957 757 989 791
rect 1023 757 1061 791
rect 1095 757 1133 791
rect 1167 757 1199 791
rect 957 751 1199 757
rect 1265 791 1507 797
rect 1265 757 1297 791
rect 1331 757 1369 791
rect 1403 757 1441 791
rect 1475 757 1507 791
rect 1265 751 1507 757
rect 1573 791 1815 797
rect 1573 757 1605 791
rect 1639 757 1677 791
rect 1711 757 1749 791
rect 1783 757 1815 791
rect 1573 751 1815 757
rect 1881 791 2123 797
rect 1881 757 1913 791
rect 1947 757 1985 791
rect 2019 757 2057 791
rect 2091 757 2123 791
rect 1881 751 2123 757
rect 2189 791 2431 797
rect 2189 757 2221 791
rect 2255 757 2293 791
rect 2327 757 2365 791
rect 2399 757 2431 791
rect 2189 751 2431 757
rect 2497 791 2739 797
rect 2497 757 2529 791
rect 2563 757 2601 791
rect 2635 757 2673 791
rect 2707 757 2739 791
rect 2497 751 2739 757
rect -2795 706 -2749 719
rect -2795 672 -2789 706
rect -2755 672 -2749 706
rect -2795 634 -2749 672
rect -2795 600 -2789 634
rect -2755 600 -2749 634
rect -2795 562 -2749 600
rect -2795 528 -2789 562
rect -2755 528 -2749 562
rect -2795 490 -2749 528
rect -2795 456 -2789 490
rect -2755 456 -2749 490
rect -2795 418 -2749 456
rect -2795 384 -2789 418
rect -2755 384 -2749 418
rect -2795 346 -2749 384
rect -2795 312 -2789 346
rect -2755 312 -2749 346
rect -2795 274 -2749 312
rect -2795 240 -2789 274
rect -2755 240 -2749 274
rect -2795 202 -2749 240
rect -2795 168 -2789 202
rect -2755 168 -2749 202
rect -2795 130 -2749 168
rect -2795 96 -2789 130
rect -2755 96 -2749 130
rect -2795 58 -2749 96
rect -2795 24 -2789 58
rect -2755 24 -2749 58
rect -2795 -14 -2749 24
rect -2795 -48 -2789 -14
rect -2755 -48 -2749 -14
rect -2795 -86 -2749 -48
rect -2795 -120 -2789 -86
rect -2755 -120 -2749 -86
rect -2795 -158 -2749 -120
rect -2795 -192 -2789 -158
rect -2755 -192 -2749 -158
rect -2795 -230 -2749 -192
rect -2795 -264 -2789 -230
rect -2755 -264 -2749 -230
rect -2795 -302 -2749 -264
rect -2795 -336 -2789 -302
rect -2755 -336 -2749 -302
rect -2795 -374 -2749 -336
rect -2795 -408 -2789 -374
rect -2755 -408 -2749 -374
rect -2795 -446 -2749 -408
rect -2795 -480 -2789 -446
rect -2755 -480 -2749 -446
rect -2795 -518 -2749 -480
rect -2795 -552 -2789 -518
rect -2755 -552 -2749 -518
rect -2795 -590 -2749 -552
rect -2795 -624 -2789 -590
rect -2755 -624 -2749 -590
rect -2795 -662 -2749 -624
rect -2795 -696 -2789 -662
rect -2755 -696 -2749 -662
rect -2795 -734 -2749 -696
rect -2795 -768 -2789 -734
rect -2755 -768 -2749 -734
rect -2795 -781 -2749 -768
rect -2487 706 -2441 719
rect -2487 672 -2481 706
rect -2447 672 -2441 706
rect -2487 634 -2441 672
rect -2487 600 -2481 634
rect -2447 600 -2441 634
rect -2487 562 -2441 600
rect -2487 528 -2481 562
rect -2447 528 -2441 562
rect -2487 490 -2441 528
rect -2487 456 -2481 490
rect -2447 456 -2441 490
rect -2487 418 -2441 456
rect -2487 384 -2481 418
rect -2447 384 -2441 418
rect -2487 346 -2441 384
rect -2487 312 -2481 346
rect -2447 312 -2441 346
rect -2487 274 -2441 312
rect -2487 240 -2481 274
rect -2447 240 -2441 274
rect -2487 202 -2441 240
rect -2487 168 -2481 202
rect -2447 168 -2441 202
rect -2487 130 -2441 168
rect -2487 96 -2481 130
rect -2447 96 -2441 130
rect -2487 58 -2441 96
rect -2487 24 -2481 58
rect -2447 24 -2441 58
rect -2487 -14 -2441 24
rect -2487 -48 -2481 -14
rect -2447 -48 -2441 -14
rect -2487 -86 -2441 -48
rect -2487 -120 -2481 -86
rect -2447 -120 -2441 -86
rect -2487 -158 -2441 -120
rect -2487 -192 -2481 -158
rect -2447 -192 -2441 -158
rect -2487 -230 -2441 -192
rect -2487 -264 -2481 -230
rect -2447 -264 -2441 -230
rect -2487 -302 -2441 -264
rect -2487 -336 -2481 -302
rect -2447 -336 -2441 -302
rect -2487 -374 -2441 -336
rect -2487 -408 -2481 -374
rect -2447 -408 -2441 -374
rect -2487 -446 -2441 -408
rect -2487 -480 -2481 -446
rect -2447 -480 -2441 -446
rect -2487 -518 -2441 -480
rect -2487 -552 -2481 -518
rect -2447 -552 -2441 -518
rect -2487 -590 -2441 -552
rect -2487 -624 -2481 -590
rect -2447 -624 -2441 -590
rect -2487 -662 -2441 -624
rect -2487 -696 -2481 -662
rect -2447 -696 -2441 -662
rect -2487 -734 -2441 -696
rect -2487 -768 -2481 -734
rect -2447 -768 -2441 -734
rect -2487 -781 -2441 -768
rect -2179 706 -2133 719
rect -2179 672 -2173 706
rect -2139 672 -2133 706
rect -2179 634 -2133 672
rect -2179 600 -2173 634
rect -2139 600 -2133 634
rect -2179 562 -2133 600
rect -2179 528 -2173 562
rect -2139 528 -2133 562
rect -2179 490 -2133 528
rect -2179 456 -2173 490
rect -2139 456 -2133 490
rect -2179 418 -2133 456
rect -2179 384 -2173 418
rect -2139 384 -2133 418
rect -2179 346 -2133 384
rect -2179 312 -2173 346
rect -2139 312 -2133 346
rect -2179 274 -2133 312
rect -2179 240 -2173 274
rect -2139 240 -2133 274
rect -2179 202 -2133 240
rect -2179 168 -2173 202
rect -2139 168 -2133 202
rect -2179 130 -2133 168
rect -2179 96 -2173 130
rect -2139 96 -2133 130
rect -2179 58 -2133 96
rect -2179 24 -2173 58
rect -2139 24 -2133 58
rect -2179 -14 -2133 24
rect -2179 -48 -2173 -14
rect -2139 -48 -2133 -14
rect -2179 -86 -2133 -48
rect -2179 -120 -2173 -86
rect -2139 -120 -2133 -86
rect -2179 -158 -2133 -120
rect -2179 -192 -2173 -158
rect -2139 -192 -2133 -158
rect -2179 -230 -2133 -192
rect -2179 -264 -2173 -230
rect -2139 -264 -2133 -230
rect -2179 -302 -2133 -264
rect -2179 -336 -2173 -302
rect -2139 -336 -2133 -302
rect -2179 -374 -2133 -336
rect -2179 -408 -2173 -374
rect -2139 -408 -2133 -374
rect -2179 -446 -2133 -408
rect -2179 -480 -2173 -446
rect -2139 -480 -2133 -446
rect -2179 -518 -2133 -480
rect -2179 -552 -2173 -518
rect -2139 -552 -2133 -518
rect -2179 -590 -2133 -552
rect -2179 -624 -2173 -590
rect -2139 -624 -2133 -590
rect -2179 -662 -2133 -624
rect -2179 -696 -2173 -662
rect -2139 -696 -2133 -662
rect -2179 -734 -2133 -696
rect -2179 -768 -2173 -734
rect -2139 -768 -2133 -734
rect -2179 -781 -2133 -768
rect -1871 706 -1825 719
rect -1871 672 -1865 706
rect -1831 672 -1825 706
rect -1871 634 -1825 672
rect -1871 600 -1865 634
rect -1831 600 -1825 634
rect -1871 562 -1825 600
rect -1871 528 -1865 562
rect -1831 528 -1825 562
rect -1871 490 -1825 528
rect -1871 456 -1865 490
rect -1831 456 -1825 490
rect -1871 418 -1825 456
rect -1871 384 -1865 418
rect -1831 384 -1825 418
rect -1871 346 -1825 384
rect -1871 312 -1865 346
rect -1831 312 -1825 346
rect -1871 274 -1825 312
rect -1871 240 -1865 274
rect -1831 240 -1825 274
rect -1871 202 -1825 240
rect -1871 168 -1865 202
rect -1831 168 -1825 202
rect -1871 130 -1825 168
rect -1871 96 -1865 130
rect -1831 96 -1825 130
rect -1871 58 -1825 96
rect -1871 24 -1865 58
rect -1831 24 -1825 58
rect -1871 -14 -1825 24
rect -1871 -48 -1865 -14
rect -1831 -48 -1825 -14
rect -1871 -86 -1825 -48
rect -1871 -120 -1865 -86
rect -1831 -120 -1825 -86
rect -1871 -158 -1825 -120
rect -1871 -192 -1865 -158
rect -1831 -192 -1825 -158
rect -1871 -230 -1825 -192
rect -1871 -264 -1865 -230
rect -1831 -264 -1825 -230
rect -1871 -302 -1825 -264
rect -1871 -336 -1865 -302
rect -1831 -336 -1825 -302
rect -1871 -374 -1825 -336
rect -1871 -408 -1865 -374
rect -1831 -408 -1825 -374
rect -1871 -446 -1825 -408
rect -1871 -480 -1865 -446
rect -1831 -480 -1825 -446
rect -1871 -518 -1825 -480
rect -1871 -552 -1865 -518
rect -1831 -552 -1825 -518
rect -1871 -590 -1825 -552
rect -1871 -624 -1865 -590
rect -1831 -624 -1825 -590
rect -1871 -662 -1825 -624
rect -1871 -696 -1865 -662
rect -1831 -696 -1825 -662
rect -1871 -734 -1825 -696
rect -1871 -768 -1865 -734
rect -1831 -768 -1825 -734
rect -1871 -781 -1825 -768
rect -1563 706 -1517 719
rect -1563 672 -1557 706
rect -1523 672 -1517 706
rect -1563 634 -1517 672
rect -1563 600 -1557 634
rect -1523 600 -1517 634
rect -1563 562 -1517 600
rect -1563 528 -1557 562
rect -1523 528 -1517 562
rect -1563 490 -1517 528
rect -1563 456 -1557 490
rect -1523 456 -1517 490
rect -1563 418 -1517 456
rect -1563 384 -1557 418
rect -1523 384 -1517 418
rect -1563 346 -1517 384
rect -1563 312 -1557 346
rect -1523 312 -1517 346
rect -1563 274 -1517 312
rect -1563 240 -1557 274
rect -1523 240 -1517 274
rect -1563 202 -1517 240
rect -1563 168 -1557 202
rect -1523 168 -1517 202
rect -1563 130 -1517 168
rect -1563 96 -1557 130
rect -1523 96 -1517 130
rect -1563 58 -1517 96
rect -1563 24 -1557 58
rect -1523 24 -1517 58
rect -1563 -14 -1517 24
rect -1563 -48 -1557 -14
rect -1523 -48 -1517 -14
rect -1563 -86 -1517 -48
rect -1563 -120 -1557 -86
rect -1523 -120 -1517 -86
rect -1563 -158 -1517 -120
rect -1563 -192 -1557 -158
rect -1523 -192 -1517 -158
rect -1563 -230 -1517 -192
rect -1563 -264 -1557 -230
rect -1523 -264 -1517 -230
rect -1563 -302 -1517 -264
rect -1563 -336 -1557 -302
rect -1523 -336 -1517 -302
rect -1563 -374 -1517 -336
rect -1563 -408 -1557 -374
rect -1523 -408 -1517 -374
rect -1563 -446 -1517 -408
rect -1563 -480 -1557 -446
rect -1523 -480 -1517 -446
rect -1563 -518 -1517 -480
rect -1563 -552 -1557 -518
rect -1523 -552 -1517 -518
rect -1563 -590 -1517 -552
rect -1563 -624 -1557 -590
rect -1523 -624 -1517 -590
rect -1563 -662 -1517 -624
rect -1563 -696 -1557 -662
rect -1523 -696 -1517 -662
rect -1563 -734 -1517 -696
rect -1563 -768 -1557 -734
rect -1523 -768 -1517 -734
rect -1563 -781 -1517 -768
rect -1255 706 -1209 719
rect -1255 672 -1249 706
rect -1215 672 -1209 706
rect -1255 634 -1209 672
rect -1255 600 -1249 634
rect -1215 600 -1209 634
rect -1255 562 -1209 600
rect -1255 528 -1249 562
rect -1215 528 -1209 562
rect -1255 490 -1209 528
rect -1255 456 -1249 490
rect -1215 456 -1209 490
rect -1255 418 -1209 456
rect -1255 384 -1249 418
rect -1215 384 -1209 418
rect -1255 346 -1209 384
rect -1255 312 -1249 346
rect -1215 312 -1209 346
rect -1255 274 -1209 312
rect -1255 240 -1249 274
rect -1215 240 -1209 274
rect -1255 202 -1209 240
rect -1255 168 -1249 202
rect -1215 168 -1209 202
rect -1255 130 -1209 168
rect -1255 96 -1249 130
rect -1215 96 -1209 130
rect -1255 58 -1209 96
rect -1255 24 -1249 58
rect -1215 24 -1209 58
rect -1255 -14 -1209 24
rect -1255 -48 -1249 -14
rect -1215 -48 -1209 -14
rect -1255 -86 -1209 -48
rect -1255 -120 -1249 -86
rect -1215 -120 -1209 -86
rect -1255 -158 -1209 -120
rect -1255 -192 -1249 -158
rect -1215 -192 -1209 -158
rect -1255 -230 -1209 -192
rect -1255 -264 -1249 -230
rect -1215 -264 -1209 -230
rect -1255 -302 -1209 -264
rect -1255 -336 -1249 -302
rect -1215 -336 -1209 -302
rect -1255 -374 -1209 -336
rect -1255 -408 -1249 -374
rect -1215 -408 -1209 -374
rect -1255 -446 -1209 -408
rect -1255 -480 -1249 -446
rect -1215 -480 -1209 -446
rect -1255 -518 -1209 -480
rect -1255 -552 -1249 -518
rect -1215 -552 -1209 -518
rect -1255 -590 -1209 -552
rect -1255 -624 -1249 -590
rect -1215 -624 -1209 -590
rect -1255 -662 -1209 -624
rect -1255 -696 -1249 -662
rect -1215 -696 -1209 -662
rect -1255 -734 -1209 -696
rect -1255 -768 -1249 -734
rect -1215 -768 -1209 -734
rect -1255 -781 -1209 -768
rect -947 706 -901 719
rect -947 672 -941 706
rect -907 672 -901 706
rect -947 634 -901 672
rect -947 600 -941 634
rect -907 600 -901 634
rect -947 562 -901 600
rect -947 528 -941 562
rect -907 528 -901 562
rect -947 490 -901 528
rect -947 456 -941 490
rect -907 456 -901 490
rect -947 418 -901 456
rect -947 384 -941 418
rect -907 384 -901 418
rect -947 346 -901 384
rect -947 312 -941 346
rect -907 312 -901 346
rect -947 274 -901 312
rect -947 240 -941 274
rect -907 240 -901 274
rect -947 202 -901 240
rect -947 168 -941 202
rect -907 168 -901 202
rect -947 130 -901 168
rect -947 96 -941 130
rect -907 96 -901 130
rect -947 58 -901 96
rect -947 24 -941 58
rect -907 24 -901 58
rect -947 -14 -901 24
rect -947 -48 -941 -14
rect -907 -48 -901 -14
rect -947 -86 -901 -48
rect -947 -120 -941 -86
rect -907 -120 -901 -86
rect -947 -158 -901 -120
rect -947 -192 -941 -158
rect -907 -192 -901 -158
rect -947 -230 -901 -192
rect -947 -264 -941 -230
rect -907 -264 -901 -230
rect -947 -302 -901 -264
rect -947 -336 -941 -302
rect -907 -336 -901 -302
rect -947 -374 -901 -336
rect -947 -408 -941 -374
rect -907 -408 -901 -374
rect -947 -446 -901 -408
rect -947 -480 -941 -446
rect -907 -480 -901 -446
rect -947 -518 -901 -480
rect -947 -552 -941 -518
rect -907 -552 -901 -518
rect -947 -590 -901 -552
rect -947 -624 -941 -590
rect -907 -624 -901 -590
rect -947 -662 -901 -624
rect -947 -696 -941 -662
rect -907 -696 -901 -662
rect -947 -734 -901 -696
rect -947 -768 -941 -734
rect -907 -768 -901 -734
rect -947 -781 -901 -768
rect -639 706 -593 719
rect -639 672 -633 706
rect -599 672 -593 706
rect -639 634 -593 672
rect -639 600 -633 634
rect -599 600 -593 634
rect -639 562 -593 600
rect -639 528 -633 562
rect -599 528 -593 562
rect -639 490 -593 528
rect -639 456 -633 490
rect -599 456 -593 490
rect -639 418 -593 456
rect -639 384 -633 418
rect -599 384 -593 418
rect -639 346 -593 384
rect -639 312 -633 346
rect -599 312 -593 346
rect -639 274 -593 312
rect -639 240 -633 274
rect -599 240 -593 274
rect -639 202 -593 240
rect -639 168 -633 202
rect -599 168 -593 202
rect -639 130 -593 168
rect -639 96 -633 130
rect -599 96 -593 130
rect -639 58 -593 96
rect -639 24 -633 58
rect -599 24 -593 58
rect -639 -14 -593 24
rect -639 -48 -633 -14
rect -599 -48 -593 -14
rect -639 -86 -593 -48
rect -639 -120 -633 -86
rect -599 -120 -593 -86
rect -639 -158 -593 -120
rect -639 -192 -633 -158
rect -599 -192 -593 -158
rect -639 -230 -593 -192
rect -639 -264 -633 -230
rect -599 -264 -593 -230
rect -639 -302 -593 -264
rect -639 -336 -633 -302
rect -599 -336 -593 -302
rect -639 -374 -593 -336
rect -639 -408 -633 -374
rect -599 -408 -593 -374
rect -639 -446 -593 -408
rect -639 -480 -633 -446
rect -599 -480 -593 -446
rect -639 -518 -593 -480
rect -639 -552 -633 -518
rect -599 -552 -593 -518
rect -639 -590 -593 -552
rect -639 -624 -633 -590
rect -599 -624 -593 -590
rect -639 -662 -593 -624
rect -639 -696 -633 -662
rect -599 -696 -593 -662
rect -639 -734 -593 -696
rect -639 -768 -633 -734
rect -599 -768 -593 -734
rect -639 -781 -593 -768
rect -331 706 -285 719
rect -331 672 -325 706
rect -291 672 -285 706
rect -331 634 -285 672
rect -331 600 -325 634
rect -291 600 -285 634
rect -331 562 -285 600
rect -331 528 -325 562
rect -291 528 -285 562
rect -331 490 -285 528
rect -331 456 -325 490
rect -291 456 -285 490
rect -331 418 -285 456
rect -331 384 -325 418
rect -291 384 -285 418
rect -331 346 -285 384
rect -331 312 -325 346
rect -291 312 -285 346
rect -331 274 -285 312
rect -331 240 -325 274
rect -291 240 -285 274
rect -331 202 -285 240
rect -331 168 -325 202
rect -291 168 -285 202
rect -331 130 -285 168
rect -331 96 -325 130
rect -291 96 -285 130
rect -331 58 -285 96
rect -331 24 -325 58
rect -291 24 -285 58
rect -331 -14 -285 24
rect -331 -48 -325 -14
rect -291 -48 -285 -14
rect -331 -86 -285 -48
rect -331 -120 -325 -86
rect -291 -120 -285 -86
rect -331 -158 -285 -120
rect -331 -192 -325 -158
rect -291 -192 -285 -158
rect -331 -230 -285 -192
rect -331 -264 -325 -230
rect -291 -264 -285 -230
rect -331 -302 -285 -264
rect -331 -336 -325 -302
rect -291 -336 -285 -302
rect -331 -374 -285 -336
rect -331 -408 -325 -374
rect -291 -408 -285 -374
rect -331 -446 -285 -408
rect -331 -480 -325 -446
rect -291 -480 -285 -446
rect -331 -518 -285 -480
rect -331 -552 -325 -518
rect -291 -552 -285 -518
rect -331 -590 -285 -552
rect -331 -624 -325 -590
rect -291 -624 -285 -590
rect -331 -662 -285 -624
rect -331 -696 -325 -662
rect -291 -696 -285 -662
rect -331 -734 -285 -696
rect -331 -768 -325 -734
rect -291 -768 -285 -734
rect -331 -781 -285 -768
rect -23 706 23 719
rect -23 672 -17 706
rect 17 672 23 706
rect -23 634 23 672
rect -23 600 -17 634
rect 17 600 23 634
rect -23 562 23 600
rect -23 528 -17 562
rect 17 528 23 562
rect -23 490 23 528
rect -23 456 -17 490
rect 17 456 23 490
rect -23 418 23 456
rect -23 384 -17 418
rect 17 384 23 418
rect -23 346 23 384
rect -23 312 -17 346
rect 17 312 23 346
rect -23 274 23 312
rect -23 240 -17 274
rect 17 240 23 274
rect -23 202 23 240
rect -23 168 -17 202
rect 17 168 23 202
rect -23 130 23 168
rect -23 96 -17 130
rect 17 96 23 130
rect -23 58 23 96
rect -23 24 -17 58
rect 17 24 23 58
rect -23 -14 23 24
rect -23 -48 -17 -14
rect 17 -48 23 -14
rect -23 -86 23 -48
rect -23 -120 -17 -86
rect 17 -120 23 -86
rect -23 -158 23 -120
rect -23 -192 -17 -158
rect 17 -192 23 -158
rect -23 -230 23 -192
rect -23 -264 -17 -230
rect 17 -264 23 -230
rect -23 -302 23 -264
rect -23 -336 -17 -302
rect 17 -336 23 -302
rect -23 -374 23 -336
rect -23 -408 -17 -374
rect 17 -408 23 -374
rect -23 -446 23 -408
rect -23 -480 -17 -446
rect 17 -480 23 -446
rect -23 -518 23 -480
rect -23 -552 -17 -518
rect 17 -552 23 -518
rect -23 -590 23 -552
rect -23 -624 -17 -590
rect 17 -624 23 -590
rect -23 -662 23 -624
rect -23 -696 -17 -662
rect 17 -696 23 -662
rect -23 -734 23 -696
rect -23 -768 -17 -734
rect 17 -768 23 -734
rect -23 -781 23 -768
rect 285 706 331 719
rect 285 672 291 706
rect 325 672 331 706
rect 285 634 331 672
rect 285 600 291 634
rect 325 600 331 634
rect 285 562 331 600
rect 285 528 291 562
rect 325 528 331 562
rect 285 490 331 528
rect 285 456 291 490
rect 325 456 331 490
rect 285 418 331 456
rect 285 384 291 418
rect 325 384 331 418
rect 285 346 331 384
rect 285 312 291 346
rect 325 312 331 346
rect 285 274 331 312
rect 285 240 291 274
rect 325 240 331 274
rect 285 202 331 240
rect 285 168 291 202
rect 325 168 331 202
rect 285 130 331 168
rect 285 96 291 130
rect 325 96 331 130
rect 285 58 331 96
rect 285 24 291 58
rect 325 24 331 58
rect 285 -14 331 24
rect 285 -48 291 -14
rect 325 -48 331 -14
rect 285 -86 331 -48
rect 285 -120 291 -86
rect 325 -120 331 -86
rect 285 -158 331 -120
rect 285 -192 291 -158
rect 325 -192 331 -158
rect 285 -230 331 -192
rect 285 -264 291 -230
rect 325 -264 331 -230
rect 285 -302 331 -264
rect 285 -336 291 -302
rect 325 -336 331 -302
rect 285 -374 331 -336
rect 285 -408 291 -374
rect 325 -408 331 -374
rect 285 -446 331 -408
rect 285 -480 291 -446
rect 325 -480 331 -446
rect 285 -518 331 -480
rect 285 -552 291 -518
rect 325 -552 331 -518
rect 285 -590 331 -552
rect 285 -624 291 -590
rect 325 -624 331 -590
rect 285 -662 331 -624
rect 285 -696 291 -662
rect 325 -696 331 -662
rect 285 -734 331 -696
rect 285 -768 291 -734
rect 325 -768 331 -734
rect 285 -781 331 -768
rect 593 706 639 719
rect 593 672 599 706
rect 633 672 639 706
rect 593 634 639 672
rect 593 600 599 634
rect 633 600 639 634
rect 593 562 639 600
rect 593 528 599 562
rect 633 528 639 562
rect 593 490 639 528
rect 593 456 599 490
rect 633 456 639 490
rect 593 418 639 456
rect 593 384 599 418
rect 633 384 639 418
rect 593 346 639 384
rect 593 312 599 346
rect 633 312 639 346
rect 593 274 639 312
rect 593 240 599 274
rect 633 240 639 274
rect 593 202 639 240
rect 593 168 599 202
rect 633 168 639 202
rect 593 130 639 168
rect 593 96 599 130
rect 633 96 639 130
rect 593 58 639 96
rect 593 24 599 58
rect 633 24 639 58
rect 593 -14 639 24
rect 593 -48 599 -14
rect 633 -48 639 -14
rect 593 -86 639 -48
rect 593 -120 599 -86
rect 633 -120 639 -86
rect 593 -158 639 -120
rect 593 -192 599 -158
rect 633 -192 639 -158
rect 593 -230 639 -192
rect 593 -264 599 -230
rect 633 -264 639 -230
rect 593 -302 639 -264
rect 593 -336 599 -302
rect 633 -336 639 -302
rect 593 -374 639 -336
rect 593 -408 599 -374
rect 633 -408 639 -374
rect 593 -446 639 -408
rect 593 -480 599 -446
rect 633 -480 639 -446
rect 593 -518 639 -480
rect 593 -552 599 -518
rect 633 -552 639 -518
rect 593 -590 639 -552
rect 593 -624 599 -590
rect 633 -624 639 -590
rect 593 -662 639 -624
rect 593 -696 599 -662
rect 633 -696 639 -662
rect 593 -734 639 -696
rect 593 -768 599 -734
rect 633 -768 639 -734
rect 593 -781 639 -768
rect 901 706 947 719
rect 901 672 907 706
rect 941 672 947 706
rect 901 634 947 672
rect 901 600 907 634
rect 941 600 947 634
rect 901 562 947 600
rect 901 528 907 562
rect 941 528 947 562
rect 901 490 947 528
rect 901 456 907 490
rect 941 456 947 490
rect 901 418 947 456
rect 901 384 907 418
rect 941 384 947 418
rect 901 346 947 384
rect 901 312 907 346
rect 941 312 947 346
rect 901 274 947 312
rect 901 240 907 274
rect 941 240 947 274
rect 901 202 947 240
rect 901 168 907 202
rect 941 168 947 202
rect 901 130 947 168
rect 901 96 907 130
rect 941 96 947 130
rect 901 58 947 96
rect 901 24 907 58
rect 941 24 947 58
rect 901 -14 947 24
rect 901 -48 907 -14
rect 941 -48 947 -14
rect 901 -86 947 -48
rect 901 -120 907 -86
rect 941 -120 947 -86
rect 901 -158 947 -120
rect 901 -192 907 -158
rect 941 -192 947 -158
rect 901 -230 947 -192
rect 901 -264 907 -230
rect 941 -264 947 -230
rect 901 -302 947 -264
rect 901 -336 907 -302
rect 941 -336 947 -302
rect 901 -374 947 -336
rect 901 -408 907 -374
rect 941 -408 947 -374
rect 901 -446 947 -408
rect 901 -480 907 -446
rect 941 -480 947 -446
rect 901 -518 947 -480
rect 901 -552 907 -518
rect 941 -552 947 -518
rect 901 -590 947 -552
rect 901 -624 907 -590
rect 941 -624 947 -590
rect 901 -662 947 -624
rect 901 -696 907 -662
rect 941 -696 947 -662
rect 901 -734 947 -696
rect 901 -768 907 -734
rect 941 -768 947 -734
rect 901 -781 947 -768
rect 1209 706 1255 719
rect 1209 672 1215 706
rect 1249 672 1255 706
rect 1209 634 1255 672
rect 1209 600 1215 634
rect 1249 600 1255 634
rect 1209 562 1255 600
rect 1209 528 1215 562
rect 1249 528 1255 562
rect 1209 490 1255 528
rect 1209 456 1215 490
rect 1249 456 1255 490
rect 1209 418 1255 456
rect 1209 384 1215 418
rect 1249 384 1255 418
rect 1209 346 1255 384
rect 1209 312 1215 346
rect 1249 312 1255 346
rect 1209 274 1255 312
rect 1209 240 1215 274
rect 1249 240 1255 274
rect 1209 202 1255 240
rect 1209 168 1215 202
rect 1249 168 1255 202
rect 1209 130 1255 168
rect 1209 96 1215 130
rect 1249 96 1255 130
rect 1209 58 1255 96
rect 1209 24 1215 58
rect 1249 24 1255 58
rect 1209 -14 1255 24
rect 1209 -48 1215 -14
rect 1249 -48 1255 -14
rect 1209 -86 1255 -48
rect 1209 -120 1215 -86
rect 1249 -120 1255 -86
rect 1209 -158 1255 -120
rect 1209 -192 1215 -158
rect 1249 -192 1255 -158
rect 1209 -230 1255 -192
rect 1209 -264 1215 -230
rect 1249 -264 1255 -230
rect 1209 -302 1255 -264
rect 1209 -336 1215 -302
rect 1249 -336 1255 -302
rect 1209 -374 1255 -336
rect 1209 -408 1215 -374
rect 1249 -408 1255 -374
rect 1209 -446 1255 -408
rect 1209 -480 1215 -446
rect 1249 -480 1255 -446
rect 1209 -518 1255 -480
rect 1209 -552 1215 -518
rect 1249 -552 1255 -518
rect 1209 -590 1255 -552
rect 1209 -624 1215 -590
rect 1249 -624 1255 -590
rect 1209 -662 1255 -624
rect 1209 -696 1215 -662
rect 1249 -696 1255 -662
rect 1209 -734 1255 -696
rect 1209 -768 1215 -734
rect 1249 -768 1255 -734
rect 1209 -781 1255 -768
rect 1517 706 1563 719
rect 1517 672 1523 706
rect 1557 672 1563 706
rect 1517 634 1563 672
rect 1517 600 1523 634
rect 1557 600 1563 634
rect 1517 562 1563 600
rect 1517 528 1523 562
rect 1557 528 1563 562
rect 1517 490 1563 528
rect 1517 456 1523 490
rect 1557 456 1563 490
rect 1517 418 1563 456
rect 1517 384 1523 418
rect 1557 384 1563 418
rect 1517 346 1563 384
rect 1517 312 1523 346
rect 1557 312 1563 346
rect 1517 274 1563 312
rect 1517 240 1523 274
rect 1557 240 1563 274
rect 1517 202 1563 240
rect 1517 168 1523 202
rect 1557 168 1563 202
rect 1517 130 1563 168
rect 1517 96 1523 130
rect 1557 96 1563 130
rect 1517 58 1563 96
rect 1517 24 1523 58
rect 1557 24 1563 58
rect 1517 -14 1563 24
rect 1517 -48 1523 -14
rect 1557 -48 1563 -14
rect 1517 -86 1563 -48
rect 1517 -120 1523 -86
rect 1557 -120 1563 -86
rect 1517 -158 1563 -120
rect 1517 -192 1523 -158
rect 1557 -192 1563 -158
rect 1517 -230 1563 -192
rect 1517 -264 1523 -230
rect 1557 -264 1563 -230
rect 1517 -302 1563 -264
rect 1517 -336 1523 -302
rect 1557 -336 1563 -302
rect 1517 -374 1563 -336
rect 1517 -408 1523 -374
rect 1557 -408 1563 -374
rect 1517 -446 1563 -408
rect 1517 -480 1523 -446
rect 1557 -480 1563 -446
rect 1517 -518 1563 -480
rect 1517 -552 1523 -518
rect 1557 -552 1563 -518
rect 1517 -590 1563 -552
rect 1517 -624 1523 -590
rect 1557 -624 1563 -590
rect 1517 -662 1563 -624
rect 1517 -696 1523 -662
rect 1557 -696 1563 -662
rect 1517 -734 1563 -696
rect 1517 -768 1523 -734
rect 1557 -768 1563 -734
rect 1517 -781 1563 -768
rect 1825 706 1871 719
rect 1825 672 1831 706
rect 1865 672 1871 706
rect 1825 634 1871 672
rect 1825 600 1831 634
rect 1865 600 1871 634
rect 1825 562 1871 600
rect 1825 528 1831 562
rect 1865 528 1871 562
rect 1825 490 1871 528
rect 1825 456 1831 490
rect 1865 456 1871 490
rect 1825 418 1871 456
rect 1825 384 1831 418
rect 1865 384 1871 418
rect 1825 346 1871 384
rect 1825 312 1831 346
rect 1865 312 1871 346
rect 1825 274 1871 312
rect 1825 240 1831 274
rect 1865 240 1871 274
rect 1825 202 1871 240
rect 1825 168 1831 202
rect 1865 168 1871 202
rect 1825 130 1871 168
rect 1825 96 1831 130
rect 1865 96 1871 130
rect 1825 58 1871 96
rect 1825 24 1831 58
rect 1865 24 1871 58
rect 1825 -14 1871 24
rect 1825 -48 1831 -14
rect 1865 -48 1871 -14
rect 1825 -86 1871 -48
rect 1825 -120 1831 -86
rect 1865 -120 1871 -86
rect 1825 -158 1871 -120
rect 1825 -192 1831 -158
rect 1865 -192 1871 -158
rect 1825 -230 1871 -192
rect 1825 -264 1831 -230
rect 1865 -264 1871 -230
rect 1825 -302 1871 -264
rect 1825 -336 1831 -302
rect 1865 -336 1871 -302
rect 1825 -374 1871 -336
rect 1825 -408 1831 -374
rect 1865 -408 1871 -374
rect 1825 -446 1871 -408
rect 1825 -480 1831 -446
rect 1865 -480 1871 -446
rect 1825 -518 1871 -480
rect 1825 -552 1831 -518
rect 1865 -552 1871 -518
rect 1825 -590 1871 -552
rect 1825 -624 1831 -590
rect 1865 -624 1871 -590
rect 1825 -662 1871 -624
rect 1825 -696 1831 -662
rect 1865 -696 1871 -662
rect 1825 -734 1871 -696
rect 1825 -768 1831 -734
rect 1865 -768 1871 -734
rect 1825 -781 1871 -768
rect 2133 706 2179 719
rect 2133 672 2139 706
rect 2173 672 2179 706
rect 2133 634 2179 672
rect 2133 600 2139 634
rect 2173 600 2179 634
rect 2133 562 2179 600
rect 2133 528 2139 562
rect 2173 528 2179 562
rect 2133 490 2179 528
rect 2133 456 2139 490
rect 2173 456 2179 490
rect 2133 418 2179 456
rect 2133 384 2139 418
rect 2173 384 2179 418
rect 2133 346 2179 384
rect 2133 312 2139 346
rect 2173 312 2179 346
rect 2133 274 2179 312
rect 2133 240 2139 274
rect 2173 240 2179 274
rect 2133 202 2179 240
rect 2133 168 2139 202
rect 2173 168 2179 202
rect 2133 130 2179 168
rect 2133 96 2139 130
rect 2173 96 2179 130
rect 2133 58 2179 96
rect 2133 24 2139 58
rect 2173 24 2179 58
rect 2133 -14 2179 24
rect 2133 -48 2139 -14
rect 2173 -48 2179 -14
rect 2133 -86 2179 -48
rect 2133 -120 2139 -86
rect 2173 -120 2179 -86
rect 2133 -158 2179 -120
rect 2133 -192 2139 -158
rect 2173 -192 2179 -158
rect 2133 -230 2179 -192
rect 2133 -264 2139 -230
rect 2173 -264 2179 -230
rect 2133 -302 2179 -264
rect 2133 -336 2139 -302
rect 2173 -336 2179 -302
rect 2133 -374 2179 -336
rect 2133 -408 2139 -374
rect 2173 -408 2179 -374
rect 2133 -446 2179 -408
rect 2133 -480 2139 -446
rect 2173 -480 2179 -446
rect 2133 -518 2179 -480
rect 2133 -552 2139 -518
rect 2173 -552 2179 -518
rect 2133 -590 2179 -552
rect 2133 -624 2139 -590
rect 2173 -624 2179 -590
rect 2133 -662 2179 -624
rect 2133 -696 2139 -662
rect 2173 -696 2179 -662
rect 2133 -734 2179 -696
rect 2133 -768 2139 -734
rect 2173 -768 2179 -734
rect 2133 -781 2179 -768
rect 2441 706 2487 719
rect 2441 672 2447 706
rect 2481 672 2487 706
rect 2441 634 2487 672
rect 2441 600 2447 634
rect 2481 600 2487 634
rect 2441 562 2487 600
rect 2441 528 2447 562
rect 2481 528 2487 562
rect 2441 490 2487 528
rect 2441 456 2447 490
rect 2481 456 2487 490
rect 2441 418 2487 456
rect 2441 384 2447 418
rect 2481 384 2487 418
rect 2441 346 2487 384
rect 2441 312 2447 346
rect 2481 312 2487 346
rect 2441 274 2487 312
rect 2441 240 2447 274
rect 2481 240 2487 274
rect 2441 202 2487 240
rect 2441 168 2447 202
rect 2481 168 2487 202
rect 2441 130 2487 168
rect 2441 96 2447 130
rect 2481 96 2487 130
rect 2441 58 2487 96
rect 2441 24 2447 58
rect 2481 24 2487 58
rect 2441 -14 2487 24
rect 2441 -48 2447 -14
rect 2481 -48 2487 -14
rect 2441 -86 2487 -48
rect 2441 -120 2447 -86
rect 2481 -120 2487 -86
rect 2441 -158 2487 -120
rect 2441 -192 2447 -158
rect 2481 -192 2487 -158
rect 2441 -230 2487 -192
rect 2441 -264 2447 -230
rect 2481 -264 2487 -230
rect 2441 -302 2487 -264
rect 2441 -336 2447 -302
rect 2481 -336 2487 -302
rect 2441 -374 2487 -336
rect 2441 -408 2447 -374
rect 2481 -408 2487 -374
rect 2441 -446 2487 -408
rect 2441 -480 2447 -446
rect 2481 -480 2487 -446
rect 2441 -518 2487 -480
rect 2441 -552 2447 -518
rect 2481 -552 2487 -518
rect 2441 -590 2487 -552
rect 2441 -624 2447 -590
rect 2481 -624 2487 -590
rect 2441 -662 2487 -624
rect 2441 -696 2447 -662
rect 2481 -696 2487 -662
rect 2441 -734 2487 -696
rect 2441 -768 2447 -734
rect 2481 -768 2487 -734
rect 2441 -781 2487 -768
rect 2749 706 2795 719
rect 2749 672 2755 706
rect 2789 672 2795 706
rect 2749 634 2795 672
rect 2749 600 2755 634
rect 2789 600 2795 634
rect 2749 562 2795 600
rect 2749 528 2755 562
rect 2789 528 2795 562
rect 2749 490 2795 528
rect 2749 456 2755 490
rect 2789 456 2795 490
rect 2749 418 2795 456
rect 2749 384 2755 418
rect 2789 384 2795 418
rect 2749 346 2795 384
rect 2749 312 2755 346
rect 2789 312 2795 346
rect 2749 274 2795 312
rect 2749 240 2755 274
rect 2789 240 2795 274
rect 2749 202 2795 240
rect 2749 168 2755 202
rect 2789 168 2795 202
rect 2749 130 2795 168
rect 2749 96 2755 130
rect 2789 96 2795 130
rect 2749 58 2795 96
rect 2749 24 2755 58
rect 2789 24 2795 58
rect 2749 -14 2795 24
rect 2749 -48 2755 -14
rect 2789 -48 2795 -14
rect 2749 -86 2795 -48
rect 2749 -120 2755 -86
rect 2789 -120 2795 -86
rect 2749 -158 2795 -120
rect 2749 -192 2755 -158
rect 2789 -192 2795 -158
rect 2749 -230 2795 -192
rect 2749 -264 2755 -230
rect 2789 -264 2795 -230
rect 2749 -302 2795 -264
rect 2749 -336 2755 -302
rect 2789 -336 2795 -302
rect 2749 -374 2795 -336
rect 2749 -408 2755 -374
rect 2789 -408 2795 -374
rect 2749 -446 2795 -408
rect 2749 -480 2755 -446
rect 2789 -480 2795 -446
rect 2749 -518 2795 -480
rect 2749 -552 2755 -518
rect 2789 -552 2795 -518
rect 2749 -590 2795 -552
rect 2749 -624 2755 -590
rect 2789 -624 2795 -590
rect 2749 -662 2795 -624
rect 2749 -696 2755 -662
rect 2789 -696 2795 -662
rect 2749 -734 2795 -696
rect 2749 -768 2755 -734
rect 2789 -768 2795 -734
rect 2749 -781 2795 -768
<< end >>
