magic
tech sky130A
magscale 1 2
timestamp 1770083657
<< pwell >>
rect 2074 974 8126 1126
rect 2074 -774 2226 974
rect 7974 -774 8126 974
rect 2074 -926 8126 -774
<< psubdiff >>
rect 2100 1067 8100 1100
rect 2100 1033 2227 1067
rect 2261 1033 2295 1067
rect 2329 1033 2363 1067
rect 2397 1033 2431 1067
rect 2465 1033 2499 1067
rect 2533 1033 2567 1067
rect 2601 1033 2635 1067
rect 2669 1033 2703 1067
rect 2737 1033 2771 1067
rect 2805 1033 2839 1067
rect 2873 1033 2907 1067
rect 2941 1033 2975 1067
rect 3009 1033 3043 1067
rect 3077 1033 3111 1067
rect 3145 1033 3179 1067
rect 3213 1033 3247 1067
rect 3281 1033 3315 1067
rect 3349 1033 3383 1067
rect 3417 1033 3451 1067
rect 3485 1033 3519 1067
rect 3553 1033 3587 1067
rect 3621 1033 3655 1067
rect 3689 1033 3723 1067
rect 3757 1033 3791 1067
rect 3825 1033 3859 1067
rect 3893 1033 3927 1067
rect 3961 1033 3995 1067
rect 4029 1033 4063 1067
rect 4097 1033 4131 1067
rect 4165 1033 4199 1067
rect 4233 1033 4267 1067
rect 4301 1033 4335 1067
rect 4369 1033 4403 1067
rect 4437 1033 4471 1067
rect 4505 1033 4539 1067
rect 4573 1033 4607 1067
rect 4641 1033 4675 1067
rect 4709 1033 4743 1067
rect 4777 1033 4811 1067
rect 4845 1033 4879 1067
rect 4913 1033 4947 1067
rect 4981 1033 5015 1067
rect 5049 1033 5083 1067
rect 5117 1033 5151 1067
rect 5185 1033 5219 1067
rect 5253 1033 5287 1067
rect 5321 1033 5355 1067
rect 5389 1033 5423 1067
rect 5457 1033 5491 1067
rect 5525 1033 5559 1067
rect 5593 1033 5627 1067
rect 5661 1033 5695 1067
rect 5729 1033 5763 1067
rect 5797 1033 5831 1067
rect 5865 1033 5899 1067
rect 5933 1033 5967 1067
rect 6001 1033 6035 1067
rect 6069 1033 6103 1067
rect 6137 1033 6171 1067
rect 6205 1033 6239 1067
rect 6273 1033 6307 1067
rect 6341 1033 6375 1067
rect 6409 1033 6443 1067
rect 6477 1033 6511 1067
rect 6545 1033 6579 1067
rect 6613 1033 6647 1067
rect 6681 1033 6715 1067
rect 6749 1033 6783 1067
rect 6817 1033 6851 1067
rect 6885 1033 6919 1067
rect 6953 1033 6987 1067
rect 7021 1033 7055 1067
rect 7089 1033 7123 1067
rect 7157 1033 7191 1067
rect 7225 1033 7259 1067
rect 7293 1033 7327 1067
rect 7361 1033 7395 1067
rect 7429 1033 7463 1067
rect 7497 1033 7531 1067
rect 7565 1033 7599 1067
rect 7633 1033 7667 1067
rect 7701 1033 7735 1067
rect 7769 1033 7803 1067
rect 7837 1033 7871 1067
rect 7905 1033 7939 1067
rect 7973 1033 8100 1067
rect 2100 1000 8100 1033
rect 2100 967 2200 1000
rect 2100 933 2133 967
rect 2167 933 2200 967
rect 2100 899 2200 933
rect 2100 865 2133 899
rect 2167 865 2200 899
rect 2100 831 2200 865
rect 2100 797 2133 831
rect 2167 797 2200 831
rect 2100 763 2200 797
rect 2100 729 2133 763
rect 2167 729 2200 763
rect 2100 695 2200 729
rect 2100 661 2133 695
rect 2167 661 2200 695
rect 2100 627 2200 661
rect 2100 593 2133 627
rect 2167 593 2200 627
rect 2100 559 2200 593
rect 2100 525 2133 559
rect 2167 525 2200 559
rect 2100 491 2200 525
rect 2100 457 2133 491
rect 2167 457 2200 491
rect 2100 423 2200 457
rect 2100 389 2133 423
rect 2167 389 2200 423
rect 2100 355 2200 389
rect 2100 321 2133 355
rect 2167 321 2200 355
rect 2100 287 2200 321
rect 2100 253 2133 287
rect 2167 253 2200 287
rect 2100 219 2200 253
rect 2100 185 2133 219
rect 2167 185 2200 219
rect 2100 151 2200 185
rect 2100 117 2133 151
rect 2167 117 2200 151
rect 2100 83 2200 117
rect 2100 49 2133 83
rect 2167 49 2200 83
rect 2100 15 2200 49
rect 2100 -19 2133 15
rect 2167 -19 2200 15
rect 2100 -53 2200 -19
rect 2100 -87 2133 -53
rect 2167 -87 2200 -53
rect 2100 -121 2200 -87
rect 2100 -155 2133 -121
rect 2167 -155 2200 -121
rect 2100 -189 2200 -155
rect 2100 -223 2133 -189
rect 2167 -223 2200 -189
rect 2100 -257 2200 -223
rect 2100 -291 2133 -257
rect 2167 -291 2200 -257
rect 2100 -325 2200 -291
rect 2100 -359 2133 -325
rect 2167 -359 2200 -325
rect 2100 -393 2200 -359
rect 2100 -427 2133 -393
rect 2167 -427 2200 -393
rect 2100 -461 2200 -427
rect 2100 -495 2133 -461
rect 2167 -495 2200 -461
rect 2100 -529 2200 -495
rect 2100 -563 2133 -529
rect 2167 -563 2200 -529
rect 2100 -597 2200 -563
rect 2100 -631 2133 -597
rect 2167 -631 2200 -597
rect 2100 -665 2200 -631
rect 2100 -699 2133 -665
rect 2167 -699 2200 -665
rect 2100 -733 2200 -699
rect 2100 -767 2133 -733
rect 2167 -767 2200 -733
rect 2100 -800 2200 -767
rect 8000 967 8100 1000
rect 8000 933 8033 967
rect 8067 933 8100 967
rect 8000 899 8100 933
rect 8000 865 8033 899
rect 8067 865 8100 899
rect 8000 831 8100 865
rect 8000 797 8033 831
rect 8067 797 8100 831
rect 8000 763 8100 797
rect 8000 729 8033 763
rect 8067 729 8100 763
rect 8000 695 8100 729
rect 8000 661 8033 695
rect 8067 661 8100 695
rect 8000 627 8100 661
rect 8000 593 8033 627
rect 8067 593 8100 627
rect 8000 559 8100 593
rect 8000 525 8033 559
rect 8067 525 8100 559
rect 8000 491 8100 525
rect 8000 457 8033 491
rect 8067 457 8100 491
rect 8000 423 8100 457
rect 8000 389 8033 423
rect 8067 389 8100 423
rect 8000 355 8100 389
rect 8000 321 8033 355
rect 8067 321 8100 355
rect 8000 287 8100 321
rect 8000 253 8033 287
rect 8067 253 8100 287
rect 8000 219 8100 253
rect 8000 185 8033 219
rect 8067 185 8100 219
rect 8000 151 8100 185
rect 8000 117 8033 151
rect 8067 117 8100 151
rect 8000 83 8100 117
rect 8000 49 8033 83
rect 8067 49 8100 83
rect 8000 15 8100 49
rect 8000 -19 8033 15
rect 8067 -19 8100 15
rect 8000 -53 8100 -19
rect 8000 -87 8033 -53
rect 8067 -87 8100 -53
rect 8000 -121 8100 -87
rect 8000 -155 8033 -121
rect 8067 -155 8100 -121
rect 8000 -189 8100 -155
rect 8000 -223 8033 -189
rect 8067 -223 8100 -189
rect 8000 -257 8100 -223
rect 8000 -291 8033 -257
rect 8067 -291 8100 -257
rect 8000 -325 8100 -291
rect 8000 -359 8033 -325
rect 8067 -359 8100 -325
rect 8000 -393 8100 -359
rect 8000 -427 8033 -393
rect 8067 -427 8100 -393
rect 8000 -461 8100 -427
rect 8000 -495 8033 -461
rect 8067 -495 8100 -461
rect 8000 -529 8100 -495
rect 8000 -563 8033 -529
rect 8067 -563 8100 -529
rect 8000 -597 8100 -563
rect 8000 -631 8033 -597
rect 8067 -631 8100 -597
rect 8000 -665 8100 -631
rect 8000 -699 8033 -665
rect 8067 -699 8100 -665
rect 8000 -733 8100 -699
rect 8000 -767 8033 -733
rect 8067 -767 8100 -733
rect 8000 -800 8100 -767
rect 2100 -833 8100 -800
rect 2100 -867 2227 -833
rect 2261 -867 2295 -833
rect 2329 -867 2363 -833
rect 2397 -867 2431 -833
rect 2465 -867 2499 -833
rect 2533 -867 2567 -833
rect 2601 -867 2635 -833
rect 2669 -867 2703 -833
rect 2737 -867 2771 -833
rect 2805 -867 2839 -833
rect 2873 -867 2907 -833
rect 2941 -867 2975 -833
rect 3009 -867 3043 -833
rect 3077 -867 3111 -833
rect 3145 -867 3179 -833
rect 3213 -867 3247 -833
rect 3281 -867 3315 -833
rect 3349 -867 3383 -833
rect 3417 -867 3451 -833
rect 3485 -867 3519 -833
rect 3553 -867 3587 -833
rect 3621 -867 3655 -833
rect 3689 -867 3723 -833
rect 3757 -867 3791 -833
rect 3825 -867 3859 -833
rect 3893 -867 3927 -833
rect 3961 -867 3995 -833
rect 4029 -867 4063 -833
rect 4097 -867 4131 -833
rect 4165 -867 4199 -833
rect 4233 -867 4267 -833
rect 4301 -867 4335 -833
rect 4369 -867 4403 -833
rect 4437 -867 4471 -833
rect 4505 -867 4539 -833
rect 4573 -867 4607 -833
rect 4641 -867 4675 -833
rect 4709 -867 4743 -833
rect 4777 -867 4811 -833
rect 4845 -867 4879 -833
rect 4913 -867 4947 -833
rect 4981 -867 5015 -833
rect 5049 -867 5083 -833
rect 5117 -867 5151 -833
rect 5185 -867 5219 -833
rect 5253 -867 5287 -833
rect 5321 -867 5355 -833
rect 5389 -867 5423 -833
rect 5457 -867 5491 -833
rect 5525 -867 5559 -833
rect 5593 -867 5627 -833
rect 5661 -867 5695 -833
rect 5729 -867 5763 -833
rect 5797 -867 5831 -833
rect 5865 -867 5899 -833
rect 5933 -867 5967 -833
rect 6001 -867 6035 -833
rect 6069 -867 6103 -833
rect 6137 -867 6171 -833
rect 6205 -867 6239 -833
rect 6273 -867 6307 -833
rect 6341 -867 6375 -833
rect 6409 -867 6443 -833
rect 6477 -867 6511 -833
rect 6545 -867 6579 -833
rect 6613 -867 6647 -833
rect 6681 -867 6715 -833
rect 6749 -867 6783 -833
rect 6817 -867 6851 -833
rect 6885 -867 6919 -833
rect 6953 -867 6987 -833
rect 7021 -867 7055 -833
rect 7089 -867 7123 -833
rect 7157 -867 7191 -833
rect 7225 -867 7259 -833
rect 7293 -867 7327 -833
rect 7361 -867 7395 -833
rect 7429 -867 7463 -833
rect 7497 -867 7531 -833
rect 7565 -867 7599 -833
rect 7633 -867 7667 -833
rect 7701 -867 7735 -833
rect 7769 -867 7803 -833
rect 7837 -867 7871 -833
rect 7905 -867 7939 -833
rect 7973 -867 8100 -833
rect 2100 -900 8100 -867
<< psubdiffcont >>
rect 2227 1033 2261 1067
rect 2295 1033 2329 1067
rect 2363 1033 2397 1067
rect 2431 1033 2465 1067
rect 2499 1033 2533 1067
rect 2567 1033 2601 1067
rect 2635 1033 2669 1067
rect 2703 1033 2737 1067
rect 2771 1033 2805 1067
rect 2839 1033 2873 1067
rect 2907 1033 2941 1067
rect 2975 1033 3009 1067
rect 3043 1033 3077 1067
rect 3111 1033 3145 1067
rect 3179 1033 3213 1067
rect 3247 1033 3281 1067
rect 3315 1033 3349 1067
rect 3383 1033 3417 1067
rect 3451 1033 3485 1067
rect 3519 1033 3553 1067
rect 3587 1033 3621 1067
rect 3655 1033 3689 1067
rect 3723 1033 3757 1067
rect 3791 1033 3825 1067
rect 3859 1033 3893 1067
rect 3927 1033 3961 1067
rect 3995 1033 4029 1067
rect 4063 1033 4097 1067
rect 4131 1033 4165 1067
rect 4199 1033 4233 1067
rect 4267 1033 4301 1067
rect 4335 1033 4369 1067
rect 4403 1033 4437 1067
rect 4471 1033 4505 1067
rect 4539 1033 4573 1067
rect 4607 1033 4641 1067
rect 4675 1033 4709 1067
rect 4743 1033 4777 1067
rect 4811 1033 4845 1067
rect 4879 1033 4913 1067
rect 4947 1033 4981 1067
rect 5015 1033 5049 1067
rect 5083 1033 5117 1067
rect 5151 1033 5185 1067
rect 5219 1033 5253 1067
rect 5287 1033 5321 1067
rect 5355 1033 5389 1067
rect 5423 1033 5457 1067
rect 5491 1033 5525 1067
rect 5559 1033 5593 1067
rect 5627 1033 5661 1067
rect 5695 1033 5729 1067
rect 5763 1033 5797 1067
rect 5831 1033 5865 1067
rect 5899 1033 5933 1067
rect 5967 1033 6001 1067
rect 6035 1033 6069 1067
rect 6103 1033 6137 1067
rect 6171 1033 6205 1067
rect 6239 1033 6273 1067
rect 6307 1033 6341 1067
rect 6375 1033 6409 1067
rect 6443 1033 6477 1067
rect 6511 1033 6545 1067
rect 6579 1033 6613 1067
rect 6647 1033 6681 1067
rect 6715 1033 6749 1067
rect 6783 1033 6817 1067
rect 6851 1033 6885 1067
rect 6919 1033 6953 1067
rect 6987 1033 7021 1067
rect 7055 1033 7089 1067
rect 7123 1033 7157 1067
rect 7191 1033 7225 1067
rect 7259 1033 7293 1067
rect 7327 1033 7361 1067
rect 7395 1033 7429 1067
rect 7463 1033 7497 1067
rect 7531 1033 7565 1067
rect 7599 1033 7633 1067
rect 7667 1033 7701 1067
rect 7735 1033 7769 1067
rect 7803 1033 7837 1067
rect 7871 1033 7905 1067
rect 7939 1033 7973 1067
rect 2133 933 2167 967
rect 2133 865 2167 899
rect 2133 797 2167 831
rect 2133 729 2167 763
rect 2133 661 2167 695
rect 2133 593 2167 627
rect 2133 525 2167 559
rect 2133 457 2167 491
rect 2133 389 2167 423
rect 2133 321 2167 355
rect 2133 253 2167 287
rect 2133 185 2167 219
rect 2133 117 2167 151
rect 2133 49 2167 83
rect 2133 -19 2167 15
rect 2133 -87 2167 -53
rect 2133 -155 2167 -121
rect 2133 -223 2167 -189
rect 2133 -291 2167 -257
rect 2133 -359 2167 -325
rect 2133 -427 2167 -393
rect 2133 -495 2167 -461
rect 2133 -563 2167 -529
rect 2133 -631 2167 -597
rect 2133 -699 2167 -665
rect 2133 -767 2167 -733
rect 8033 933 8067 967
rect 8033 865 8067 899
rect 8033 797 8067 831
rect 8033 729 8067 763
rect 8033 661 8067 695
rect 8033 593 8067 627
rect 8033 525 8067 559
rect 8033 457 8067 491
rect 8033 389 8067 423
rect 8033 321 8067 355
rect 8033 253 8067 287
rect 8033 185 8067 219
rect 8033 117 8067 151
rect 8033 49 8067 83
rect 8033 -19 8067 15
rect 8033 -87 8067 -53
rect 8033 -155 8067 -121
rect 8033 -223 8067 -189
rect 8033 -291 8067 -257
rect 8033 -359 8067 -325
rect 8033 -427 8067 -393
rect 8033 -495 8067 -461
rect 8033 -563 8067 -529
rect 8033 -631 8067 -597
rect 8033 -699 8067 -665
rect 8033 -767 8067 -733
rect 2227 -867 2261 -833
rect 2295 -867 2329 -833
rect 2363 -867 2397 -833
rect 2431 -867 2465 -833
rect 2499 -867 2533 -833
rect 2567 -867 2601 -833
rect 2635 -867 2669 -833
rect 2703 -867 2737 -833
rect 2771 -867 2805 -833
rect 2839 -867 2873 -833
rect 2907 -867 2941 -833
rect 2975 -867 3009 -833
rect 3043 -867 3077 -833
rect 3111 -867 3145 -833
rect 3179 -867 3213 -833
rect 3247 -867 3281 -833
rect 3315 -867 3349 -833
rect 3383 -867 3417 -833
rect 3451 -867 3485 -833
rect 3519 -867 3553 -833
rect 3587 -867 3621 -833
rect 3655 -867 3689 -833
rect 3723 -867 3757 -833
rect 3791 -867 3825 -833
rect 3859 -867 3893 -833
rect 3927 -867 3961 -833
rect 3995 -867 4029 -833
rect 4063 -867 4097 -833
rect 4131 -867 4165 -833
rect 4199 -867 4233 -833
rect 4267 -867 4301 -833
rect 4335 -867 4369 -833
rect 4403 -867 4437 -833
rect 4471 -867 4505 -833
rect 4539 -867 4573 -833
rect 4607 -867 4641 -833
rect 4675 -867 4709 -833
rect 4743 -867 4777 -833
rect 4811 -867 4845 -833
rect 4879 -867 4913 -833
rect 4947 -867 4981 -833
rect 5015 -867 5049 -833
rect 5083 -867 5117 -833
rect 5151 -867 5185 -833
rect 5219 -867 5253 -833
rect 5287 -867 5321 -833
rect 5355 -867 5389 -833
rect 5423 -867 5457 -833
rect 5491 -867 5525 -833
rect 5559 -867 5593 -833
rect 5627 -867 5661 -833
rect 5695 -867 5729 -833
rect 5763 -867 5797 -833
rect 5831 -867 5865 -833
rect 5899 -867 5933 -833
rect 5967 -867 6001 -833
rect 6035 -867 6069 -833
rect 6103 -867 6137 -833
rect 6171 -867 6205 -833
rect 6239 -867 6273 -833
rect 6307 -867 6341 -833
rect 6375 -867 6409 -833
rect 6443 -867 6477 -833
rect 6511 -867 6545 -833
rect 6579 -867 6613 -833
rect 6647 -867 6681 -833
rect 6715 -867 6749 -833
rect 6783 -867 6817 -833
rect 6851 -867 6885 -833
rect 6919 -867 6953 -833
rect 6987 -867 7021 -833
rect 7055 -867 7089 -833
rect 7123 -867 7157 -833
rect 7191 -867 7225 -833
rect 7259 -867 7293 -833
rect 7327 -867 7361 -833
rect 7395 -867 7429 -833
rect 7463 -867 7497 -833
rect 7531 -867 7565 -833
rect 7599 -867 7633 -833
rect 7667 -867 7701 -833
rect 7735 -867 7769 -833
rect 7803 -867 7837 -833
rect 7871 -867 7905 -833
rect 7939 -867 7973 -833
<< locali >>
rect 2100 1067 8100 1100
rect 2100 1033 2227 1067
rect 2261 1033 2295 1067
rect 2329 1033 2363 1067
rect 2397 1033 2431 1067
rect 2465 1033 2499 1067
rect 2533 1033 2567 1067
rect 2601 1033 2635 1067
rect 2669 1033 2703 1067
rect 2737 1033 2771 1067
rect 2805 1033 2839 1067
rect 2873 1033 2907 1067
rect 2941 1033 2975 1067
rect 3009 1033 3043 1067
rect 3077 1033 3111 1067
rect 3145 1033 3179 1067
rect 3213 1033 3247 1067
rect 3281 1033 3315 1067
rect 3349 1033 3383 1067
rect 3417 1033 3451 1067
rect 3485 1033 3519 1067
rect 3553 1033 3587 1067
rect 3621 1033 3655 1067
rect 3689 1033 3723 1067
rect 3757 1033 3791 1067
rect 3825 1033 3859 1067
rect 3893 1033 3927 1067
rect 3961 1033 3995 1067
rect 4029 1033 4063 1067
rect 4097 1033 4131 1067
rect 4165 1033 4199 1067
rect 4233 1033 4267 1067
rect 4301 1033 4335 1067
rect 4369 1033 4403 1067
rect 4437 1033 4471 1067
rect 4505 1033 4539 1067
rect 4573 1033 4607 1067
rect 4641 1033 4675 1067
rect 4709 1033 4743 1067
rect 4777 1033 4811 1067
rect 4845 1033 4879 1067
rect 4913 1033 4947 1067
rect 4981 1033 5015 1067
rect 5049 1033 5083 1067
rect 5117 1033 5151 1067
rect 5185 1033 5219 1067
rect 5253 1033 5287 1067
rect 5321 1033 5355 1067
rect 5389 1033 5423 1067
rect 5457 1033 5491 1067
rect 5525 1033 5559 1067
rect 5593 1033 5627 1067
rect 5661 1033 5695 1067
rect 5729 1033 5763 1067
rect 5797 1033 5831 1067
rect 5865 1033 5899 1067
rect 5933 1033 5967 1067
rect 6001 1033 6035 1067
rect 6069 1033 6103 1067
rect 6137 1033 6171 1067
rect 6205 1033 6239 1067
rect 6273 1033 6307 1067
rect 6341 1033 6375 1067
rect 6409 1033 6443 1067
rect 6477 1033 6511 1067
rect 6545 1033 6579 1067
rect 6613 1033 6647 1067
rect 6681 1033 6715 1067
rect 6749 1033 6783 1067
rect 6817 1033 6851 1067
rect 6885 1033 6919 1067
rect 6953 1033 6987 1067
rect 7021 1033 7055 1067
rect 7089 1033 7123 1067
rect 7157 1033 7191 1067
rect 7225 1033 7259 1067
rect 7293 1033 7327 1067
rect 7361 1033 7395 1067
rect 7429 1033 7463 1067
rect 7497 1033 7531 1067
rect 7565 1033 7599 1067
rect 7633 1033 7667 1067
rect 7701 1033 7735 1067
rect 7769 1033 7803 1067
rect 7837 1033 7871 1067
rect 7905 1033 7939 1067
rect 7973 1033 8100 1067
rect 2100 1000 8100 1033
rect 2100 967 2200 1000
rect 2100 933 2133 967
rect 2167 933 2200 967
rect 2100 899 2200 933
rect 2100 865 2133 899
rect 2167 865 2200 899
rect 8000 967 8100 1000
rect 8000 933 8033 967
rect 8067 933 8100 967
rect 8000 899 8100 933
rect 2100 831 2200 865
rect 2100 797 2133 831
rect 2167 797 2200 831
rect 2100 763 2200 797
rect 2100 729 2133 763
rect 2167 729 2200 763
rect 2100 695 2200 729
rect 2100 661 2133 695
rect 2167 661 2200 695
rect 2100 627 2200 661
rect 2100 593 2133 627
rect 2167 593 2200 627
rect 2100 559 2200 593
rect 2100 525 2133 559
rect 2167 525 2200 559
rect 2100 491 2200 525
rect 2100 457 2133 491
rect 2167 457 2200 491
rect 2100 423 2200 457
rect 2100 389 2133 423
rect 2167 389 2200 423
rect 2100 355 2200 389
rect 2100 321 2133 355
rect 2167 321 2200 355
rect 2100 287 2200 321
rect 2100 253 2133 287
rect 2167 253 2200 287
rect 2100 219 2200 253
rect 2100 185 2133 219
rect 2167 185 2200 219
rect 2100 151 2200 185
rect 2100 117 2133 151
rect 2167 117 2200 151
rect 2100 83 2200 117
rect 2100 49 2133 83
rect 2167 49 2200 83
rect 2100 15 2200 49
rect 2100 -19 2133 15
rect 2167 -19 2200 15
rect 2100 -53 2200 -19
rect 2100 -87 2133 -53
rect 2167 -87 2200 -53
rect 2100 -121 2200 -87
rect 2100 -155 2133 -121
rect 2167 -155 2200 -121
rect 2100 -189 2200 -155
rect 2100 -223 2133 -189
rect 2167 -223 2200 -189
rect 2100 -257 2200 -223
rect 2100 -291 2133 -257
rect 2167 -291 2200 -257
rect 2100 -325 2200 -291
rect 2100 -359 2133 -325
rect 2167 -359 2200 -325
rect 2100 -393 2200 -359
rect 2100 -427 2133 -393
rect 2167 -427 2200 -393
rect 2100 -461 2200 -427
rect 2100 -495 2133 -461
rect 2167 -495 2200 -461
rect 2100 -529 2200 -495
rect 2100 -563 2133 -529
rect 2167 -563 2200 -529
rect 2100 -597 2200 -563
rect 2100 -631 2133 -597
rect 2167 -631 2200 -597
rect 2100 -665 2200 -631
rect 2100 -699 2133 -665
rect 2167 -699 2200 -665
rect 2100 -733 2200 -699
rect 2340 167 2620 880
rect 2340 133 2453 167
rect 2487 133 2620 167
rect 2340 67 2620 133
rect 2340 33 2453 67
rect 2487 33 2620 67
rect 2340 -33 2620 33
rect 2340 -67 2453 -33
rect 2487 -67 2620 -33
rect 2340 -700 2620 -67
rect 2100 -767 2133 -733
rect 2167 -767 2200 -733
rect 2100 -800 2200 -767
rect 2880 -800 3000 800
rect 3500 -800 3620 800
rect 4120 -800 4240 800
rect 4720 -800 4840 800
rect 5340 -800 5460 800
rect 5960 -800 6080 800
rect 6580 -800 6700 800
rect 7200 -800 7320 800
rect 7580 167 7860 880
rect 7580 133 7693 167
rect 7727 133 7860 167
rect 7580 67 7860 133
rect 7580 33 7693 67
rect 7727 33 7860 67
rect 7580 -33 7860 33
rect 7580 -67 7693 -33
rect 7727 -67 7860 -33
rect 7580 -700 7860 -67
rect 8000 865 8033 899
rect 8067 865 8100 899
rect 8000 831 8100 865
rect 8000 797 8033 831
rect 8067 797 8100 831
rect 8000 763 8100 797
rect 8000 729 8033 763
rect 8067 729 8100 763
rect 8000 695 8100 729
rect 8000 661 8033 695
rect 8067 661 8100 695
rect 8000 627 8100 661
rect 8000 593 8033 627
rect 8067 593 8100 627
rect 8000 559 8100 593
rect 8000 525 8033 559
rect 8067 525 8100 559
rect 8000 491 8100 525
rect 8000 457 8033 491
rect 8067 457 8100 491
rect 8000 423 8100 457
rect 8000 389 8033 423
rect 8067 389 8100 423
rect 8000 355 8100 389
rect 8000 321 8033 355
rect 8067 321 8100 355
rect 8000 287 8100 321
rect 8000 253 8033 287
rect 8067 253 8100 287
rect 8000 219 8100 253
rect 8000 185 8033 219
rect 8067 185 8100 219
rect 8000 151 8100 185
rect 8000 117 8033 151
rect 8067 117 8100 151
rect 8000 83 8100 117
rect 8000 49 8033 83
rect 8067 49 8100 83
rect 8000 15 8100 49
rect 8000 -19 8033 15
rect 8067 -19 8100 15
rect 8000 -53 8100 -19
rect 8000 -87 8033 -53
rect 8067 -87 8100 -53
rect 8000 -121 8100 -87
rect 8000 -155 8033 -121
rect 8067 -155 8100 -121
rect 8000 -189 8100 -155
rect 8000 -223 8033 -189
rect 8067 -223 8100 -189
rect 8000 -257 8100 -223
rect 8000 -291 8033 -257
rect 8067 -291 8100 -257
rect 8000 -325 8100 -291
rect 8000 -359 8033 -325
rect 8067 -359 8100 -325
rect 8000 -393 8100 -359
rect 8000 -427 8033 -393
rect 8067 -427 8100 -393
rect 8000 -461 8100 -427
rect 8000 -495 8033 -461
rect 8067 -495 8100 -461
rect 8000 -529 8100 -495
rect 8000 -563 8033 -529
rect 8067 -563 8100 -529
rect 8000 -597 8100 -563
rect 8000 -631 8033 -597
rect 8067 -631 8100 -597
rect 8000 -665 8100 -631
rect 8000 -699 8033 -665
rect 8067 -699 8100 -665
rect 8000 -733 8100 -699
rect 8000 -767 8033 -733
rect 8067 -767 8100 -733
rect 8000 -800 8100 -767
rect 2100 -833 8100 -800
rect 2100 -867 2133 -833
rect 2167 -867 2227 -833
rect 2261 -867 2295 -833
rect 2329 -867 2363 -833
rect 2397 -867 2431 -833
rect 2465 -867 2499 -833
rect 2533 -867 2567 -833
rect 2601 -867 2635 -833
rect 2669 -867 2703 -833
rect 2737 -867 2771 -833
rect 2805 -867 2839 -833
rect 2873 -867 2907 -833
rect 2941 -867 2975 -833
rect 3009 -867 3043 -833
rect 3077 -867 3111 -833
rect 3145 -867 3179 -833
rect 3213 -867 3247 -833
rect 3281 -867 3315 -833
rect 3349 -867 3383 -833
rect 3417 -867 3451 -833
rect 3485 -867 3519 -833
rect 3553 -867 3587 -833
rect 3621 -867 3655 -833
rect 3689 -867 3723 -833
rect 3757 -867 3791 -833
rect 3825 -867 3859 -833
rect 3893 -867 3927 -833
rect 3961 -867 3995 -833
rect 4029 -867 4063 -833
rect 4097 -867 4131 -833
rect 4165 -867 4199 -833
rect 4233 -867 4267 -833
rect 4301 -867 4335 -833
rect 4369 -867 4403 -833
rect 4437 -867 4471 -833
rect 4505 -867 4539 -833
rect 4573 -867 4607 -833
rect 4641 -867 4675 -833
rect 4709 -867 4743 -833
rect 4777 -867 4811 -833
rect 4845 -867 4879 -833
rect 4913 -867 4947 -833
rect 4981 -867 5015 -833
rect 5049 -867 5083 -833
rect 5117 -867 5151 -833
rect 5185 -867 5219 -833
rect 5253 -867 5287 -833
rect 5321 -867 5355 -833
rect 5389 -867 5423 -833
rect 5457 -867 5491 -833
rect 5525 -867 5559 -833
rect 5593 -867 5627 -833
rect 5661 -867 5695 -833
rect 5729 -867 5763 -833
rect 5797 -867 5831 -833
rect 5865 -867 5899 -833
rect 5933 -867 5967 -833
rect 6001 -867 6035 -833
rect 6069 -867 6103 -833
rect 6137 -867 6171 -833
rect 6205 -867 6239 -833
rect 6273 -867 6307 -833
rect 6341 -867 6375 -833
rect 6409 -867 6443 -833
rect 6477 -867 6511 -833
rect 6545 -867 6579 -833
rect 6613 -867 6647 -833
rect 6681 -867 6715 -833
rect 6749 -867 6783 -833
rect 6817 -867 6851 -833
rect 6885 -867 6919 -833
rect 6953 -867 6987 -833
rect 7021 -867 7055 -833
rect 7089 -867 7123 -833
rect 7157 -867 7191 -833
rect 7225 -867 7259 -833
rect 7293 -867 7327 -833
rect 7361 -867 7395 -833
rect 7429 -867 7463 -833
rect 7497 -867 7531 -833
rect 7565 -867 7599 -833
rect 7633 -867 7667 -833
rect 7701 -867 7735 -833
rect 7769 -867 7803 -833
rect 7837 -867 7871 -833
rect 7905 -867 7939 -833
rect 7973 -867 8100 -833
rect 2100 -900 8100 -867
<< viali >>
rect 2453 133 2487 167
rect 2453 33 2487 67
rect 2453 -67 2487 -33
rect 7693 133 7727 167
rect 7693 33 7727 67
rect 7693 -67 7727 -33
rect 2133 -867 2167 -833
<< metal1 >>
rect 2660 860 7540 940
rect 1800 176 2100 200
rect 1800 124 1824 176
rect 1876 124 1924 176
rect 1976 124 2024 176
rect 2076 124 2100 176
rect 1800 76 2100 124
rect 1800 24 1824 76
rect 1876 24 1924 76
rect 1976 24 2024 76
rect 2076 24 2100 76
rect 1800 -24 2100 24
rect 1800 -76 1824 -24
rect 1876 -76 1924 -24
rect 1976 -76 2024 -24
rect 2076 -76 2100 -24
rect 1800 -100 2100 -76
rect 2420 176 2520 200
rect 2420 124 2444 176
rect 2496 124 2520 176
rect 2420 76 2520 124
rect 2420 24 2444 76
rect 2496 24 2520 76
rect 2420 -24 2520 24
rect 2420 -76 2444 -24
rect 2496 -76 2520 -24
rect 2420 -100 2520 -76
rect 3180 -324 3320 860
rect 3820 176 3920 200
rect 3820 124 3844 176
rect 3896 124 3920 176
rect 3820 76 3920 124
rect 3820 24 3844 76
rect 3896 24 3920 76
rect 3820 -24 3920 24
rect 3820 -76 3844 -24
rect 3896 -76 3920 -24
rect 3820 -100 3920 -76
rect 3180 -376 3224 -324
rect 3276 -376 3320 -324
rect 3180 -424 3320 -376
rect 3180 -476 3224 -424
rect 3276 -476 3320 -424
rect 3180 -524 3320 -476
rect 3180 -576 3224 -524
rect 3276 -576 3320 -524
rect 3180 -700 3320 -576
rect 4420 -324 4560 860
rect 5060 176 5160 200
rect 5060 124 5084 176
rect 5136 124 5160 176
rect 5060 76 5160 124
rect 5060 24 5084 76
rect 5136 24 5160 76
rect 5060 -24 5160 24
rect 5060 -76 5084 -24
rect 5136 -76 5160 -24
rect 5060 -100 5160 -76
rect 4420 -376 4464 -324
rect 4516 -376 4560 -324
rect 4420 -424 4560 -376
rect 4420 -476 4464 -424
rect 4516 -476 4560 -424
rect 4420 -524 4560 -476
rect 4420 -576 4464 -524
rect 4516 -576 4560 -524
rect 4420 -700 4560 -576
rect 5640 -324 5780 860
rect 6280 176 6380 200
rect 6280 124 6304 176
rect 6356 124 6380 176
rect 6280 76 6380 124
rect 6280 24 6304 76
rect 6356 24 6380 76
rect 6280 -24 6380 24
rect 6280 -76 6304 -24
rect 6356 -76 6380 -24
rect 6280 -100 6380 -76
rect 5640 -376 5684 -324
rect 5736 -376 5780 -324
rect 5640 -424 5780 -376
rect 5640 -476 5684 -424
rect 5736 -476 5780 -424
rect 5640 -524 5780 -476
rect 5640 -576 5684 -524
rect 5736 -576 5780 -524
rect 5640 -700 5780 -576
rect 6860 -324 7000 860
rect 7660 176 7760 200
rect 7660 124 7684 176
rect 7736 124 7760 176
rect 7660 76 7760 124
rect 7660 24 7684 76
rect 7736 24 7760 76
rect 7660 -24 7760 24
rect 7660 -76 7684 -24
rect 7736 -76 7760 -24
rect 7660 -100 7760 -76
rect 8100 176 8400 200
rect 8100 124 8124 176
rect 8176 124 8224 176
rect 8276 124 8324 176
rect 8376 124 8400 176
rect 8100 76 8400 124
rect 8100 24 8124 76
rect 8176 24 8224 76
rect 8276 24 8324 76
rect 8376 24 8400 76
rect 8100 -24 8400 24
rect 8100 -76 8124 -24
rect 8176 -76 8224 -24
rect 8276 -76 8324 -24
rect 8376 -76 8400 -24
rect 8100 -100 8400 -76
rect 6860 -376 6904 -324
rect 6956 -376 7000 -324
rect 6860 -424 7000 -376
rect 6860 -476 6904 -424
rect 6956 -476 7000 -424
rect 6860 -524 7000 -476
rect 6860 -576 6904 -524
rect 6956 -576 7000 -524
rect 6860 -700 7000 -576
rect 2100 -833 2200 -800
rect 2100 -867 2133 -833
rect 2167 -867 2200 -833
rect 2100 -900 2200 -867
rect 5000 -1624 5200 -1600
rect 5000 -1676 5024 -1624
rect 5076 -1676 5124 -1624
rect 5176 -1676 5200 -1624
rect 5000 -1724 5200 -1676
rect 5000 -1776 5024 -1724
rect 5076 -1776 5124 -1724
rect 5176 -1776 5200 -1724
rect 5000 -1800 5200 -1776
<< via1 >>
rect 1824 124 1876 176
rect 1924 124 1976 176
rect 2024 124 2076 176
rect 1824 24 1876 76
rect 1924 24 1976 76
rect 2024 24 2076 76
rect 1824 -76 1876 -24
rect 1924 -76 1976 -24
rect 2024 -76 2076 -24
rect 2444 167 2496 176
rect 2444 133 2453 167
rect 2453 133 2487 167
rect 2487 133 2496 167
rect 2444 124 2496 133
rect 2444 67 2496 76
rect 2444 33 2453 67
rect 2453 33 2487 67
rect 2487 33 2496 67
rect 2444 24 2496 33
rect 2444 -33 2496 -24
rect 2444 -67 2453 -33
rect 2453 -67 2487 -33
rect 2487 -67 2496 -33
rect 2444 -76 2496 -67
rect 3844 124 3896 176
rect 3844 24 3896 76
rect 3844 -76 3896 -24
rect 3224 -376 3276 -324
rect 3224 -476 3276 -424
rect 3224 -576 3276 -524
rect 5084 124 5136 176
rect 5084 24 5136 76
rect 5084 -76 5136 -24
rect 4464 -376 4516 -324
rect 4464 -476 4516 -424
rect 4464 -576 4516 -524
rect 6304 124 6356 176
rect 6304 24 6356 76
rect 6304 -76 6356 -24
rect 5684 -376 5736 -324
rect 5684 -476 5736 -424
rect 5684 -576 5736 -524
rect 7684 167 7736 176
rect 7684 133 7693 167
rect 7693 133 7727 167
rect 7727 133 7736 167
rect 7684 124 7736 133
rect 7684 67 7736 76
rect 7684 33 7693 67
rect 7693 33 7727 67
rect 7727 33 7736 67
rect 7684 24 7736 33
rect 7684 -33 7736 -24
rect 7684 -67 7693 -33
rect 7693 -67 7727 -33
rect 7727 -67 7736 -33
rect 7684 -76 7736 -67
rect 8124 124 8176 176
rect 8224 124 8276 176
rect 8324 124 8376 176
rect 8124 24 8176 76
rect 8224 24 8276 76
rect 8324 24 8376 76
rect 8124 -76 8176 -24
rect 8224 -76 8276 -24
rect 8324 -76 8376 -24
rect 6904 -376 6956 -324
rect 6904 -476 6956 -424
rect 6904 -576 6956 -524
rect 5024 -1676 5076 -1624
rect 5124 -1676 5176 -1624
rect 5024 -1776 5076 -1724
rect 5124 -1776 5176 -1724
<< metal2 >>
rect 1800 176 8400 200
rect 1800 124 1824 176
rect 1876 124 1924 176
rect 1976 124 2024 176
rect 2076 124 2444 176
rect 2496 124 3844 176
rect 3896 124 5084 176
rect 5136 124 6304 176
rect 6356 124 7684 176
rect 7736 124 8124 176
rect 8176 124 8224 176
rect 8276 124 8324 176
rect 8376 124 8400 176
rect 1800 76 8400 124
rect 1800 24 1824 76
rect 1876 24 1924 76
rect 1976 24 2024 76
rect 2076 24 2444 76
rect 2496 24 3844 76
rect 3896 24 5084 76
rect 5136 24 6304 76
rect 6356 24 7684 76
rect 7736 24 8124 76
rect 8176 24 8224 76
rect 8276 24 8324 76
rect 8376 24 8400 76
rect 1800 -24 8400 24
rect 1800 -76 1824 -24
rect 1876 -76 1924 -24
rect 1976 -76 2024 -24
rect 2076 -76 2444 -24
rect 2496 -76 3844 -24
rect 3896 -76 5084 -24
rect 5136 -76 6304 -24
rect 6356 -76 7684 -24
rect 7736 -76 8124 -24
rect 8176 -76 8224 -24
rect 8276 -76 8324 -24
rect 8376 -76 8400 -24
rect 1800 -100 8400 -76
rect 3100 -324 7100 -300
rect 3100 -376 3224 -324
rect 3276 -376 4464 -324
rect 4516 -376 5684 -324
rect 5736 -376 6904 -324
rect 6956 -376 7100 -324
rect 3100 -424 7100 -376
rect 3100 -476 3224 -424
rect 3276 -476 4464 -424
rect 4516 -476 5684 -424
rect 5736 -476 6904 -424
rect 6956 -476 7100 -424
rect 3100 -524 7100 -476
rect 3100 -576 3224 -524
rect 3276 -576 4464 -524
rect 4516 -576 5684 -524
rect 5736 -576 6904 -524
rect 6956 -576 7100 -524
rect 3100 -600 7100 -576
rect 5000 -1624 5200 -600
rect 5000 -1676 5024 -1624
rect 5076 -1676 5124 -1624
rect 5176 -1676 5200 -1624
rect 5000 -1724 5200 -1676
rect 5000 -1776 5024 -1724
rect 5076 -1776 5124 -1724
rect 5176 -1776 5200 -1724
rect 5000 -1800 5200 -1776
use sky130_fd_pr__nfet_g5v0d10v5_7GKDBD  XM6
timestamp 1770083657
transform 1 0 5101 0 1 107
box -2827 -807 2827 807
<< labels >>
flabel metal1 s 5000 -1800 5200 -1600 0 FreeSans 320 0 0 0 IBIAS
port 1 nsew
flabel metal1 s 1860 -40 2060 160 0 FreeSans 320 0 0 0 S
port 2 nsew
flabel metal1 s 2100 -900 2200 -800 0 FreeSans 320 0 0 0 VSS
port 3 nsew
<< end >>
