* SPICE3 file created from 1st-stage.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_1_RK594X m3_120_n5200# m3_n5492_n5200# c1_160_n5160#
+ c1_n5452_n5160# VSUBS
X0 c1_n5452_n5160# m3_n5492_n5200# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X1 c1_n5452_n5160# m3_n5492_n5200# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X2 c1_160_n5160# m3_120_n5200# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X3 c1_160_n5160# m3_120_n5200# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
C0 m3_n5492_n5200# c1_160_n5160# 2.13703f
C1 m3_n5492_n5200# c1_n5452_n5160# 0.11107p
C2 m3_120_n5200# c1_160_n5160# 0.11107p
C3 m3_n5492_n5200# m3_120_n5200# 2.60505f
C4 c1_160_n5160# VSUBS 2.41009f
C5 c1_n5452_n5160# VSUBS 3.9139f
C6 m3_120_n5200# VSUBS 24.0617f
C7 m3_n5492_n5200# VSUBS 22.4584f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7 a_n29_n444# a_n187_n444# a_29_n532# a_n129_n532#
+ a_129_n444# VSUBS
X0 a_129_n444# a_29_n532# a_n29_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.3775 pd=10.08 as=0.68875 ps=5.04 w=4.75 l=0.5
X1 a_n29_n444# a_n129_n532# a_n187_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=1.3775 ps=10.08 w=4.75 l=0.5
C0 a_n29_n444# a_129_n444# 0.42382f
C1 a_n187_n444# a_n29_n444# 0.42382f
C2 a_n129_n532# a_n29_n444# 0.06273f
C3 a_29_n532# a_129_n444# 0.06273f
C4 a_n129_n532# a_n187_n444# 0.06273f
C5 a_29_n532# a_n29_n444# 0.06273f
C6 a_n129_n532# a_29_n532# 0.05942f
C7 a_129_n444# VSUBS 0.45597f
C8 a_n29_n444# VSUBS 0.10803f
C9 a_n187_n444# VSUBS 0.45597f
C10 a_29_n532# VSUBS 0.25901f
C11 a_n129_n532# VSUBS 0.25901f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_838SN6 a_n187_n506# a_129_n506# a_29_n532# a_n129_n532#
+ a_n29_n506# VSUBS
X0 a_129_n506# a_29_n532# a_n29_n506# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.3775 pd=10.08 as=0.68875 ps=5.04 w=4.75 l=0.5
X1 a_n29_n506# a_n129_n532# a_n187_n506# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=1.3775 ps=10.08 w=4.75 l=0.5
C0 a_n29_n506# a_129_n506# 0.42382f
C1 a_n187_n506# a_n29_n506# 0.42382f
C2 a_n129_n532# a_n29_n506# 0.06273f
C3 a_29_n532# a_129_n506# 0.06273f
C4 a_n129_n532# a_n187_n506# 0.06273f
C5 a_29_n532# a_n29_n506# 0.06273f
C6 a_n129_n532# a_29_n532# 0.05942f
C7 a_129_n506# VSUBS 0.45597f
C8 a_n29_n506# VSUBS 0.10803f
C9 a_n187_n506# VSUBS 0.45597f
C10 a_29_n532# VSUBS 0.25901f
C11 a_n129_n532# VSUBS 0.25901f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DQUD5W a_n953_n781# a_2185_n807# a_n587_n807#
+ a_645_n807# a_29_n807# a_2435_n781# a_n2185_n781# a_1261_n807# a_1569_n807# a_279_n781#
+ a_895_n781# a_n2435_n807# a_n1261_n781# a_1511_n781# a_1819_n781# a_n1569_n781#
+ a_n29_n781# a_n645_n781# a_n1511_n807# a_n279_n807# a_n1819_n807# a_n895_n807# a_337_n807#
+ a_953_n807# a_2127_n781# a_n2493_n781# a_587_n781# a_1877_n807# a_n2127_n807# a_1203_n781#
+ a_n1877_n781# a_n337_n781# a_n1203_n807# VSUBS
X0 a_1511_n781# a_1261_n807# a_1203_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X1 a_n1261_n781# a_n1511_n807# a_n1569_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X2 a_n1877_n781# a_n2127_n807# a_n2185_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X3 a_895_n781# a_645_n807# a_587_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X4 a_n1569_n781# a_n1819_n807# a_n1877_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X5 a_n645_n781# a_n895_n807# a_n953_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X6 a_1819_n781# a_1569_n807# a_1511_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X7 a_n29_n781# a_n279_n807# a_n337_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X8 a_n953_n781# a_n1203_n807# a_n1261_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X9 a_2435_n781# a_2185_n807# a_2127_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=1.25
X10 a_n2185_n781# a_n2435_n807# a_n2493_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=1.25
X11 a_1203_n781# a_953_n807# a_895_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X12 a_587_n781# a_337_n807# a_279_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X13 a_2127_n781# a_1877_n807# a_1819_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X14 a_n337_n781# a_n587_n807# a_n645_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X15 a_279_n781# a_29_n807# a_n29_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
C0 a_n587_n807# a_n279_n807# 0.05942f
C1 a_n1819_n807# a_n1569_n781# 0.19032f
C2 a_n1511_n807# a_n1261_n781# 0.19032f
C3 a_n337_n781# a_n279_n807# 0.19032f
C4 a_1511_n781# a_1261_n807# 0.19032f
C5 a_895_n781# a_645_n807# 0.19032f
C6 a_n895_n807# a_n645_n781# 0.19032f
C7 a_n1877_n781# a_n2185_n781# 0.34377f
C8 a_1877_n807# a_2185_n807# 0.05942f
C9 a_337_n807# a_645_n807# 0.05942f
C10 a_n1511_n807# a_n1203_n807# 0.05942f
C11 a_1569_n807# a_1511_n781# 0.19032f
C12 a_587_n781# a_645_n807# 0.19032f
C13 a_1877_n807# a_1819_n781# 0.19032f
C14 a_2127_n781# a_2435_n781# 0.34377f
C15 a_n1877_n781# a_n2127_n807# 0.19032f
C16 a_n953_n781# a_n1261_n781# 0.34377f
C17 a_n1819_n807# a_n1511_n807# 0.05942f
C18 a_1203_n781# a_1511_n781# 0.34377f
C19 a_n953_n781# a_n1203_n807# 0.19032f
C20 a_895_n781# a_953_n807# 0.19032f
C21 a_n587_n807# a_n645_n781# 0.19032f
C22 a_2185_n807# a_2435_n781# 0.19032f
C23 a_n337_n781# a_n29_n781# 0.34377f
C24 a_29_n807# a_n279_n807# 0.05942f
C25 a_1203_n781# a_895_n781# 0.34377f
C26 a_1877_n807# a_1569_n807# 0.05942f
C27 a_1569_n807# a_1819_n781# 0.19032f
C28 a_n337_n781# a_n645_n781# 0.34377f
C29 a_n29_n781# a_n279_n807# 0.19032f
C30 a_n1877_n781# a_n1569_n781# 0.34377f
C31 a_n587_n807# a_n895_n807# 0.05942f
C32 a_29_n807# a_279_n781# 0.19032f
C33 a_1569_n807# a_1261_n807# 0.05942f
C34 a_n29_n781# a_279_n781# 0.34377f
C35 a_645_n807# a_953_n807# 0.05942f
C36 a_337_n807# a_279_n781# 0.19032f
C37 a_n1203_n807# a_n895_n807# 0.05942f
C38 a_279_n781# a_587_n781# 0.34377f
C39 a_n2185_n781# a_n2435_n807# 0.19032f
C40 a_29_n807# a_n29_n781# 0.19032f
C41 a_953_n807# a_1261_n807# 0.05942f
C42 a_n2127_n807# a_n1819_n807# 0.05942f
C43 a_337_n807# a_29_n807# 0.05942f
C44 a_n1261_n781# a_n1569_n781# 0.34377f
C45 a_n953_n781# a_n645_n781# 0.34377f
C46 a_1203_n781# a_1261_n807# 0.19032f
C47 a_587_n781# a_895_n781# 0.34377f
C48 a_337_n807# a_587_n781# 0.19032f
C49 a_2127_n781# a_2185_n807# 0.19032f
C50 a_n2185_n781# a_n2493_n781# 0.34377f
C51 a_n2185_n781# a_n2127_n807# 0.19032f
C52 a_n2435_n807# a_n2493_n781# 0.19032f
C53 a_n2435_n807# a_n2127_n807# 0.05942f
C54 a_n1511_n807# a_n1569_n781# 0.19032f
C55 a_n337_n781# a_n587_n807# 0.19032f
C56 a_1819_n781# a_1511_n781# 0.34377f
C57 a_n1203_n807# a_n1261_n781# 0.19032f
C58 a_n1877_n781# a_n1819_n807# 0.19032f
C59 a_1877_n807# a_2127_n781# 0.19032f
C60 a_1203_n781# a_953_n807# 0.19032f
C61 a_1819_n781# a_2127_n781# 0.34377f
C62 a_n953_n781# a_n895_n807# 0.19032f
C63 a_2435_n781# VSUBS 0.75893f
C64 a_2127_n781# VSUBS 0.26915f
C65 a_1819_n781# VSUBS 0.26915f
C66 a_1511_n781# VSUBS 0.26915f
C67 a_1203_n781# VSUBS 0.26915f
C68 a_895_n781# VSUBS 0.26915f
C69 a_587_n781# VSUBS 0.26915f
C70 a_279_n781# VSUBS 0.26915f
C71 a_n29_n781# VSUBS 0.26915f
C72 a_n337_n781# VSUBS 0.26915f
C73 a_n645_n781# VSUBS 0.26915f
C74 a_n953_n781# VSUBS 0.26915f
C75 a_n1261_n781# VSUBS 0.26915f
C76 a_n1569_n781# VSUBS 0.26915f
C77 a_n1877_n781# VSUBS 0.26915f
C78 a_n2185_n781# VSUBS 0.26915f
C79 a_n2493_n781# VSUBS 0.75893f
C80 a_2185_n807# VSUBS 0.56406f
C81 a_1877_n807# VSUBS 0.52924f
C82 a_1569_n807# VSUBS 0.52924f
C83 a_1261_n807# VSUBS 0.52924f
C84 a_953_n807# VSUBS 0.52924f
C85 a_645_n807# VSUBS 0.52924f
C86 a_337_n807# VSUBS 0.52924f
C87 a_29_n807# VSUBS 0.52924f
C88 a_n279_n807# VSUBS 0.52924f
C89 a_n587_n807# VSUBS 0.52924f
C90 a_n895_n807# VSUBS 0.52924f
C91 a_n1203_n807# VSUBS 0.52924f
C92 a_n1511_n807# VSUBS 0.52924f
C93 a_n1819_n807# VSUBS 0.52924f
C94 a_n2127_n807# VSUBS 0.52924f
C95 a_n2435_n807# VSUBS 0.56406f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DNNC3W a_29_n807# a_n129_n807# a_n29_n781# a_n187_n781#
+ a_129_n781# VSUBS
X0 a_n29_n781# a_n129_n807# a_n187_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=0.5
X1 a_129_n781# a_29_n807# a_n29_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=0.5
C0 a_129_n781# a_29_n807# 0.0968f
C1 a_n29_n781# a_129_n781# 0.66815f
C2 a_n129_n807# a_29_n807# 0.05942f
C3 a_n129_n807# a_n29_n781# 0.0968f
C4 a_n129_n807# a_n187_n781# 0.0968f
C5 a_n29_n781# a_29_n807# 0.0968f
C6 a_n187_n781# a_n29_n781# 0.66815f
C7 a_129_n781# VSUBS 0.7007f
C8 a_n29_n781# VSUBS 0.1527f
C9 a_n187_n781# VSUBS 0.7007f
C10 a_29_n807# VSUBS 0.25717f
C11 a_n129_n807# VSUBS 0.25717f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_DETAA8 a_587_n964# a_1203_n964# a_337_n1061#
+ a_n279_n1061# a_953_n1061# a_n895_n1061# a_n1203_n1061# a_n337_n964# a_n953_n964#
+ a_29_n1061# w_n1297_n1064# a_279_n964# a_895_n964# a_n1261_n964# a_645_n1061# a_n587_n1061#
+ a_n645_n964# a_n29_n964# VSUBS
X0 a_895_n964# a_645_n1061# a_587_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X1 a_n645_n964# a_n895_n1061# a_n953_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X2 a_n29_n964# a_n279_n1061# a_n337_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X3 a_n953_n964# a_n1203_n1061# a_n1261_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1.25
X4 a_1203_n964# a_953_n1061# a_895_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1.25
X5 a_587_n964# a_337_n1061# a_279_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X6 a_n337_n964# a_n587_n1061# a_n645_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X7 a_279_n964# a_29_n1061# a_n29_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
C0 w_n1297_n1064# a_953_n1061# 0.13293f
C1 a_n645_n964# w_n1297_n1064# 0.00517f
C2 a_n895_n1061# a_n953_n964# 0.25181f
C3 a_279_n964# a_587_n964# 0.45807f
C4 a_n29_n964# a_n279_n1061# 0.25181f
C5 a_587_n964# a_645_n1061# 0.25181f
C6 a_279_n964# a_337_n1061# 0.25181f
C7 a_279_n964# a_29_n1061# 0.25181f
C8 a_337_n1061# a_645_n1061# 0.0619f
C9 a_n587_n1061# a_n279_n1061# 0.0619f
C10 a_n337_n964# a_n279_n1061# 0.25181f
C11 w_n1297_n1064# a_n29_n964# 0.00517f
C12 a_587_n964# a_895_n964# 0.45807f
C13 w_n1297_n1064# a_n1203_n1061# 0.13293f
C14 a_29_n1061# a_n279_n1061# 0.0619f
C15 w_n1297_n1064# a_n1261_n964# 0.02956f
C16 w_n1297_n1064# a_587_n964# 0.00517f
C17 a_n645_n964# a_n587_n1061# 0.25181f
C18 a_n645_n964# a_n337_n964# 0.45807f
C19 w_n1297_n1064# a_n587_n1061# 0.12683f
C20 w_n1297_n1064# a_n337_n964# 0.00517f
C21 a_n645_n964# a_n953_n964# 0.45807f
C22 w_n1297_n1064# a_337_n1061# 0.12683f
C23 w_n1297_n1064# a_n953_n964# 0.00517f
C24 w_n1297_n1064# a_29_n1061# 0.12683f
C25 a_n645_n964# a_n895_n1061# 0.25181f
C26 a_n337_n964# a_n29_n964# 0.45807f
C27 a_n1261_n964# a_n1203_n1061# 0.25181f
C28 w_n1297_n1064# a_n895_n1061# 0.12683f
C29 a_n29_n964# a_29_n1061# 0.25181f
C30 a_895_n964# a_645_n1061# 0.25181f
C31 a_n1203_n1061# a_n953_n964# 0.25181f
C32 a_953_n1061# a_645_n1061# 0.0619f
C33 a_n337_n964# a_n587_n1061# 0.25181f
C34 a_1203_n964# a_895_n964# 0.45807f
C35 a_587_n964# a_337_n1061# 0.25181f
C36 a_n1261_n964# a_n953_n964# 0.45807f
C37 a_279_n964# w_n1297_n1064# 0.00517f
C38 a_1203_n964# a_953_n1061# 0.25181f
C39 w_n1297_n1064# a_645_n1061# 0.12683f
C40 a_1203_n964# w_n1297_n1064# 0.02956f
C41 a_337_n1061# a_29_n1061# 0.0619f
C42 a_895_n964# a_953_n1061# 0.25181f
C43 w_n1297_n1064# a_n279_n1061# 0.12683f
C44 a_n895_n1061# a_n1203_n1061# 0.0619f
C45 w_n1297_n1064# a_895_n964# 0.00517f
C46 a_n895_n1061# a_n587_n1061# 0.0619f
C47 a_279_n964# a_n29_n964# 0.45807f
C48 a_1203_n964# VSUBS 0.97158f
C49 a_895_n964# VSUBS 0.34405f
C50 a_587_n964# VSUBS 0.34405f
C51 a_279_n964# VSUBS 0.34405f
C52 a_n29_n964# VSUBS 0.34405f
C53 a_n337_n964# VSUBS 0.34405f
C54 a_n645_n964# VSUBS 0.34405f
C55 a_n953_n964# VSUBS 0.34405f
C56 a_n1261_n964# VSUBS 0.97158f
C57 a_953_n1061# VSUBS 0.44026f
C58 a_645_n1061# VSUBS 0.40993f
C59 a_337_n1061# VSUBS 0.40993f
C60 a_29_n1061# VSUBS 0.40993f
C61 a_n279_n1061# VSUBS 0.40993f
C62 a_n587_n1061# VSUBS 0.40993f
C63 a_n895_n1061# VSUBS 0.40993f
C64 a_n1203_n1061# VSUBS 0.44026f
C65 w_n1297_n1064# VSUBS 16.8247f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_686LYQ a_n587_n807# a_587_n719# a_29_n807# a_n337_n719#
+ a_n279_n807# a_337_n807# a_279_n719# a_n29_n719# a_n645_n719# VSUBS
X0 a_n29_n719# a_n279_n807# a_n337_n719# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X1 a_587_n719# a_337_n807# a_279_n719# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=1.25
X2 a_n337_n719# a_n587_n807# a_n645_n719# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=1.25
X3 a_279_n719# a_29_n807# a_n29_n719# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
C0 a_279_n719# a_n29_n719# 0.34377f
C1 a_29_n807# a_337_n807# 0.05942f
C2 a_n279_n807# a_n337_n719# 0.19032f
C3 a_n337_n719# a_n587_n807# 0.19032f
C4 a_n337_n719# a_n29_n719# 0.34377f
C5 a_279_n719# a_587_n719# 0.34377f
C6 a_29_n807# a_n279_n807# 0.05942f
C7 a_n645_n719# a_n587_n807# 0.19032f
C8 a_279_n719# a_337_n807# 0.19032f
C9 a_29_n807# a_n29_n719# 0.19032f
C10 a_29_n807# a_279_n719# 0.19032f
C11 a_n279_n807# a_n587_n807# 0.05942f
C12 a_n279_n807# a_n29_n719# 0.19032f
C13 a_n337_n719# a_n645_n719# 0.34377f
C14 a_587_n719# a_337_n807# 0.19032f
C15 a_587_n719# VSUBS 0.75893f
C16 a_279_n719# VSUBS 0.26915f
C17 a_n29_n719# VSUBS 0.26915f
C18 a_n337_n719# VSUBS 0.26915f
C19 a_n645_n719# VSUBS 0.75893f
C20 a_337_n807# VSUBS 0.56406f
C21 a_29_n807# VSUBS 0.52924f
C22 a_n279_n807# VSUBS 0.52924f
C23 a_n587_n807# VSUBS 0.56406f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y a_29_n1001# w_n223_n1004# a_n129_n1001#
+ a_n29_n904# a_n187_n904# a_129_n904# VSUBS
X0 a_129_n904# a_29_n1001# a_n29_n904# w_n223_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=2.726 pd=19.38 as=1.363 ps=9.69 w=9.4 l=0.5
X1 a_n29_n904# a_n129_n1001# a_n187_n904# w_n223_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=2.726 ps=19.38 w=9.4 l=0.5
C0 a_29_n1001# w_n223_n1004# 0.07336f
C1 a_n29_n904# a_129_n904# 0.83696f
C2 a_n187_n904# a_n29_n904# 0.83696f
C3 a_n129_n1001# a_n187_n904# 0.12034f
C4 a_n129_n1001# a_n29_n904# 0.12034f
C5 w_n223_n1004# a_129_n904# 0.02814f
C6 w_n223_n1004# a_n187_n904# 0.02814f
C7 w_n223_n1004# a_n29_n904# 0.0052f
C8 w_n223_n1004# a_n129_n1001# 0.07336f
C9 a_29_n1001# a_129_n904# 0.12034f
C10 a_29_n1001# a_n29_n904# 0.12034f
C11 a_29_n1001# a_n129_n1001# 0.0619f
C12 a_129_n904# VSUBS 0.84164f
C13 a_n29_n904# VSUBS 0.17835f
C14 a_n187_n904# VSUBS 0.84164f
C15 a_29_n1001# VSUBS 0.18948f
C16 a_n129_n1001# VSUBS 0.18948f
C17 w_n223_n1004# VSUBS 2.7322f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Y7F49Y a_n337_n904# a_n1203_n1001# a_n953_n904#
+ a_2185_n1001# a_29_n1001# w_n2529_n1004# a_n2185_n904# a_2435_n904# a_n2435_n1001#
+ a_279_n904# a_1877_n1001# a_895_n904# a_1261_n1001# a_1511_n904# a_n1261_n904# a_n1569_n904#
+ a_1819_n904# a_645_n1001# a_n587_n1001# a_n1511_n1001# a_n29_n904# a_n645_n904#
+ a_2127_n904# a_n2493_n904# a_n2127_n1001# a_1569_n1001# a_587_n904# a_1203_n904#
+ a_n1877_n904# a_953_n1001# a_337_n1001# a_n279_n1001# a_n895_n1001# a_n1819_n1001#
+ VSUBS
X0 a_n1877_n904# a_n2127_n1001# a_n2185_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X1 a_895_n904# a_645_n1001# a_587_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X2 a_n1569_n904# a_n1819_n1001# a_n1877_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X3 a_n645_n904# a_n895_n1001# a_n953_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X4 a_1819_n904# a_1569_n1001# a_1511_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X5 a_n29_n904# a_n279_n1001# a_n337_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X6 a_n2185_n904# a_n2435_n1001# a_n2493_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=2.726 ps=19.38 w=9.4 l=1.25
X7 a_n953_n904# a_n1203_n1001# a_n1261_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X8 a_1203_n904# a_953_n1001# a_895_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X9 a_2435_n904# a_2185_n1001# a_2127_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=2.726 pd=19.38 as=1.363 ps=9.69 w=9.4 l=1.25
X10 a_587_n904# a_337_n1001# a_279_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X11 a_2127_n904# a_1877_n1001# a_1819_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X12 a_n337_n904# a_n587_n1001# a_n645_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X13 a_279_n904# a_29_n1001# a_n29_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X14 a_n1261_n904# a_n1511_n1001# a_n1569_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X15 a_1511_n904# a_1261_n1001# a_1203_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
C0 w_n2529_n1004# a_895_n904# 0.00341f
C1 a_n953_n904# w_n2529_n1004# 0.00341f
C2 a_587_n904# a_895_n904# 0.34564f
C3 a_279_n904# w_n2529_n1004# 0.00341f
C4 a_1569_n1001# w_n2529_n1004# 0.12683f
C5 a_279_n904# a_587_n904# 0.34564f
C6 a_1877_n1001# a_2185_n1001# 0.0619f
C7 a_279_n904# a_337_n1001# 0.19111f
C8 a_n953_n904# a_n895_n1001# 0.19111f
C9 a_1203_n904# a_895_n904# 0.34564f
C10 a_1261_n1001# a_1511_n904# 0.19111f
C11 a_279_n904# a_29_n1001# 0.19111f
C12 a_1569_n1001# a_1819_n904# 0.19111f
C13 a_1569_n1001# a_1877_n1001# 0.0619f
C14 w_n2529_n1004# a_2435_n904# 0.02194f
C15 w_n2529_n1004# a_1511_n904# 0.00341f
C16 a_n2127_n1001# a_n1877_n904# 0.19111f
C17 a_n2127_n1001# w_n2529_n1004# 0.12683f
C18 a_2127_n904# a_2435_n904# 0.34564f
C19 a_n1569_n904# a_n1819_n1001# 0.19111f
C20 w_n2529_n1004# a_645_n1001# 0.12683f
C21 a_587_n904# a_645_n1001# 0.19111f
C22 a_1511_n904# a_1203_n904# 0.34564f
C23 a_n29_n904# w_n2529_n1004# 0.00341f
C24 a_337_n1001# a_645_n1001# 0.0619f
C25 a_1819_n904# a_1511_n904# 0.34564f
C26 a_n2435_n1001# a_n2185_n904# 0.19111f
C27 a_n587_n1001# a_n279_n1001# 0.0619f
C28 a_n1569_n904# a_n1511_n1001# 0.19111f
C29 a_2435_n904# a_2185_n1001# 0.19111f
C30 w_n2529_n1004# a_n279_n1001# 0.12683f
C31 a_n645_n904# a_n337_n904# 0.34564f
C32 a_n29_n904# a_29_n1001# 0.19111f
C33 a_1261_n1001# a_953_n1001# 0.0619f
C34 a_n587_n1001# a_n337_n904# 0.19111f
C35 a_n1511_n1001# a_n1203_n1001# 0.0619f
C36 a_n1569_n904# a_n1261_n904# 0.34564f
C37 w_n2529_n1004# a_n337_n904# 0.00341f
C38 a_29_n1001# a_n279_n1001# 0.0619f
C39 a_n1819_n1001# a_n1511_n1001# 0.0619f
C40 a_n2493_n904# a_n2185_n904# 0.34564f
C41 w_n2529_n1004# a_953_n1001# 0.12683f
C42 a_1569_n1001# a_1511_n904# 0.19111f
C43 a_895_n904# a_645_n1001# 0.19111f
C44 a_n2185_n904# a_n1877_n904# 0.34564f
C45 w_n2529_n1004# a_n2185_n904# 0.00341f
C46 a_n1203_n1001# a_n1261_n904# 0.19111f
C47 a_1203_n904# a_953_n1001# 0.19111f
C48 a_n1569_n904# a_n1877_n904# 0.34564f
C49 a_n1569_n904# w_n2529_n1004# 0.00341f
C50 a_n29_n904# a_279_n904# 0.34564f
C51 w_n2529_n1004# a_n1203_n1001# 0.12683f
C52 a_n1819_n1001# a_n1877_n904# 0.19111f
C53 w_n2529_n1004# a_n1819_n1001# 0.12683f
C54 a_n1511_n1001# a_n1261_n904# 0.19111f
C55 a_n1203_n1001# a_n895_n1001# 0.0619f
C56 a_953_n1001# a_895_n904# 0.19111f
C57 a_n2435_n1001# a_n2493_n904# 0.19111f
C58 w_n2529_n1004# a_n1511_n1001# 0.12683f
C59 w_n2529_n1004# a_n2435_n1001# 0.13293f
C60 w_n2529_n1004# a_n1261_n904# 0.00341f
C61 a_n29_n904# a_n279_n1001# 0.19111f
C62 a_n645_n904# a_n587_n1001# 0.19111f
C63 a_n953_n904# a_n1203_n1001# 0.19111f
C64 w_n2529_n1004# a_1261_n1001# 0.12683f
C65 a_n645_n904# w_n2529_n1004# 0.00341f
C66 w_n2529_n1004# a_n2493_n904# 0.02194f
C67 a_953_n1001# a_645_n1001# 0.0619f
C68 a_n2127_n1001# a_n2185_n904# 0.19111f
C69 w_n2529_n1004# a_n587_n1001# 0.12683f
C70 a_n29_n904# a_n337_n904# 0.34564f
C71 a_n645_n904# a_n895_n1001# 0.19111f
C72 w_n2529_n1004# a_n1877_n904# 0.00341f
C73 a_1261_n1001# a_1203_n904# 0.19111f
C74 w_n2529_n1004# a_587_n904# 0.00341f
C75 a_n587_n1001# a_n895_n1001# 0.0619f
C76 w_n2529_n1004# a_2127_n904# 0.00341f
C77 a_n279_n1001# a_n337_n904# 0.19111f
C78 w_n2529_n1004# a_337_n1001# 0.12683f
C79 a_337_n1001# a_587_n904# 0.19111f
C80 w_n2529_n1004# a_n895_n1001# 0.12683f
C81 w_n2529_n1004# a_1203_n904# 0.00341f
C82 w_n2529_n1004# a_29_n1001# 0.12683f
C83 a_n2127_n1001# a_n1819_n1001# 0.0619f
C84 a_1819_n904# w_n2529_n1004# 0.00341f
C85 w_n2529_n1004# a_1877_n1001# 0.12683f
C86 a_337_n1001# a_29_n1001# 0.0619f
C87 a_1819_n904# a_2127_n904# 0.34564f
C88 a_n953_n904# a_n1261_n904# 0.34564f
C89 a_2127_n904# a_1877_n1001# 0.19111f
C90 w_n2529_n1004# a_2185_n1001# 0.13293f
C91 a_2127_n904# a_2185_n1001# 0.19111f
C92 a_n953_n904# a_n645_n904# 0.34564f
C93 a_1569_n1001# a_1261_n1001# 0.0619f
C94 a_1819_n904# a_1877_n1001# 0.19111f
C95 a_n2127_n1001# a_n2435_n1001# 0.0619f
C96 a_2435_n904# VSUBS 0.72996f
C97 a_2127_n904# VSUBS 0.25611f
C98 a_1819_n904# VSUBS 0.25611f
C99 a_1511_n904# VSUBS 0.25611f
C100 a_1203_n904# VSUBS 0.25611f
C101 a_895_n904# VSUBS 0.25611f
C102 a_587_n904# VSUBS 0.25611f
C103 a_279_n904# VSUBS 0.25611f
C104 a_n29_n904# VSUBS 0.25611f
C105 a_n337_n904# VSUBS 0.25611f
C106 a_n645_n904# VSUBS 0.25611f
C107 a_n953_n904# VSUBS 0.25611f
C108 a_n1261_n904# VSUBS 0.25611f
C109 a_n1569_n904# VSUBS 0.25611f
C110 a_n1877_n904# VSUBS 0.25611f
C111 a_n2185_n904# VSUBS 0.25611f
C112 a_n2493_n904# VSUBS 0.72996f
C113 a_2185_n1001# VSUBS 0.44026f
C114 a_1877_n1001# VSUBS 0.40993f
C115 a_1569_n1001# VSUBS 0.40993f
C116 a_1261_n1001# VSUBS 0.40993f
C117 a_953_n1001# VSUBS 0.40993f
C118 a_645_n1001# VSUBS 0.40993f
C119 a_337_n1001# VSUBS 0.40993f
C120 a_29_n1001# VSUBS 0.40993f
C121 a_n279_n1001# VSUBS 0.40993f
C122 a_n587_n1001# VSUBS 0.40993f
C123 a_n895_n1001# VSUBS 0.40993f
C124 a_n1203_n1001# VSUBS 0.40993f
C125 a_n1511_n1001# VSUBS 0.40993f
C126 a_n1819_n1001# VSUBS 0.40993f
C127 a_n2127_n1001# VSUBS 0.40993f
C128 a_n2435_n1001# VSUBS 0.44026f
C129 w_n2529_n1004# VSUBS 30.9853f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AXYYHE w_n303_n564# a_n267_n464# a_29_n561# a_209_n464#
+ a_n29_n464# a_n209_n561# VSUBS
X0 a_n29_n464# a_n209_n561# a_n267_n464# w_n303_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.9
X1 a_209_n464# a_29_n561# a_n29_n464# w_n303_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.9
C0 a_n29_n464# a_209_n464# 0.29682f
C1 a_n267_n464# a_n29_n464# 0.29682f
C2 a_n267_n464# a_n209_n561# 0.10455f
C3 a_n29_n464# w_n303_n564# 0.00519f
C4 a_n209_n561# w_n303_n564# 0.10539f
C5 a_29_n561# a_n29_n464# 0.10455f
C6 a_29_n561# a_n209_n561# 0.0619f
C7 a_n29_n464# a_n209_n561# 0.10455f
C8 a_209_n464# w_n303_n564# 0.01763f
C9 a_29_n561# a_209_n464# 0.10455f
C10 a_n267_n464# w_n303_n564# 0.01763f
C11 a_29_n561# w_n303_n564# 0.10539f
C12 a_209_n464# VSUBS 0.4826f
C13 a_n29_n464# VSUBS 0.15094f
C14 a_n267_n464# VSUBS 0.4826f
C15 a_29_n561# VSUBS 0.32575f
C16 a_n209_n561# VSUBS 0.32575f
C17 w_n303_n564# VSUBS 2.11252f
.ends

.subckt x1st-stage VP VN IBIAS VSS OUT VDD
Xsky130_fd_pr__cap_mim_m3_1_RK594X_0 m1_7460_n3800# m1_7460_n3800# m1_8320_n4220#
+ m1_8320_n4220# VSS sky130_fd_pr__cap_mim_m3_1_RK594X
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_5 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_2 m1_7460_n3800# m1_7460_n3800# VN VN li_9700_n5600#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_6 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_3 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
XXM24 VSS IBIAS IBIAS IBIAS IBIAS IBIAS VSS IBIAS IBIAS VSS VSS IBIAS IBIAS VSS li_9700_n5600#
+ VSS IBIAS li_9700_n5600# IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS VSS IBIAS li_9700_n5600#
+ IBIAS IBIAS IBIAS li_9700_n5600# VSS IBIAS VSS sky130_fd_pr__nfet_g5v0d10v5_DQUD5W
XXM25 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_DNNC3W
Xsky130_fd_pr__cap_mim_m3_1_RK594X_1 m1_7460_n3800# m1_7460_n3800# m1_8320_n4220#
+ m1_8320_n4220# VSS sky130_fd_pr__cap_mim_m3_1_RK594X
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7 li_9700_n5600# m1_7460_n3800# VN VN m1_7460_n3800#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_8 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_4 m1_10280_n4680# m1_10280_n4680# VP VP li_9700_n5600#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
XXM27 OUT OUT m1_7460_n3800# m1_7460_n3800# m1_7460_n3800# m1_7460_n3800# m1_7460_n3800#
+ VDD VDD m1_7460_n3800# VDD VDD VDD OUT m1_7460_n3800# m1_7460_n3800# OUT OUT VSS
+ sky130_fd_pr__pfet_g5v0d10v5_DETAA8
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_9 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_5 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
XXM28 IBIAS OUT IBIAS VSS IBIAS IBIAS VSS OUT OUT VSS sky130_fd_pr__nfet_g5v0d10v5_686LYQ
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_6 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_DNNC3W_0 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_DNNC3W
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_7 m1_10280_n4680# m1_10280_n4680# VP VP li_9700_n5600#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_8 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__pfet_g5v0d10v5_DU7D3Y_0 VDD VDD VDD VDD VDD VDD VSS sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_9 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_686LYQ_0 IBIAS OUT IBIAS VSS IBIAS IBIAS VSS OUT OUT
+ VSS sky130_fd_pr__nfet_g5v0d10v5_686LYQ
XXM2 VDD m1_10280_n4680# VDD m1_10280_n4680# m1_10280_n4680# VDD VDD m1_10280_n4680#
+ m1_10280_n4680# VDD m1_10280_n4680# VDD m1_10280_n4680# VDD m1_10280_n4680# VDD
+ m1_7460_n3800# m1_10280_n4680# m1_10280_n4680# m1_10280_n4680# m1_10280_n4680# m1_7460_n3800#
+ VDD m1_10280_n4680# m1_10280_n4680# m1_10280_n4680# m1_7460_n3800# m1_10280_n4680#
+ m1_7460_n3800# m1_10280_n4680# m1_10280_n4680# m1_10280_n4680# m1_10280_n4680# m1_10280_n4680#
+ VSS sky130_fd_pr__pfet_g5v0d10v5_Y7F49Y
XXM4 VDD VDD VDD VDD VDD VDD VSS sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y
Xsky130_fd_pr__pfet_g5v0d10v5_DETAA8_0 OUT OUT m1_7460_n3800# m1_7460_n3800# m1_7460_n3800#
+ m1_7460_n3800# m1_7460_n3800# VDD VDD m1_7460_n3800# VDD VDD VDD OUT m1_7460_n3800#
+ m1_7460_n3800# OUT OUT VSS sky130_fd_pr__pfet_g5v0d10v5_DETAA8
Xsky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0 VDD m1_8320_n4220# VSS m1_8320_n4220# OUT VSS
+ VSS sky130_fd_pr__pfet_g5v0d10v5_AXYYHE
Xsky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1 VDD m1_8320_n4220# VSS m1_8320_n4220# OUT VSS
+ VSS sky130_fd_pr__pfet_g5v0d10v5_AXYYHE
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10 li_9700_n5600# m1_10280_n4680# VP VP m1_10280_n4680#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_11 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_0 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_1 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2 li_9700_n5600# m1_10280_n4680# VP VP m1_10280_n4680#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_3 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_10 m1_7460_n3800# m1_7460_n3800# VN VN li_9700_n5600#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_0 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4 li_9700_n5600# m1_7460_n3800# VN VN m1_7460_n3800#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_11 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_1 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
C0 VDD m1_10280_n4680# 24.65616f
C1 VN IBIAS 1.04429f
C2 m1_8320_n4220# VP 0.10106f
C3 VDD m1_7460_n3800# 32.61767f
C4 a_17500_n7340# li_9700_n5600# 0.00143f
C5 VDD a_7360_n3320# 1.62535f
C6 VN VP 7.73234f
C7 a_18890_n7340# IBIAS 0.02687f
C8 OUT li_9700_n5600# 0.01117f
C9 OUT a_19390_n3320# 0.11581f
C10 VDD a_16800_n3320# 1.57554f
C11 a_8320_n5020# IBIAS 0
C12 OUT a_18500_n4990# 0.03399f
C13 VDD a_17500_n7340# 0
C14 m1_8320_n4220# m1_10280_n4680# 0
C15 a_8920_n5020# IBIAS 0
C16 m1_7460_n3800# m1_8320_n4220# 6.41884f
C17 VN m1_10280_n4680# 1.03165f
C18 VDD OUT 8.9719f
C19 m1_10280_n4680# a_17900_n4990# 0
C20 a_7360_n3320# m1_8320_n4220# 0.00245f
C21 m1_7460_n3800# VN 2.34721f
C22 m1_7460_n3800# a_17900_n4990# 0.0109f
C23 m1_7460_n3800# a_18890_n7340# 0.00777f
C24 VDD a_7840_n7320# 0.01447f
C25 m1_8320_n4220# a_17500_n7340# 0.00308f
C26 a_9950_n3320# m1_10280_n4680# 0.0049f
C27 m1_7460_n3800# a_8320_n5020# 0.00261f
C28 VN a_17500_n7340# 0.02278f
C29 a_9230_n7320# IBIAS 0.03414f
C30 m1_7460_n3800# a_9950_n3320# 0.04409f
C31 m1_8320_n4220# OUT 6.36335f
C32 a_8920_n5020# m1_10280_n4680# 0
C33 m1_7460_n3800# a_8920_n5020# 0.00993f
C34 VN OUT 1.0288f
C35 a_9230_n7320# VP 0.02057f
C36 a_18890_n7340# a_17500_n7340# 0.01812f
C37 OUT a_17900_n4990# 0.02228f
C38 VDD li_9700_n5600# 0.10708f
C39 VDD a_19390_n3320# 1.61879f
C40 OUT a_18890_n7340# 0.16217f
C41 m1_8320_n4220# a_7840_n7320# 0.00986f
C42 VDD a_18500_n4990# 0.80948f
C43 VN a_7840_n7320# 0
C44 OUT a_8320_n5020# 0.0357f
C45 a_9230_n7320# m1_10280_n4680# 0
C46 a_9950_n3320# OUT 0.117f
C47 IBIAS VP 1.03049f
C48 m1_7460_n3800# a_9230_n7320# 0.00141f
C49 OUT a_8920_n5020# 0.01991f
C50 m1_8320_n4220# li_9700_n5600# 0.00805f
C51 m1_8320_n4220# a_19390_n3320# 0.00245f
C52 VN li_9700_n5600# 7.23164f
C53 a_17900_n4990# li_9700_n5600# 0
C54 m1_8320_n4220# a_18500_n4990# 0.06986f
C55 IBIAS m1_10280_n4680# 0.23417f
C56 a_17900_n4990# a_18500_n4990# 0.02883f
C57 m1_7460_n3800# IBIAS 0.16844f
C58 VDD m1_8320_n4220# 4.41391f
C59 m1_10280_n4680# VP 1.85645f
C60 OUT a_9230_n7320# 0.16185f
C61 VDD VN 0.33524f
C62 m1_7460_n3800# VP 2.03905f
C63 VDD a_17900_n4990# 0.72612f
C64 a_8920_n5020# li_9700_n5600# 0
C65 VDD a_18890_n7340# 0.01405f
C66 a_17500_n7340# IBIAS 0.03437f
C67 a_7840_n7320# a_9230_n7320# 0.01812f
C68 VDD a_8320_n5020# 0.77301f
C69 OUT IBIAS 3.54922f
C70 VDD a_9950_n3320# 1.58528f
C71 m1_7460_n3800# m1_10280_n4680# 13.76171f
C72 VN m1_8320_n4220# 0.10069f
C73 VDD a_8920_n5020# 0.75752f
C74 m1_8320_n4220# a_17900_n4990# 0.06122f
C75 OUT VP 0.93708f
C76 m1_7460_n3800# a_7360_n3320# 0.07501f
C77 a_16800_n3320# m1_10280_n4680# 0.00476f
C78 m1_8320_n4220# a_18890_n7340# 0.00982f
C79 a_9230_n7320# li_9700_n5600# 0.00143f
C80 a_7840_n7320# IBIAS 0.02676f
C81 m1_7460_n3800# a_16800_n3320# 0.04657f
C82 VN a_18890_n7340# 0
C83 a_17500_n7340# m1_10280_n4680# 0.00103f
C84 m1_8320_n4220# a_8320_n5020# 0.07283f
C85 m1_7460_n3800# a_17500_n7340# 0.00137f
C86 OUT m1_10280_n4680# 0.16505f
C87 m1_8320_n4220# a_8920_n5020# 0.06092f
C88 VDD a_9230_n7320# 0.00137f
C89 m1_7460_n3800# OUT 5.89997f
C90 IBIAS li_9700_n5600# 5.45001f
C91 a_7360_n3320# OUT 0.11783f
C92 VP li_9700_n5600# 7.48119f
C93 IBIAS a_18500_n4990# 0
C94 a_16800_n3320# OUT 0.11914f
C95 m1_7460_n3800# a_7840_n7320# 0.01389f
C96 OUT a_17500_n7340# 0.15796f
C97 a_8920_n5020# a_8320_n5020# 0.02883f
C98 VDD IBIAS 0.37869f
C99 m1_8320_n4220# a_9230_n7320# 0.00311f
C100 VDD VP 0.42134f
C101 m1_10280_n4680# li_9700_n5600# 5.46013f
C102 VN a_9230_n7320# 0.00277f
C103 m1_7460_n3800# li_9700_n5600# 4.9898f
C104 m1_7460_n3800# a_19390_n3320# 0.05674f
C105 OUT a_7840_n7320# 0.1653f
C106 m1_7460_n3800# a_18500_n4990# 0.00583f
C107 m1_8320_n4220# IBIAS 0.58635f
C108 a_18890_n7340# VSS 1.46251f 
C109 a_17500_n7340# VSS 1.4904f
C110 a_18500_n4990# VSS 0.04329f 
C111 a_17900_n4990# VSS 0.09855f 
C112 a_9230_n7320# VSS 1.46852f 
C113 a_7840_n7320# VSS 1.48112f 
C114 a_8920_n5020# VSS 0.10741f 
C115 a_8320_n5020# VSS 0.0446f 
C116 a_19390_n3320# VSS 0.08083f 
C117 a_16800_n3320# VSS 0.04815f 
C118 a_9950_n3320# VSS 0.04836f 
C119 a_7360_n3320# VSS 0.08311f 
C120 VP VSS 7.38831f
C121 VDD VSS 0.17127p
C122 OUT VSS 21.76822f
C123 m1_10280_n4680# VSS 14.71998f
C124 m1_8320_n4220# VSS 21.12795f
C125 li_9700_n5600# VSS 28.38409f
C126 IBIAS VSS 43.2622f
C127 m1_7460_n3800# VSS 0.12166p
C128 VN VSS 7.51773f
.ends

