magic
tech sky130A
magscale 1 2
timestamp 1770000594
<< nwell >>
rect 1240 -160 7440 2340
<< nsubdiff >>
rect 1300 2280 7400 2300
rect 1300 2220 1420 2280
rect 7280 2220 7400 2280
rect 1300 2200 7400 2220
rect 1300 2180 1400 2200
rect 1300 20 1320 2180
rect 1380 20 1400 2180
rect 1300 0 1400 20
rect 7300 2180 7400 2200
rect 7300 20 7320 2180
rect 7380 20 7400 2180
rect 7300 0 7400 20
rect 1300 -20 7400 0
rect 1300 -80 1420 -20
rect 7280 -80 7400 -20
rect 1300 -100 7400 -80
<< nsubdiffcont >>
rect 1420 2220 7280 2280
rect 1320 20 1380 2180
rect 7320 20 7380 2180
rect 1420 -80 7280 -20
<< locali >>
rect 1300 2280 7400 2300
rect 1300 2220 1420 2280
rect 7280 2220 7400 2280
rect 1300 2200 7400 2220
rect 1300 2180 1400 2200
rect 1300 20 1320 2180
rect 1380 20 1400 2180
rect 1560 160 1860 2080
rect 2120 200 2240 2200
rect 2740 200 2860 2200
rect 3040 160 3160 2080
rect 3360 200 3480 2200
rect 3960 200 4080 2200
rect 4280 260 4400 2080
rect 4200 160 4500 260
rect 4580 200 4700 2200
rect 5200 200 5320 2200
rect 5500 160 5620 2080
rect 5820 200 5940 2200
rect 6440 200 6560 2200
rect 7300 2180 7400 2200
rect 6800 160 7100 2080
rect 1560 140 7100 160
rect 1560 80 4300 140
rect 4200 60 4300 80
rect 4380 80 7100 140
rect 4380 60 4500 80
rect 4200 40 4500 60
rect 1300 0 1400 20
rect 7300 20 7320 2180
rect 7380 20 7400 2180
rect 7300 0 7400 20
rect 1300 -20 7400 0
rect 1300 -80 1320 -20
rect 1380 -80 1420 -20
rect 7280 -80 7400 -20
rect 1300 -100 7400 -80
rect 4200 -280 4220 -220
rect 4280 -280 4320 -220
rect 4380 -280 4420 -220
rect 4480 -280 4500 -220
rect 4200 -320 4500 -280
rect 4200 -380 4220 -320
rect 4280 -380 4320 -320
rect 4380 -380 4420 -320
rect 4480 -380 4500 -320
rect 4200 -420 4500 -380
rect 4200 -480 4220 -420
rect 4280 -480 4320 -420
rect 4380 -480 4420 -420
rect 4480 -480 4500 -420
rect 4200 -500 4500 -480
<< viali >>
rect 4300 60 4380 140
rect 1320 -80 1380 -20
rect 4220 -280 4280 -220
rect 4320 -280 4380 -220
rect 4420 -280 4480 -220
rect 4220 -380 4280 -320
rect 4320 -380 4380 -320
rect 4420 -380 4480 -320
rect 4220 -480 4280 -420
rect 4320 -480 4380 -420
rect 4420 -480 4480 -420
<< metal1 >>
rect 900 1280 1200 1300
rect 900 1220 920 1280
rect 980 1220 1020 1280
rect 1080 1220 1120 1280
rect 1180 1220 1200 1280
rect 900 1180 1200 1220
rect 900 1120 920 1180
rect 980 1120 1020 1180
rect 1080 1120 1120 1180
rect 1180 1120 1200 1180
rect 900 1080 1200 1120
rect 900 1020 920 1080
rect 980 1020 1020 1080
rect 1080 1020 1120 1080
rect 1180 1020 1200 1080
rect 900 1000 1200 1020
rect 2400 1280 2600 1300
rect 2400 1220 2420 1280
rect 2480 1220 2520 1280
rect 2580 1220 2600 1280
rect 2400 1180 2600 1220
rect 2400 1120 2420 1180
rect 2480 1120 2520 1180
rect 2580 1120 2600 1180
rect 2400 1080 2600 1120
rect 2400 1020 2420 1080
rect 2480 1020 2520 1080
rect 2580 1020 2600 1080
rect 2400 1000 2600 1020
rect 3600 1280 3800 1300
rect 3600 1220 3620 1280
rect 3680 1220 3720 1280
rect 3780 1220 3800 1280
rect 3600 1180 3800 1220
rect 3600 1120 3620 1180
rect 3680 1120 3720 1180
rect 3780 1120 3800 1180
rect 3600 1080 3800 1120
rect 3600 1020 3620 1080
rect 3680 1020 3720 1080
rect 3780 1020 3800 1080
rect 3600 1000 3800 1020
rect 4860 1280 5060 1300
rect 4860 1220 4880 1280
rect 4940 1220 4980 1280
rect 5040 1220 5060 1280
rect 4860 1180 5060 1220
rect 4860 1120 4880 1180
rect 4940 1120 4980 1180
rect 5040 1120 5060 1180
rect 4860 1080 5060 1120
rect 4860 1020 4880 1080
rect 4940 1020 4980 1080
rect 5040 1020 5060 1080
rect 4860 1000 5060 1020
rect 6100 1280 6300 1300
rect 6100 1220 6120 1280
rect 6180 1220 6220 1280
rect 6280 1220 6300 1280
rect 6100 1180 6300 1220
rect 6100 1120 6120 1180
rect 6180 1120 6220 1180
rect 6280 1120 6300 1180
rect 6100 1080 6300 1120
rect 6100 1020 6120 1080
rect 6180 1020 6220 1080
rect 6280 1020 6300 1080
rect 6100 1000 6300 1020
rect 7500 1280 7800 1300
rect 7500 1220 7520 1280
rect 7580 1220 7620 1280
rect 7680 1220 7720 1280
rect 7780 1220 7800 1280
rect 7500 1180 7800 1220
rect 7500 1120 7520 1180
rect 7580 1120 7620 1180
rect 7680 1120 7720 1180
rect 7780 1120 7800 1180
rect 7500 1080 7800 1120
rect 7500 1020 7520 1080
rect 7580 1020 7620 1080
rect 7680 1020 7720 1080
rect 7780 1020 7800 1080
rect 7500 1000 7800 1020
rect 4200 140 4500 260
rect 4200 60 4300 140
rect 4380 60 4500 140
rect 1300 -20 1400 0
rect 1300 -80 1320 -20
rect 1380 -80 1400 -20
rect 1300 -100 1400 -80
rect 4200 -220 4500 60
rect 4200 -280 4220 -220
rect 4280 -280 4320 -220
rect 4380 -280 4420 -220
rect 4480 -280 4500 -220
rect 4200 -320 4500 -280
rect 4200 -380 4220 -320
rect 4280 -380 4320 -320
rect 4380 -380 4420 -320
rect 4480 -380 4500 -320
rect 4200 -420 4500 -380
rect 4200 -480 4220 -420
rect 4280 -480 4320 -420
rect 4380 -480 4420 -420
rect 4480 -480 4500 -420
rect 4200 -500 4500 -480
<< via1 >>
rect 920 1220 980 1280
rect 1020 1220 1080 1280
rect 1120 1220 1180 1280
rect 920 1120 980 1180
rect 1020 1120 1080 1180
rect 1120 1120 1180 1180
rect 920 1020 980 1080
rect 1020 1020 1080 1080
rect 1120 1020 1180 1080
rect 2420 1220 2480 1280
rect 2520 1220 2580 1280
rect 2420 1120 2480 1180
rect 2520 1120 2580 1180
rect 2420 1020 2480 1080
rect 2520 1020 2580 1080
rect 3620 1220 3680 1280
rect 3720 1220 3780 1280
rect 3620 1120 3680 1180
rect 3720 1120 3780 1180
rect 3620 1020 3680 1080
rect 3720 1020 3780 1080
rect 4880 1220 4940 1280
rect 4980 1220 5040 1280
rect 4880 1120 4940 1180
rect 4980 1120 5040 1180
rect 4880 1020 4940 1080
rect 4980 1020 5040 1080
rect 6120 1220 6180 1280
rect 6220 1220 6280 1280
rect 6120 1120 6180 1180
rect 6220 1120 6280 1180
rect 6120 1020 6180 1080
rect 6220 1020 6280 1080
rect 7520 1220 7580 1280
rect 7620 1220 7680 1280
rect 7720 1220 7780 1280
rect 7520 1120 7580 1180
rect 7620 1120 7680 1180
rect 7720 1120 7780 1180
rect 7520 1020 7580 1080
rect 7620 1020 7680 1080
rect 7720 1020 7780 1080
<< metal2 >>
rect 900 1280 7800 1300
rect 900 1220 920 1280
rect 980 1220 1020 1280
rect 1080 1220 1120 1280
rect 1180 1220 2420 1280
rect 2480 1220 2520 1280
rect 2580 1220 3620 1280
rect 3680 1220 3720 1280
rect 3780 1220 4880 1280
rect 4940 1220 4980 1280
rect 5040 1220 6120 1280
rect 6180 1220 6220 1280
rect 6280 1220 7520 1280
rect 7580 1220 7620 1280
rect 7680 1220 7720 1280
rect 7780 1220 7800 1280
rect 900 1180 7800 1220
rect 900 1120 920 1180
rect 980 1120 1020 1180
rect 1080 1120 1120 1180
rect 1180 1120 2420 1180
rect 2480 1120 2520 1180
rect 2580 1120 3620 1180
rect 3680 1120 3720 1180
rect 3780 1120 4880 1180
rect 4940 1120 4980 1180
rect 5040 1120 6120 1180
rect 6180 1120 6220 1180
rect 6280 1120 7520 1180
rect 7580 1120 7620 1180
rect 7680 1120 7720 1180
rect 7780 1120 7800 1180
rect 900 1080 7800 1120
rect 900 1020 920 1080
rect 980 1020 1020 1080
rect 1080 1020 1120 1080
rect 1180 1020 2420 1080
rect 2480 1020 2520 1080
rect 2580 1020 3620 1080
rect 3680 1020 3720 1080
rect 3780 1020 4880 1080
rect 4940 1020 4980 1080
rect 5040 1020 6120 1080
rect 6180 1020 6220 1080
rect 6280 1020 7520 1080
rect 7580 1020 7620 1080
rect 7680 1020 7720 1080
rect 7780 1020 7800 1080
rect 900 1000 7800 1020
use sky130_fd_pr__pfet_g5v0d10v5_ZPXM7F  XM2
timestamp 1769999431
transform 1 0 4337 0 1 1104
box -2867 -1004 2867 1042
<< labels >>
flabel metal1 1300 -100 1400 0 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1000 1100 1100 1200 0 FreeSans 256 0 0 0 D2
port 2 nsew
flabel metal1 4300 -400 4400 -300 0 FreeSans 256 0 0 0 D1
port 1 nsew
<< end >>
