magic
tech sky130A
magscale 1 2
timestamp 1769169801
<< nwell >>
rect -1461 -2415 1461 2415
<< mvpmos >>
rect -1203 118 -953 2118
rect -895 118 -645 2118
rect -587 118 -337 2118
rect -279 118 -29 2118
rect 29 118 279 2118
rect 337 118 587 2118
rect 645 118 895 2118
rect 953 118 1203 2118
rect -1203 -2118 -953 -118
rect -895 -2118 -645 -118
rect -587 -2118 -337 -118
rect -279 -2118 -29 -118
rect 29 -2118 279 -118
rect 337 -2118 587 -118
rect 645 -2118 895 -118
rect 953 -2118 1203 -118
<< mvpdiff >>
rect -1261 2106 -1203 2118
rect -1261 130 -1249 2106
rect -1215 130 -1203 2106
rect -1261 118 -1203 130
rect -953 2106 -895 2118
rect -953 130 -941 2106
rect -907 130 -895 2106
rect -953 118 -895 130
rect -645 2106 -587 2118
rect -645 130 -633 2106
rect -599 130 -587 2106
rect -645 118 -587 130
rect -337 2106 -279 2118
rect -337 130 -325 2106
rect -291 130 -279 2106
rect -337 118 -279 130
rect -29 2106 29 2118
rect -29 130 -17 2106
rect 17 130 29 2106
rect -29 118 29 130
rect 279 2106 337 2118
rect 279 130 291 2106
rect 325 130 337 2106
rect 279 118 337 130
rect 587 2106 645 2118
rect 587 130 599 2106
rect 633 130 645 2106
rect 587 118 645 130
rect 895 2106 953 2118
rect 895 130 907 2106
rect 941 130 953 2106
rect 895 118 953 130
rect 1203 2106 1261 2118
rect 1203 130 1215 2106
rect 1249 130 1261 2106
rect 1203 118 1261 130
rect -1261 -130 -1203 -118
rect -1261 -2106 -1249 -130
rect -1215 -2106 -1203 -130
rect -1261 -2118 -1203 -2106
rect -953 -130 -895 -118
rect -953 -2106 -941 -130
rect -907 -2106 -895 -130
rect -953 -2118 -895 -2106
rect -645 -130 -587 -118
rect -645 -2106 -633 -130
rect -599 -2106 -587 -130
rect -645 -2118 -587 -2106
rect -337 -130 -279 -118
rect -337 -2106 -325 -130
rect -291 -2106 -279 -130
rect -337 -2118 -279 -2106
rect -29 -130 29 -118
rect -29 -2106 -17 -130
rect 17 -2106 29 -130
rect -29 -2118 29 -2106
rect 279 -130 337 -118
rect 279 -2106 291 -130
rect 325 -2106 337 -130
rect 279 -2118 337 -2106
rect 587 -130 645 -118
rect 587 -2106 599 -130
rect 633 -2106 645 -130
rect 587 -2118 645 -2106
rect 895 -130 953 -118
rect 895 -2106 907 -130
rect 941 -2106 953 -130
rect 895 -2118 953 -2106
rect 1203 -130 1261 -118
rect 1203 -2106 1215 -130
rect 1249 -2106 1261 -130
rect 1203 -2118 1261 -2106
<< mvpdiffc >>
rect -1249 130 -1215 2106
rect -941 130 -907 2106
rect -633 130 -599 2106
rect -325 130 -291 2106
rect -17 130 17 2106
rect 291 130 325 2106
rect 599 130 633 2106
rect 907 130 941 2106
rect 1215 130 1249 2106
rect -1249 -2106 -1215 -130
rect -941 -2106 -907 -130
rect -633 -2106 -599 -130
rect -325 -2106 -291 -130
rect -17 -2106 17 -130
rect 291 -2106 325 -130
rect 599 -2106 633 -130
rect 907 -2106 941 -130
rect 1215 -2106 1249 -130
<< mvnsubdiff >>
rect -1395 2337 1395 2349
rect -1395 2303 -1287 2337
rect 1287 2303 1395 2337
rect -1395 2291 1395 2303
rect -1395 2241 -1337 2291
rect -1395 -2241 -1383 2241
rect -1349 -2241 -1337 2241
rect 1337 2241 1395 2291
rect -1395 -2291 -1337 -2241
rect 1337 -2241 1349 2241
rect 1383 -2241 1395 2241
rect 1337 -2291 1395 -2241
rect -1395 -2303 1395 -2291
rect -1395 -2337 -1287 -2303
rect 1287 -2337 1395 -2303
rect -1395 -2349 1395 -2337
<< mvnsubdiffcont >>
rect -1287 2303 1287 2337
rect -1383 -2241 -1349 2241
rect 1349 -2241 1383 2241
rect -1287 -2337 1287 -2303
<< poly >>
rect -1203 2199 -953 2215
rect -1203 2165 -1187 2199
rect -969 2165 -953 2199
rect -1203 2118 -953 2165
rect -895 2199 -645 2215
rect -895 2165 -879 2199
rect -661 2165 -645 2199
rect -895 2118 -645 2165
rect -587 2199 -337 2215
rect -587 2165 -571 2199
rect -353 2165 -337 2199
rect -587 2118 -337 2165
rect -279 2199 -29 2215
rect -279 2165 -263 2199
rect -45 2165 -29 2199
rect -279 2118 -29 2165
rect 29 2199 279 2215
rect 29 2165 45 2199
rect 263 2165 279 2199
rect 29 2118 279 2165
rect 337 2199 587 2215
rect 337 2165 353 2199
rect 571 2165 587 2199
rect 337 2118 587 2165
rect 645 2199 895 2215
rect 645 2165 661 2199
rect 879 2165 895 2199
rect 645 2118 895 2165
rect 953 2199 1203 2215
rect 953 2165 969 2199
rect 1187 2165 1203 2199
rect 953 2118 1203 2165
rect -1203 71 -953 118
rect -1203 37 -1187 71
rect -969 37 -953 71
rect -1203 21 -953 37
rect -895 71 -645 118
rect -895 37 -879 71
rect -661 37 -645 71
rect -895 21 -645 37
rect -587 71 -337 118
rect -587 37 -571 71
rect -353 37 -337 71
rect -587 21 -337 37
rect -279 71 -29 118
rect -279 37 -263 71
rect -45 37 -29 71
rect -279 21 -29 37
rect 29 71 279 118
rect 29 37 45 71
rect 263 37 279 71
rect 29 21 279 37
rect 337 71 587 118
rect 337 37 353 71
rect 571 37 587 71
rect 337 21 587 37
rect 645 71 895 118
rect 645 37 661 71
rect 879 37 895 71
rect 645 21 895 37
rect 953 71 1203 118
rect 953 37 969 71
rect 1187 37 1203 71
rect 953 21 1203 37
rect -1203 -37 -953 -21
rect -1203 -71 -1187 -37
rect -969 -71 -953 -37
rect -1203 -118 -953 -71
rect -895 -37 -645 -21
rect -895 -71 -879 -37
rect -661 -71 -645 -37
rect -895 -118 -645 -71
rect -587 -37 -337 -21
rect -587 -71 -571 -37
rect -353 -71 -337 -37
rect -587 -118 -337 -71
rect -279 -37 -29 -21
rect -279 -71 -263 -37
rect -45 -71 -29 -37
rect -279 -118 -29 -71
rect 29 -37 279 -21
rect 29 -71 45 -37
rect 263 -71 279 -37
rect 29 -118 279 -71
rect 337 -37 587 -21
rect 337 -71 353 -37
rect 571 -71 587 -37
rect 337 -118 587 -71
rect 645 -37 895 -21
rect 645 -71 661 -37
rect 879 -71 895 -37
rect 645 -118 895 -71
rect 953 -37 1203 -21
rect 953 -71 969 -37
rect 1187 -71 1203 -37
rect 953 -118 1203 -71
rect -1203 -2165 -953 -2118
rect -1203 -2199 -1187 -2165
rect -969 -2199 -953 -2165
rect -1203 -2215 -953 -2199
rect -895 -2165 -645 -2118
rect -895 -2199 -879 -2165
rect -661 -2199 -645 -2165
rect -895 -2215 -645 -2199
rect -587 -2165 -337 -2118
rect -587 -2199 -571 -2165
rect -353 -2199 -337 -2165
rect -587 -2215 -337 -2199
rect -279 -2165 -29 -2118
rect -279 -2199 -263 -2165
rect -45 -2199 -29 -2165
rect -279 -2215 -29 -2199
rect 29 -2165 279 -2118
rect 29 -2199 45 -2165
rect 263 -2199 279 -2165
rect 29 -2215 279 -2199
rect 337 -2165 587 -2118
rect 337 -2199 353 -2165
rect 571 -2199 587 -2165
rect 337 -2215 587 -2199
rect 645 -2165 895 -2118
rect 645 -2199 661 -2165
rect 879 -2199 895 -2165
rect 645 -2215 895 -2199
rect 953 -2165 1203 -2118
rect 953 -2199 969 -2165
rect 1187 -2199 1203 -2165
rect 953 -2215 1203 -2199
<< polycont >>
rect -1187 2165 -969 2199
rect -879 2165 -661 2199
rect -571 2165 -353 2199
rect -263 2165 -45 2199
rect 45 2165 263 2199
rect 353 2165 571 2199
rect 661 2165 879 2199
rect 969 2165 1187 2199
rect -1187 37 -969 71
rect -879 37 -661 71
rect -571 37 -353 71
rect -263 37 -45 71
rect 45 37 263 71
rect 353 37 571 71
rect 661 37 879 71
rect 969 37 1187 71
rect -1187 -71 -969 -37
rect -879 -71 -661 -37
rect -571 -71 -353 -37
rect -263 -71 -45 -37
rect 45 -71 263 -37
rect 353 -71 571 -37
rect 661 -71 879 -37
rect 969 -71 1187 -37
rect -1187 -2199 -969 -2165
rect -879 -2199 -661 -2165
rect -571 -2199 -353 -2165
rect -263 -2199 -45 -2165
rect 45 -2199 263 -2165
rect 353 -2199 571 -2165
rect 661 -2199 879 -2165
rect 969 -2199 1187 -2165
<< locali >>
rect -1383 2303 -1287 2337
rect 1287 2303 1383 2337
rect -1383 2241 -1349 2303
rect 1349 2241 1383 2303
rect -1203 2165 -1187 2199
rect -969 2165 -953 2199
rect -895 2165 -879 2199
rect -661 2165 -645 2199
rect -587 2165 -571 2199
rect -353 2165 -337 2199
rect -279 2165 -263 2199
rect -45 2165 -29 2199
rect 29 2165 45 2199
rect 263 2165 279 2199
rect 337 2165 353 2199
rect 571 2165 587 2199
rect 645 2165 661 2199
rect 879 2165 895 2199
rect 953 2165 969 2199
rect 1187 2165 1203 2199
rect -1249 2106 -1215 2122
rect -1249 114 -1215 130
rect -941 2106 -907 2122
rect -941 114 -907 130
rect -633 2106 -599 2122
rect -633 114 -599 130
rect -325 2106 -291 2122
rect -325 114 -291 130
rect -17 2106 17 2122
rect -17 114 17 130
rect 291 2106 325 2122
rect 291 114 325 130
rect 599 2106 633 2122
rect 599 114 633 130
rect 907 2106 941 2122
rect 907 114 941 130
rect 1215 2106 1249 2122
rect 1215 114 1249 130
rect -1203 37 -1187 71
rect -969 37 -953 71
rect -895 37 -879 71
rect -661 37 -645 71
rect -587 37 -571 71
rect -353 37 -337 71
rect -279 37 -263 71
rect -45 37 -29 71
rect 29 37 45 71
rect 263 37 279 71
rect 337 37 353 71
rect 571 37 587 71
rect 645 37 661 71
rect 879 37 895 71
rect 953 37 969 71
rect 1187 37 1203 71
rect -1203 -71 -1187 -37
rect -969 -71 -953 -37
rect -895 -71 -879 -37
rect -661 -71 -645 -37
rect -587 -71 -571 -37
rect -353 -71 -337 -37
rect -279 -71 -263 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 263 -71 279 -37
rect 337 -71 353 -37
rect 571 -71 587 -37
rect 645 -71 661 -37
rect 879 -71 895 -37
rect 953 -71 969 -37
rect 1187 -71 1203 -37
rect -1249 -130 -1215 -114
rect -1249 -2122 -1215 -2106
rect -941 -130 -907 -114
rect -941 -2122 -907 -2106
rect -633 -130 -599 -114
rect -633 -2122 -599 -2106
rect -325 -130 -291 -114
rect -325 -2122 -291 -2106
rect -17 -130 17 -114
rect -17 -2122 17 -2106
rect 291 -130 325 -114
rect 291 -2122 325 -2106
rect 599 -130 633 -114
rect 599 -2122 633 -2106
rect 907 -130 941 -114
rect 907 -2122 941 -2106
rect 1215 -130 1249 -114
rect 1215 -2122 1249 -2106
rect -1203 -2199 -1187 -2165
rect -969 -2199 -953 -2165
rect -895 -2199 -879 -2165
rect -661 -2199 -645 -2165
rect -587 -2199 -571 -2165
rect -353 -2199 -337 -2165
rect -279 -2199 -263 -2165
rect -45 -2199 -29 -2165
rect 29 -2199 45 -2165
rect 263 -2199 279 -2165
rect 337 -2199 353 -2165
rect 571 -2199 587 -2165
rect 645 -2199 661 -2165
rect 879 -2199 895 -2165
rect 953 -2199 969 -2165
rect 1187 -2199 1203 -2165
rect -1383 -2303 -1349 -2241
rect 1349 -2303 1383 -2241
rect -1383 -2337 -1287 -2303
rect 1287 -2337 1383 -2303
<< viali >>
rect -1187 2165 -969 2199
rect -879 2165 -661 2199
rect -571 2165 -353 2199
rect -263 2165 -45 2199
rect 45 2165 263 2199
rect 353 2165 571 2199
rect 661 2165 879 2199
rect 969 2165 1187 2199
rect -1249 130 -1215 2106
rect -941 130 -907 2106
rect -633 130 -599 2106
rect -325 130 -291 2106
rect -17 130 17 2106
rect 291 130 325 2106
rect 599 130 633 2106
rect 907 130 941 2106
rect 1215 130 1249 2106
rect -1187 37 -969 71
rect -879 37 -661 71
rect -571 37 -353 71
rect -263 37 -45 71
rect 45 37 263 71
rect 353 37 571 71
rect 661 37 879 71
rect 969 37 1187 71
rect -1187 -71 -969 -37
rect -879 -71 -661 -37
rect -571 -71 -353 -37
rect -263 -71 -45 -37
rect 45 -71 263 -37
rect 353 -71 571 -37
rect 661 -71 879 -37
rect 969 -71 1187 -37
rect -1249 -2106 -1215 -130
rect -941 -2106 -907 -130
rect -633 -2106 -599 -130
rect -325 -2106 -291 -130
rect -17 -2106 17 -130
rect 291 -2106 325 -130
rect 599 -2106 633 -130
rect 907 -2106 941 -130
rect 1215 -2106 1249 -130
rect -1187 -2199 -969 -2165
rect -879 -2199 -661 -2165
rect -571 -2199 -353 -2165
rect -263 -2199 -45 -2165
rect 45 -2199 263 -2165
rect 353 -2199 571 -2165
rect 661 -2199 879 -2165
rect 969 -2199 1187 -2165
<< metal1 >>
rect -1199 2199 -957 2205
rect -1199 2165 -1187 2199
rect -969 2165 -957 2199
rect -1199 2159 -957 2165
rect -891 2199 -649 2205
rect -891 2165 -879 2199
rect -661 2165 -649 2199
rect -891 2159 -649 2165
rect -583 2199 -341 2205
rect -583 2165 -571 2199
rect -353 2165 -341 2199
rect -583 2159 -341 2165
rect -275 2199 -33 2205
rect -275 2165 -263 2199
rect -45 2165 -33 2199
rect -275 2159 -33 2165
rect 33 2199 275 2205
rect 33 2165 45 2199
rect 263 2165 275 2199
rect 33 2159 275 2165
rect 341 2199 583 2205
rect 341 2165 353 2199
rect 571 2165 583 2199
rect 341 2159 583 2165
rect 649 2199 891 2205
rect 649 2165 661 2199
rect 879 2165 891 2199
rect 649 2159 891 2165
rect 957 2199 1199 2205
rect 957 2165 969 2199
rect 1187 2165 1199 2199
rect 957 2159 1199 2165
rect -1255 2106 -1209 2118
rect -1255 130 -1249 2106
rect -1215 130 -1209 2106
rect -1255 118 -1209 130
rect -947 2106 -901 2118
rect -947 130 -941 2106
rect -907 130 -901 2106
rect -947 118 -901 130
rect -639 2106 -593 2118
rect -639 130 -633 2106
rect -599 130 -593 2106
rect -639 118 -593 130
rect -331 2106 -285 2118
rect -331 130 -325 2106
rect -291 130 -285 2106
rect -331 118 -285 130
rect -23 2106 23 2118
rect -23 130 -17 2106
rect 17 130 23 2106
rect -23 118 23 130
rect 285 2106 331 2118
rect 285 130 291 2106
rect 325 130 331 2106
rect 285 118 331 130
rect 593 2106 639 2118
rect 593 130 599 2106
rect 633 130 639 2106
rect 593 118 639 130
rect 901 2106 947 2118
rect 901 130 907 2106
rect 941 130 947 2106
rect 901 118 947 130
rect 1209 2106 1255 2118
rect 1209 130 1215 2106
rect 1249 130 1255 2106
rect 1209 118 1255 130
rect -1199 71 -957 77
rect -1199 37 -1187 71
rect -969 37 -957 71
rect -1199 31 -957 37
rect -891 71 -649 77
rect -891 37 -879 71
rect -661 37 -649 71
rect -891 31 -649 37
rect -583 71 -341 77
rect -583 37 -571 71
rect -353 37 -341 71
rect -583 31 -341 37
rect -275 71 -33 77
rect -275 37 -263 71
rect -45 37 -33 71
rect -275 31 -33 37
rect 33 71 275 77
rect 33 37 45 71
rect 263 37 275 71
rect 33 31 275 37
rect 341 71 583 77
rect 341 37 353 71
rect 571 37 583 71
rect 341 31 583 37
rect 649 71 891 77
rect 649 37 661 71
rect 879 37 891 71
rect 649 31 891 37
rect 957 71 1199 77
rect 957 37 969 71
rect 1187 37 1199 71
rect 957 31 1199 37
rect -1199 -37 -957 -31
rect -1199 -71 -1187 -37
rect -969 -71 -957 -37
rect -1199 -77 -957 -71
rect -891 -37 -649 -31
rect -891 -71 -879 -37
rect -661 -71 -649 -37
rect -891 -77 -649 -71
rect -583 -37 -341 -31
rect -583 -71 -571 -37
rect -353 -71 -341 -37
rect -583 -77 -341 -71
rect -275 -37 -33 -31
rect -275 -71 -263 -37
rect -45 -71 -33 -37
rect -275 -77 -33 -71
rect 33 -37 275 -31
rect 33 -71 45 -37
rect 263 -71 275 -37
rect 33 -77 275 -71
rect 341 -37 583 -31
rect 341 -71 353 -37
rect 571 -71 583 -37
rect 341 -77 583 -71
rect 649 -37 891 -31
rect 649 -71 661 -37
rect 879 -71 891 -37
rect 649 -77 891 -71
rect 957 -37 1199 -31
rect 957 -71 969 -37
rect 1187 -71 1199 -37
rect 957 -77 1199 -71
rect -1255 -130 -1209 -118
rect -1255 -2106 -1249 -130
rect -1215 -2106 -1209 -130
rect -1255 -2118 -1209 -2106
rect -947 -130 -901 -118
rect -947 -2106 -941 -130
rect -907 -2106 -901 -130
rect -947 -2118 -901 -2106
rect -639 -130 -593 -118
rect -639 -2106 -633 -130
rect -599 -2106 -593 -130
rect -639 -2118 -593 -2106
rect -331 -130 -285 -118
rect -331 -2106 -325 -130
rect -291 -2106 -285 -130
rect -331 -2118 -285 -2106
rect -23 -130 23 -118
rect -23 -2106 -17 -130
rect 17 -2106 23 -130
rect -23 -2118 23 -2106
rect 285 -130 331 -118
rect 285 -2106 291 -130
rect 325 -2106 331 -130
rect 285 -2118 331 -2106
rect 593 -130 639 -118
rect 593 -2106 599 -130
rect 633 -2106 639 -130
rect 593 -2118 639 -2106
rect 901 -130 947 -118
rect 901 -2106 907 -130
rect 941 -2106 947 -130
rect 901 -2118 947 -2106
rect 1209 -130 1255 -118
rect 1209 -2106 1215 -130
rect 1249 -2106 1255 -130
rect 1209 -2118 1255 -2106
rect -1199 -2165 -957 -2159
rect -1199 -2199 -1187 -2165
rect -969 -2199 -957 -2165
rect -1199 -2205 -957 -2199
rect -891 -2165 -649 -2159
rect -891 -2199 -879 -2165
rect -661 -2199 -649 -2165
rect -891 -2205 -649 -2199
rect -583 -2165 -341 -2159
rect -583 -2199 -571 -2165
rect -353 -2199 -341 -2165
rect -583 -2205 -341 -2199
rect -275 -2165 -33 -2159
rect -275 -2199 -263 -2165
rect -45 -2199 -33 -2165
rect -275 -2205 -33 -2199
rect 33 -2165 275 -2159
rect 33 -2199 45 -2165
rect 263 -2199 275 -2165
rect 33 -2205 275 -2199
rect 341 -2165 583 -2159
rect 341 -2199 353 -2165
rect 571 -2199 583 -2165
rect 341 -2205 583 -2199
rect 649 -2165 891 -2159
rect 649 -2199 661 -2165
rect 879 -2199 891 -2165
rect 649 -2205 891 -2199
rect 957 -2165 1199 -2159
rect 957 -2199 969 -2165
rect 1187 -2199 1199 -2165
rect 957 -2205 1199 -2199
<< properties >>
string FIXED_BBOX -1366 -2320 1366 2320
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 1.25 m 2 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
