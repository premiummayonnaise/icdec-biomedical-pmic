magic
tech sky130A
magscale 1 2
timestamp 1769411983
<< pwell >>
rect -1463 -729 1463 729
<< mvnmos >>
rect -1235 -471 -1135 471
rect -1077 -471 -977 471
rect -919 -471 -819 471
rect -761 -471 -661 471
rect -603 -471 -503 471
rect -445 -471 -345 471
rect -287 -471 -187 471
rect -129 -471 -29 471
rect 29 -471 129 471
rect 187 -471 287 471
rect 345 -471 445 471
rect 503 -471 603 471
rect 661 -471 761 471
rect 819 -471 919 471
rect 977 -471 1077 471
rect 1135 -471 1235 471
<< mvndiff >>
rect -1293 459 -1235 471
rect -1293 -459 -1281 459
rect -1247 -459 -1235 459
rect -1293 -471 -1235 -459
rect -1135 459 -1077 471
rect -1135 -459 -1123 459
rect -1089 -459 -1077 459
rect -1135 -471 -1077 -459
rect -977 459 -919 471
rect -977 -459 -965 459
rect -931 -459 -919 459
rect -977 -471 -919 -459
rect -819 459 -761 471
rect -819 -459 -807 459
rect -773 -459 -761 459
rect -819 -471 -761 -459
rect -661 459 -603 471
rect -661 -459 -649 459
rect -615 -459 -603 459
rect -661 -471 -603 -459
rect -503 459 -445 471
rect -503 -459 -491 459
rect -457 -459 -445 459
rect -503 -471 -445 -459
rect -345 459 -287 471
rect -345 -459 -333 459
rect -299 -459 -287 459
rect -345 -471 -287 -459
rect -187 459 -129 471
rect -187 -459 -175 459
rect -141 -459 -129 459
rect -187 -471 -129 -459
rect -29 459 29 471
rect -29 -459 -17 459
rect 17 -459 29 459
rect -29 -471 29 -459
rect 129 459 187 471
rect 129 -459 141 459
rect 175 -459 187 459
rect 129 -471 187 -459
rect 287 459 345 471
rect 287 -459 299 459
rect 333 -459 345 459
rect 287 -471 345 -459
rect 445 459 503 471
rect 445 -459 457 459
rect 491 -459 503 459
rect 445 -471 503 -459
rect 603 459 661 471
rect 603 -459 615 459
rect 649 -459 661 459
rect 603 -471 661 -459
rect 761 459 819 471
rect 761 -459 773 459
rect 807 -459 819 459
rect 761 -471 819 -459
rect 919 459 977 471
rect 919 -459 931 459
rect 965 -459 977 459
rect 919 -471 977 -459
rect 1077 459 1135 471
rect 1077 -459 1089 459
rect 1123 -459 1135 459
rect 1077 -471 1135 -459
rect 1235 459 1293 471
rect 1235 -459 1247 459
rect 1281 -459 1293 459
rect 1235 -471 1293 -459
<< mvndiffc >>
rect -1281 -459 -1247 459
rect -1123 -459 -1089 459
rect -965 -459 -931 459
rect -807 -459 -773 459
rect -649 -459 -615 459
rect -491 -459 -457 459
rect -333 -459 -299 459
rect -175 -459 -141 459
rect -17 -459 17 459
rect 141 -459 175 459
rect 299 -459 333 459
rect 457 -459 491 459
rect 615 -459 649 459
rect 773 -459 807 459
rect 931 -459 965 459
rect 1089 -459 1123 459
rect 1247 -459 1281 459
<< mvpsubdiff >>
rect -1427 681 1427 693
rect -1427 647 -1319 681
rect 1319 647 1427 681
rect -1427 635 1427 647
rect -1427 585 -1369 635
rect -1427 -585 -1415 585
rect -1381 -585 -1369 585
rect 1369 585 1427 635
rect -1427 -635 -1369 -585
rect 1369 -585 1381 585
rect 1415 -585 1427 585
rect 1369 -635 1427 -585
rect -1427 -647 1427 -635
rect -1427 -681 -1319 -647
rect 1319 -681 1427 -647
rect -1427 -693 1427 -681
<< mvpsubdiffcont >>
rect -1319 647 1319 681
rect -1415 -585 -1381 585
rect 1381 -585 1415 585
rect -1319 -681 1319 -647
<< poly >>
rect -1235 543 -1135 559
rect -1235 509 -1219 543
rect -1151 509 -1135 543
rect -1235 471 -1135 509
rect -1077 543 -977 559
rect -1077 509 -1061 543
rect -993 509 -977 543
rect -1077 471 -977 509
rect -919 543 -819 559
rect -919 509 -903 543
rect -835 509 -819 543
rect -919 471 -819 509
rect -761 543 -661 559
rect -761 509 -745 543
rect -677 509 -661 543
rect -761 471 -661 509
rect -603 543 -503 559
rect -603 509 -587 543
rect -519 509 -503 543
rect -603 471 -503 509
rect -445 543 -345 559
rect -445 509 -429 543
rect -361 509 -345 543
rect -445 471 -345 509
rect -287 543 -187 559
rect -287 509 -271 543
rect -203 509 -187 543
rect -287 471 -187 509
rect -129 543 -29 559
rect -129 509 -113 543
rect -45 509 -29 543
rect -129 471 -29 509
rect 29 543 129 559
rect 29 509 45 543
rect 113 509 129 543
rect 29 471 129 509
rect 187 543 287 559
rect 187 509 203 543
rect 271 509 287 543
rect 187 471 287 509
rect 345 543 445 559
rect 345 509 361 543
rect 429 509 445 543
rect 345 471 445 509
rect 503 543 603 559
rect 503 509 519 543
rect 587 509 603 543
rect 503 471 603 509
rect 661 543 761 559
rect 661 509 677 543
rect 745 509 761 543
rect 661 471 761 509
rect 819 543 919 559
rect 819 509 835 543
rect 903 509 919 543
rect 819 471 919 509
rect 977 543 1077 559
rect 977 509 993 543
rect 1061 509 1077 543
rect 977 471 1077 509
rect 1135 543 1235 559
rect 1135 509 1151 543
rect 1219 509 1235 543
rect 1135 471 1235 509
rect -1235 -509 -1135 -471
rect -1235 -543 -1219 -509
rect -1151 -543 -1135 -509
rect -1235 -559 -1135 -543
rect -1077 -509 -977 -471
rect -1077 -543 -1061 -509
rect -993 -543 -977 -509
rect -1077 -559 -977 -543
rect -919 -509 -819 -471
rect -919 -543 -903 -509
rect -835 -543 -819 -509
rect -919 -559 -819 -543
rect -761 -509 -661 -471
rect -761 -543 -745 -509
rect -677 -543 -661 -509
rect -761 -559 -661 -543
rect -603 -509 -503 -471
rect -603 -543 -587 -509
rect -519 -543 -503 -509
rect -603 -559 -503 -543
rect -445 -509 -345 -471
rect -445 -543 -429 -509
rect -361 -543 -345 -509
rect -445 -559 -345 -543
rect -287 -509 -187 -471
rect -287 -543 -271 -509
rect -203 -543 -187 -509
rect -287 -559 -187 -543
rect -129 -509 -29 -471
rect -129 -543 -113 -509
rect -45 -543 -29 -509
rect -129 -559 -29 -543
rect 29 -509 129 -471
rect 29 -543 45 -509
rect 113 -543 129 -509
rect 29 -559 129 -543
rect 187 -509 287 -471
rect 187 -543 203 -509
rect 271 -543 287 -509
rect 187 -559 287 -543
rect 345 -509 445 -471
rect 345 -543 361 -509
rect 429 -543 445 -509
rect 345 -559 445 -543
rect 503 -509 603 -471
rect 503 -543 519 -509
rect 587 -543 603 -509
rect 503 -559 603 -543
rect 661 -509 761 -471
rect 661 -543 677 -509
rect 745 -543 761 -509
rect 661 -559 761 -543
rect 819 -509 919 -471
rect 819 -543 835 -509
rect 903 -543 919 -509
rect 819 -559 919 -543
rect 977 -509 1077 -471
rect 977 -543 993 -509
rect 1061 -543 1077 -509
rect 977 -559 1077 -543
rect 1135 -509 1235 -471
rect 1135 -543 1151 -509
rect 1219 -543 1235 -509
rect 1135 -559 1235 -543
<< polycont >>
rect -1219 509 -1151 543
rect -1061 509 -993 543
rect -903 509 -835 543
rect -745 509 -677 543
rect -587 509 -519 543
rect -429 509 -361 543
rect -271 509 -203 543
rect -113 509 -45 543
rect 45 509 113 543
rect 203 509 271 543
rect 361 509 429 543
rect 519 509 587 543
rect 677 509 745 543
rect 835 509 903 543
rect 993 509 1061 543
rect 1151 509 1219 543
rect -1219 -543 -1151 -509
rect -1061 -543 -993 -509
rect -903 -543 -835 -509
rect -745 -543 -677 -509
rect -587 -543 -519 -509
rect -429 -543 -361 -509
rect -271 -543 -203 -509
rect -113 -543 -45 -509
rect 45 -543 113 -509
rect 203 -543 271 -509
rect 361 -543 429 -509
rect 519 -543 587 -509
rect 677 -543 745 -509
rect 835 -543 903 -509
rect 993 -543 1061 -509
rect 1151 -543 1219 -509
<< locali >>
rect -1415 647 -1319 681
rect 1319 647 1415 681
rect -1415 585 -1381 647
rect 1381 585 1415 647
rect -1235 509 -1219 543
rect -1151 509 -1135 543
rect -1077 509 -1061 543
rect -993 509 -977 543
rect -919 509 -903 543
rect -835 509 -819 543
rect -761 509 -745 543
rect -677 509 -661 543
rect -603 509 -587 543
rect -519 509 -503 543
rect -445 509 -429 543
rect -361 509 -345 543
rect -287 509 -271 543
rect -203 509 -187 543
rect -129 509 -113 543
rect -45 509 -29 543
rect 29 509 45 543
rect 113 509 129 543
rect 187 509 203 543
rect 271 509 287 543
rect 345 509 361 543
rect 429 509 445 543
rect 503 509 519 543
rect 587 509 603 543
rect 661 509 677 543
rect 745 509 761 543
rect 819 509 835 543
rect 903 509 919 543
rect 977 509 993 543
rect 1061 509 1077 543
rect 1135 509 1151 543
rect 1219 509 1235 543
rect -1281 459 -1247 475
rect -1281 -475 -1247 -459
rect -1123 459 -1089 475
rect -1123 -475 -1089 -459
rect -965 459 -931 475
rect -965 -475 -931 -459
rect -807 459 -773 475
rect -807 -475 -773 -459
rect -649 459 -615 475
rect -649 -475 -615 -459
rect -491 459 -457 475
rect -491 -475 -457 -459
rect -333 459 -299 475
rect -333 -475 -299 -459
rect -175 459 -141 475
rect -175 -475 -141 -459
rect -17 459 17 475
rect -17 -475 17 -459
rect 141 459 175 475
rect 141 -475 175 -459
rect 299 459 333 475
rect 299 -475 333 -459
rect 457 459 491 475
rect 457 -475 491 -459
rect 615 459 649 475
rect 615 -475 649 -459
rect 773 459 807 475
rect 773 -475 807 -459
rect 931 459 965 475
rect 931 -475 965 -459
rect 1089 459 1123 475
rect 1089 -475 1123 -459
rect 1247 459 1281 475
rect 1247 -475 1281 -459
rect -1235 -543 -1219 -509
rect -1151 -543 -1135 -509
rect -1077 -543 -1061 -509
rect -993 -543 -977 -509
rect -919 -543 -903 -509
rect -835 -543 -819 -509
rect -761 -543 -745 -509
rect -677 -543 -661 -509
rect -603 -543 -587 -509
rect -519 -543 -503 -509
rect -445 -543 -429 -509
rect -361 -543 -345 -509
rect -287 -543 -271 -509
rect -203 -543 -187 -509
rect -129 -543 -113 -509
rect -45 -543 -29 -509
rect 29 -543 45 -509
rect 113 -543 129 -509
rect 187 -543 203 -509
rect 271 -543 287 -509
rect 345 -543 361 -509
rect 429 -543 445 -509
rect 503 -543 519 -509
rect 587 -543 603 -509
rect 661 -543 677 -509
rect 745 -543 761 -509
rect 819 -543 835 -509
rect 903 -543 919 -509
rect 977 -543 993 -509
rect 1061 -543 1077 -509
rect 1135 -543 1151 -509
rect 1219 -543 1235 -509
rect -1415 -647 -1381 -585
rect 1381 -647 1415 -585
rect -1415 -681 -1319 -647
rect 1319 -681 1415 -647
<< viali >>
rect -1219 509 -1151 543
rect -1061 509 -993 543
rect -903 509 -835 543
rect -745 509 -677 543
rect -587 509 -519 543
rect -429 509 -361 543
rect -271 509 -203 543
rect -113 509 -45 543
rect 45 509 113 543
rect 203 509 271 543
rect 361 509 429 543
rect 519 509 587 543
rect 677 509 745 543
rect 835 509 903 543
rect 993 509 1061 543
rect 1151 509 1219 543
rect -1281 -459 -1247 459
rect -1123 -459 -1089 459
rect -965 -459 -931 459
rect -807 -459 -773 459
rect -649 -459 -615 459
rect -491 -459 -457 459
rect -333 -459 -299 459
rect -175 -459 -141 459
rect -17 -459 17 459
rect 141 -459 175 459
rect 299 -459 333 459
rect 457 -459 491 459
rect 615 -459 649 459
rect 773 -459 807 459
rect 931 -459 965 459
rect 1089 -459 1123 459
rect 1247 -459 1281 459
rect -1219 -543 -1151 -509
rect -1061 -543 -993 -509
rect -903 -543 -835 -509
rect -745 -543 -677 -509
rect -587 -543 -519 -509
rect -429 -543 -361 -509
rect -271 -543 -203 -509
rect -113 -543 -45 -509
rect 45 -543 113 -509
rect 203 -543 271 -509
rect 361 -543 429 -509
rect 519 -543 587 -509
rect 677 -543 745 -509
rect 835 -543 903 -509
rect 993 -543 1061 -509
rect 1151 -543 1219 -509
<< metal1 >>
rect -1231 543 -1139 549
rect -1231 509 -1219 543
rect -1151 509 -1139 543
rect -1231 503 -1139 509
rect -1073 543 -981 549
rect -1073 509 -1061 543
rect -993 509 -981 543
rect -1073 503 -981 509
rect -915 543 -823 549
rect -915 509 -903 543
rect -835 509 -823 543
rect -915 503 -823 509
rect -757 543 -665 549
rect -757 509 -745 543
rect -677 509 -665 543
rect -757 503 -665 509
rect -599 543 -507 549
rect -599 509 -587 543
rect -519 509 -507 543
rect -599 503 -507 509
rect -441 543 -349 549
rect -441 509 -429 543
rect -361 509 -349 543
rect -441 503 -349 509
rect -283 543 -191 549
rect -283 509 -271 543
rect -203 509 -191 543
rect -283 503 -191 509
rect -125 543 -33 549
rect -125 509 -113 543
rect -45 509 -33 543
rect -125 503 -33 509
rect 33 543 125 549
rect 33 509 45 543
rect 113 509 125 543
rect 33 503 125 509
rect 191 543 283 549
rect 191 509 203 543
rect 271 509 283 543
rect 191 503 283 509
rect 349 543 441 549
rect 349 509 361 543
rect 429 509 441 543
rect 349 503 441 509
rect 507 543 599 549
rect 507 509 519 543
rect 587 509 599 543
rect 507 503 599 509
rect 665 543 757 549
rect 665 509 677 543
rect 745 509 757 543
rect 665 503 757 509
rect 823 543 915 549
rect 823 509 835 543
rect 903 509 915 543
rect 823 503 915 509
rect 981 543 1073 549
rect 981 509 993 543
rect 1061 509 1073 543
rect 981 503 1073 509
rect 1139 543 1231 549
rect 1139 509 1151 543
rect 1219 509 1231 543
rect 1139 503 1231 509
rect -1287 459 -1241 471
rect -1287 -459 -1281 459
rect -1247 -459 -1241 459
rect -1287 -471 -1241 -459
rect -1129 459 -1083 471
rect -1129 -459 -1123 459
rect -1089 -459 -1083 459
rect -1129 -471 -1083 -459
rect -971 459 -925 471
rect -971 -459 -965 459
rect -931 -459 -925 459
rect -971 -471 -925 -459
rect -813 459 -767 471
rect -813 -459 -807 459
rect -773 -459 -767 459
rect -813 -471 -767 -459
rect -655 459 -609 471
rect -655 -459 -649 459
rect -615 -459 -609 459
rect -655 -471 -609 -459
rect -497 459 -451 471
rect -497 -459 -491 459
rect -457 -459 -451 459
rect -497 -471 -451 -459
rect -339 459 -293 471
rect -339 -459 -333 459
rect -299 -459 -293 459
rect -339 -471 -293 -459
rect -181 459 -135 471
rect -181 -459 -175 459
rect -141 -459 -135 459
rect -181 -471 -135 -459
rect -23 459 23 471
rect -23 -459 -17 459
rect 17 -459 23 459
rect -23 -471 23 -459
rect 135 459 181 471
rect 135 -459 141 459
rect 175 -459 181 459
rect 135 -471 181 -459
rect 293 459 339 471
rect 293 -459 299 459
rect 333 -459 339 459
rect 293 -471 339 -459
rect 451 459 497 471
rect 451 -459 457 459
rect 491 -459 497 459
rect 451 -471 497 -459
rect 609 459 655 471
rect 609 -459 615 459
rect 649 -459 655 459
rect 609 -471 655 -459
rect 767 459 813 471
rect 767 -459 773 459
rect 807 -459 813 459
rect 767 -471 813 -459
rect 925 459 971 471
rect 925 -459 931 459
rect 965 -459 971 459
rect 925 -471 971 -459
rect 1083 459 1129 471
rect 1083 -459 1089 459
rect 1123 -459 1129 459
rect 1083 -471 1129 -459
rect 1241 459 1287 471
rect 1241 -459 1247 459
rect 1281 -459 1287 459
rect 1241 -471 1287 -459
rect -1231 -509 -1139 -503
rect -1231 -543 -1219 -509
rect -1151 -543 -1139 -509
rect -1231 -549 -1139 -543
rect -1073 -509 -981 -503
rect -1073 -543 -1061 -509
rect -993 -543 -981 -509
rect -1073 -549 -981 -543
rect -915 -509 -823 -503
rect -915 -543 -903 -509
rect -835 -543 -823 -509
rect -915 -549 -823 -543
rect -757 -509 -665 -503
rect -757 -543 -745 -509
rect -677 -543 -665 -509
rect -757 -549 -665 -543
rect -599 -509 -507 -503
rect -599 -543 -587 -509
rect -519 -543 -507 -509
rect -599 -549 -507 -543
rect -441 -509 -349 -503
rect -441 -543 -429 -509
rect -361 -543 -349 -509
rect -441 -549 -349 -543
rect -283 -509 -191 -503
rect -283 -543 -271 -509
rect -203 -543 -191 -509
rect -283 -549 -191 -543
rect -125 -509 -33 -503
rect -125 -543 -113 -509
rect -45 -543 -33 -509
rect -125 -549 -33 -543
rect 33 -509 125 -503
rect 33 -543 45 -509
rect 113 -543 125 -509
rect 33 -549 125 -543
rect 191 -509 283 -503
rect 191 -543 203 -509
rect 271 -543 283 -509
rect 191 -549 283 -543
rect 349 -509 441 -503
rect 349 -543 361 -509
rect 429 -543 441 -509
rect 349 -549 441 -543
rect 507 -509 599 -503
rect 507 -543 519 -509
rect 587 -543 599 -509
rect 507 -549 599 -543
rect 665 -509 757 -503
rect 665 -543 677 -509
rect 745 -543 757 -509
rect 665 -549 757 -543
rect 823 -509 915 -503
rect 823 -543 835 -509
rect 903 -543 915 -509
rect 823 -549 915 -543
rect 981 -509 1073 -503
rect 981 -543 993 -509
rect 1061 -543 1073 -509
rect 981 -549 1073 -543
rect 1139 -509 1231 -503
rect 1139 -543 1151 -509
rect 1219 -543 1231 -509
rect 1139 -549 1231 -543
<< properties >>
string FIXED_BBOX -1398 -664 1398 664
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.7125 l 0.5 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
