magic
tech sky130A
magscale 1 2
timestamp 1770083657
<< pwell >>
rect -371 -470 371 532
<< mvnmos >>
rect -287 -444 -187 506
rect -129 -444 -29 506
rect 29 -444 129 506
rect 187 -444 287 506
<< mvndiff >>
rect -345 388 -287 506
rect -345 354 -333 388
rect -299 354 -287 388
rect -345 320 -287 354
rect -345 286 -333 320
rect -299 286 -287 320
rect -345 252 -287 286
rect -345 218 -333 252
rect -299 218 -287 252
rect -345 184 -287 218
rect -345 150 -333 184
rect -299 150 -287 184
rect -345 116 -287 150
rect -345 82 -333 116
rect -299 82 -287 116
rect -345 48 -287 82
rect -345 14 -333 48
rect -299 14 -287 48
rect -345 -20 -287 14
rect -345 -54 -333 -20
rect -299 -54 -287 -20
rect -345 -88 -287 -54
rect -345 -122 -333 -88
rect -299 -122 -287 -88
rect -345 -156 -287 -122
rect -345 -190 -333 -156
rect -299 -190 -287 -156
rect -345 -224 -287 -190
rect -345 -258 -333 -224
rect -299 -258 -287 -224
rect -345 -292 -287 -258
rect -345 -326 -333 -292
rect -299 -326 -287 -292
rect -345 -444 -287 -326
rect -187 388 -129 506
rect -187 354 -175 388
rect -141 354 -129 388
rect -187 320 -129 354
rect -187 286 -175 320
rect -141 286 -129 320
rect -187 252 -129 286
rect -187 218 -175 252
rect -141 218 -129 252
rect -187 184 -129 218
rect -187 150 -175 184
rect -141 150 -129 184
rect -187 116 -129 150
rect -187 82 -175 116
rect -141 82 -129 116
rect -187 48 -129 82
rect -187 14 -175 48
rect -141 14 -129 48
rect -187 -20 -129 14
rect -187 -54 -175 -20
rect -141 -54 -129 -20
rect -187 -88 -129 -54
rect -187 -122 -175 -88
rect -141 -122 -129 -88
rect -187 -156 -129 -122
rect -187 -190 -175 -156
rect -141 -190 -129 -156
rect -187 -224 -129 -190
rect -187 -258 -175 -224
rect -141 -258 -129 -224
rect -187 -292 -129 -258
rect -187 -326 -175 -292
rect -141 -326 -129 -292
rect -187 -444 -129 -326
rect -29 388 29 506
rect -29 354 -17 388
rect 17 354 29 388
rect -29 320 29 354
rect -29 286 -17 320
rect 17 286 29 320
rect -29 252 29 286
rect -29 218 -17 252
rect 17 218 29 252
rect -29 184 29 218
rect -29 150 -17 184
rect 17 150 29 184
rect -29 116 29 150
rect -29 82 -17 116
rect 17 82 29 116
rect -29 48 29 82
rect -29 14 -17 48
rect 17 14 29 48
rect -29 -20 29 14
rect -29 -54 -17 -20
rect 17 -54 29 -20
rect -29 -88 29 -54
rect -29 -122 -17 -88
rect 17 -122 29 -88
rect -29 -156 29 -122
rect -29 -190 -17 -156
rect 17 -190 29 -156
rect -29 -224 29 -190
rect -29 -258 -17 -224
rect 17 -258 29 -224
rect -29 -292 29 -258
rect -29 -326 -17 -292
rect 17 -326 29 -292
rect -29 -444 29 -326
rect 129 388 187 506
rect 129 354 141 388
rect 175 354 187 388
rect 129 320 187 354
rect 129 286 141 320
rect 175 286 187 320
rect 129 252 187 286
rect 129 218 141 252
rect 175 218 187 252
rect 129 184 187 218
rect 129 150 141 184
rect 175 150 187 184
rect 129 116 187 150
rect 129 82 141 116
rect 175 82 187 116
rect 129 48 187 82
rect 129 14 141 48
rect 175 14 187 48
rect 129 -20 187 14
rect 129 -54 141 -20
rect 175 -54 187 -20
rect 129 -88 187 -54
rect 129 -122 141 -88
rect 175 -122 187 -88
rect 129 -156 187 -122
rect 129 -190 141 -156
rect 175 -190 187 -156
rect 129 -224 187 -190
rect 129 -258 141 -224
rect 175 -258 187 -224
rect 129 -292 187 -258
rect 129 -326 141 -292
rect 175 -326 187 -292
rect 129 -444 187 -326
rect 287 388 345 506
rect 287 354 299 388
rect 333 354 345 388
rect 287 320 345 354
rect 287 286 299 320
rect 333 286 345 320
rect 287 252 345 286
rect 287 218 299 252
rect 333 218 345 252
rect 287 184 345 218
rect 287 150 299 184
rect 333 150 345 184
rect 287 116 345 150
rect 287 82 299 116
rect 333 82 345 116
rect 287 48 345 82
rect 287 14 299 48
rect 333 14 345 48
rect 287 -20 345 14
rect 287 -54 299 -20
rect 333 -54 345 -20
rect 287 -88 345 -54
rect 287 -122 299 -88
rect 333 -122 345 -88
rect 287 -156 345 -122
rect 287 -190 299 -156
rect 333 -190 345 -156
rect 287 -224 345 -190
rect 287 -258 299 -224
rect 333 -258 345 -224
rect 287 -292 345 -258
rect 287 -326 299 -292
rect 333 -326 345 -292
rect 287 -444 345 -326
<< mvndiffc >>
rect -333 354 -299 388
rect -333 286 -299 320
rect -333 218 -299 252
rect -333 150 -299 184
rect -333 82 -299 116
rect -333 14 -299 48
rect -333 -54 -299 -20
rect -333 -122 -299 -88
rect -333 -190 -299 -156
rect -333 -258 -299 -224
rect -333 -326 -299 -292
rect -175 354 -141 388
rect -175 286 -141 320
rect -175 218 -141 252
rect -175 150 -141 184
rect -175 82 -141 116
rect -175 14 -141 48
rect -175 -54 -141 -20
rect -175 -122 -141 -88
rect -175 -190 -141 -156
rect -175 -258 -141 -224
rect -175 -326 -141 -292
rect -17 354 17 388
rect -17 286 17 320
rect -17 218 17 252
rect -17 150 17 184
rect -17 82 17 116
rect -17 14 17 48
rect -17 -54 17 -20
rect -17 -122 17 -88
rect -17 -190 17 -156
rect -17 -258 17 -224
rect -17 -326 17 -292
rect 141 354 175 388
rect 141 286 175 320
rect 141 218 175 252
rect 141 150 175 184
rect 141 82 175 116
rect 141 14 175 48
rect 141 -54 175 -20
rect 141 -122 175 -88
rect 141 -190 175 -156
rect 141 -258 175 -224
rect 141 -326 175 -292
rect 299 354 333 388
rect 299 286 333 320
rect 299 218 333 252
rect 299 150 333 184
rect 299 82 333 116
rect 299 14 333 48
rect 299 -54 333 -20
rect 299 -122 333 -88
rect 299 -190 333 -156
rect 299 -258 333 -224
rect 299 -326 333 -292
<< poly >>
rect -287 506 -187 532
rect -129 506 -29 532
rect 29 506 129 532
rect 187 506 287 532
rect -287 -482 -187 -444
rect -287 -516 -254 -482
rect -220 -516 -187 -482
rect -287 -532 -187 -516
rect -129 -482 -29 -444
rect -129 -516 -96 -482
rect -62 -516 -29 -482
rect -129 -532 -29 -516
rect 29 -482 129 -444
rect 29 -516 62 -482
rect 96 -516 129 -482
rect 29 -532 129 -516
rect 187 -482 287 -444
rect 187 -516 220 -482
rect 254 -516 287 -482
rect 187 -532 287 -516
<< polycont >>
rect -254 -516 -220 -482
rect -96 -516 -62 -482
rect 62 -516 96 -482
rect 220 -516 254 -482
<< locali >>
rect -333 480 -299 494
rect -333 408 -299 446
rect -17 480 17 494
rect -333 336 -299 354
rect -333 264 -299 286
rect -333 192 -299 218
rect -333 120 -299 150
rect -333 48 -299 82
rect -333 -20 -299 14
rect -333 -88 -299 -58
rect -333 -156 -299 -130
rect -333 -224 -299 -202
rect -333 -292 -299 -274
rect -333 -384 -299 -346
rect -175 388 -141 417
rect -175 320 -141 338
rect -175 252 -141 266
rect -175 184 -141 194
rect -175 116 -141 122
rect -175 48 -141 50
rect -175 12 -141 14
rect -175 -60 -141 -54
rect -175 -132 -141 -122
rect -175 -204 -141 -190
rect -175 -276 -141 -258
rect -175 -355 -141 -326
rect -17 408 17 446
rect 299 480 333 494
rect -17 336 17 354
rect -17 264 17 286
rect -17 192 17 218
rect -17 120 17 150
rect -17 48 17 82
rect -17 -20 17 14
rect -17 -88 17 -58
rect -17 -156 17 -130
rect -17 -224 17 -202
rect -17 -292 17 -274
rect -333 -432 -299 -418
rect -17 -384 17 -346
rect 141 388 175 417
rect 141 320 175 338
rect 141 252 175 266
rect 141 184 175 194
rect 141 116 175 122
rect 141 48 175 50
rect 141 12 175 14
rect 141 -60 175 -54
rect 141 -132 175 -122
rect 141 -204 175 -190
rect 141 -276 175 -258
rect 141 -355 175 -326
rect 299 408 333 446
rect 299 336 333 354
rect 299 264 333 286
rect 299 192 333 218
rect 299 120 333 150
rect 299 48 333 82
rect 299 -20 333 14
rect 299 -88 333 -58
rect 299 -156 333 -130
rect 299 -224 333 -202
rect 299 -292 333 -274
rect -17 -432 17 -418
rect 299 -384 333 -346
rect 299 -432 333 -418
rect -287 -516 -254 -482
rect -220 -516 -187 -482
rect -129 -516 -96 -482
rect -62 -516 -29 -482
rect 29 -516 62 -482
rect 96 -516 129 -482
rect 187 -516 220 -482
rect 254 -516 287 -482
<< viali >>
rect -333 446 -299 480
rect -17 446 17 480
rect -333 388 -299 408
rect -333 374 -299 388
rect -333 320 -299 336
rect -333 302 -299 320
rect -333 252 -299 264
rect -333 230 -299 252
rect -333 184 -299 192
rect -333 158 -299 184
rect -333 116 -299 120
rect -333 86 -299 116
rect -333 14 -299 48
rect -333 -54 -299 -24
rect -333 -58 -299 -54
rect -333 -122 -299 -96
rect -333 -130 -299 -122
rect -333 -190 -299 -168
rect -333 -202 -299 -190
rect -333 -258 -299 -240
rect -333 -274 -299 -258
rect -333 -326 -299 -312
rect -333 -346 -299 -326
rect -175 354 -141 372
rect -175 338 -141 354
rect -175 286 -141 300
rect -175 266 -141 286
rect -175 218 -141 228
rect -175 194 -141 218
rect -175 150 -141 156
rect -175 122 -141 150
rect -175 82 -141 84
rect -175 50 -141 82
rect -175 -20 -141 12
rect -175 -22 -141 -20
rect -175 -88 -141 -60
rect -175 -94 -141 -88
rect -175 -156 -141 -132
rect -175 -166 -141 -156
rect -175 -224 -141 -204
rect -175 -238 -141 -224
rect -175 -292 -141 -276
rect -175 -310 -141 -292
rect 299 446 333 480
rect -17 388 17 408
rect -17 374 17 388
rect -17 320 17 336
rect -17 302 17 320
rect -17 252 17 264
rect -17 230 17 252
rect -17 184 17 192
rect -17 158 17 184
rect -17 116 17 120
rect -17 86 17 116
rect -17 14 17 48
rect -17 -54 17 -24
rect -17 -58 17 -54
rect -17 -122 17 -96
rect -17 -130 17 -122
rect -17 -190 17 -168
rect -17 -202 17 -190
rect -17 -258 17 -240
rect -17 -274 17 -258
rect -17 -326 17 -312
rect -17 -346 17 -326
rect -333 -418 -299 -384
rect 141 354 175 372
rect 141 338 175 354
rect 141 286 175 300
rect 141 266 175 286
rect 141 218 175 228
rect 141 194 175 218
rect 141 150 175 156
rect 141 122 175 150
rect 141 82 175 84
rect 141 50 175 82
rect 141 -20 175 12
rect 141 -22 175 -20
rect 141 -88 175 -60
rect 141 -94 175 -88
rect 141 -156 175 -132
rect 141 -166 175 -156
rect 141 -224 175 -204
rect 141 -238 175 -224
rect 141 -292 175 -276
rect 141 -310 175 -292
rect 299 388 333 408
rect 299 374 333 388
rect 299 320 333 336
rect 299 302 333 320
rect 299 252 333 264
rect 299 230 333 252
rect 299 184 333 192
rect 299 158 333 184
rect 299 116 333 120
rect 299 86 333 116
rect 299 14 333 48
rect 299 -54 333 -24
rect 299 -58 333 -54
rect 299 -122 333 -96
rect 299 -130 333 -122
rect 299 -190 333 -168
rect 299 -202 333 -190
rect 299 -258 333 -240
rect 299 -274 333 -258
rect 299 -326 333 -312
rect 299 -346 333 -326
rect -17 -418 17 -384
rect 299 -418 333 -384
rect -254 -516 -220 -482
rect -96 -516 -62 -482
rect 62 -516 96 -482
rect 220 -516 254 -482
<< metal1 >>
rect -339 480 -293 506
rect -339 446 -333 480
rect -299 446 -293 480
rect -339 408 -293 446
rect -23 480 23 506
rect -23 446 -17 480
rect 17 446 23 480
rect -339 374 -333 408
rect -299 374 -293 408
rect -339 336 -293 374
rect -339 302 -333 336
rect -299 302 -293 336
rect -339 264 -293 302
rect -339 230 -333 264
rect -299 230 -293 264
rect -339 192 -293 230
rect -339 158 -333 192
rect -299 158 -293 192
rect -339 120 -293 158
rect -339 86 -333 120
rect -299 86 -293 120
rect -339 48 -293 86
rect -339 14 -333 48
rect -299 14 -293 48
rect -339 -24 -293 14
rect -339 -58 -333 -24
rect -299 -58 -293 -24
rect -339 -96 -293 -58
rect -339 -130 -333 -96
rect -299 -130 -293 -96
rect -339 -168 -293 -130
rect -339 -202 -333 -168
rect -299 -202 -293 -168
rect -339 -240 -293 -202
rect -339 -274 -333 -240
rect -299 -274 -293 -240
rect -339 -312 -293 -274
rect -339 -346 -333 -312
rect -299 -346 -293 -312
rect -339 -384 -293 -346
rect -181 372 -135 413
rect -181 338 -175 372
rect -141 338 -135 372
rect -181 300 -135 338
rect -181 266 -175 300
rect -141 266 -135 300
rect -181 228 -135 266
rect -181 194 -175 228
rect -141 194 -135 228
rect -181 156 -135 194
rect -181 122 -175 156
rect -141 122 -135 156
rect -181 84 -135 122
rect -181 50 -175 84
rect -141 50 -135 84
rect -181 12 -135 50
rect -181 -22 -175 12
rect -141 -22 -135 12
rect -181 -60 -135 -22
rect -181 -94 -175 -60
rect -141 -94 -135 -60
rect -181 -132 -135 -94
rect -181 -166 -175 -132
rect -141 -166 -135 -132
rect -181 -204 -135 -166
rect -181 -238 -175 -204
rect -141 -238 -135 -204
rect -181 -276 -135 -238
rect -181 -310 -175 -276
rect -141 -310 -135 -276
rect -181 -351 -135 -310
rect -23 408 23 446
rect 293 480 339 506
rect 293 446 299 480
rect 333 446 339 480
rect -23 374 -17 408
rect 17 374 23 408
rect -23 336 23 374
rect -23 302 -17 336
rect 17 302 23 336
rect -23 264 23 302
rect -23 230 -17 264
rect 17 230 23 264
rect -23 192 23 230
rect -23 158 -17 192
rect 17 158 23 192
rect -23 120 23 158
rect -23 86 -17 120
rect 17 86 23 120
rect -23 48 23 86
rect -23 14 -17 48
rect 17 14 23 48
rect -23 -24 23 14
rect -23 -58 -17 -24
rect 17 -58 23 -24
rect -23 -96 23 -58
rect -23 -130 -17 -96
rect 17 -130 23 -96
rect -23 -168 23 -130
rect -23 -202 -17 -168
rect 17 -202 23 -168
rect -23 -240 23 -202
rect -23 -274 -17 -240
rect 17 -274 23 -240
rect -23 -312 23 -274
rect -23 -346 -17 -312
rect 17 -346 23 -312
rect -339 -418 -333 -384
rect -299 -418 -293 -384
rect -339 -444 -293 -418
rect -23 -384 23 -346
rect 135 372 181 413
rect 135 338 141 372
rect 175 338 181 372
rect 135 300 181 338
rect 135 266 141 300
rect 175 266 181 300
rect 135 228 181 266
rect 135 194 141 228
rect 175 194 181 228
rect 135 156 181 194
rect 135 122 141 156
rect 175 122 181 156
rect 135 84 181 122
rect 135 50 141 84
rect 175 50 181 84
rect 135 12 181 50
rect 135 -22 141 12
rect 175 -22 181 12
rect 135 -60 181 -22
rect 135 -94 141 -60
rect 175 -94 181 -60
rect 135 -132 181 -94
rect 135 -166 141 -132
rect 175 -166 181 -132
rect 135 -204 181 -166
rect 135 -238 141 -204
rect 175 -238 181 -204
rect 135 -276 181 -238
rect 135 -310 141 -276
rect 175 -310 181 -276
rect 135 -351 181 -310
rect 293 408 339 446
rect 293 374 299 408
rect 333 374 339 408
rect 293 336 339 374
rect 293 302 299 336
rect 333 302 339 336
rect 293 264 339 302
rect 293 230 299 264
rect 333 230 339 264
rect 293 192 339 230
rect 293 158 299 192
rect 333 158 339 192
rect 293 120 339 158
rect 293 86 299 120
rect 333 86 339 120
rect 293 48 339 86
rect 293 14 299 48
rect 333 14 339 48
rect 293 -24 339 14
rect 293 -58 299 -24
rect 333 -58 339 -24
rect 293 -96 339 -58
rect 293 -130 299 -96
rect 333 -130 339 -96
rect 293 -168 339 -130
rect 293 -202 299 -168
rect 333 -202 339 -168
rect 293 -240 339 -202
rect 293 -274 299 -240
rect 333 -274 339 -240
rect 293 -312 339 -274
rect 293 -346 299 -312
rect 333 -346 339 -312
rect -23 -418 -17 -384
rect 17 -418 23 -384
rect -23 -444 23 -418
rect 293 -384 339 -346
rect 293 -418 299 -384
rect 333 -418 339 -384
rect 293 -444 339 -418
rect -283 -482 -191 -476
rect -283 -516 -254 -482
rect -220 -516 -191 -482
rect -283 -522 -191 -516
rect -125 -482 -33 -476
rect -125 -516 -96 -482
rect -62 -516 -33 -482
rect -125 -522 -33 -516
rect 33 -482 125 -476
rect 33 -516 62 -482
rect 96 -516 125 -482
rect 33 -522 125 -516
rect 191 -482 283 -476
rect 191 -516 220 -482
rect 254 -516 283 -482
rect 191 -522 283 -516
<< end >>
