magic
tech sky130A
magscale 1 2
timestamp 1770222546
<< metal3 >>
rect -5492 5172 -120 5200
rect -5492 148 -204 5172
rect -140 148 -120 5172
rect -5492 120 -120 148
rect 120 5172 5492 5200
rect 120 148 5408 5172
rect 5472 148 5492 5172
rect 120 120 5492 148
rect -5492 -148 -120 -120
rect -5492 -5172 -204 -148
rect -140 -5172 -120 -148
rect -5492 -5200 -120 -5172
rect 120 -148 5492 -120
rect 120 -5172 5408 -148
rect 5472 -5172 5492 -148
rect 120 -5200 5492 -5172
<< via3 >>
rect -204 148 -140 5172
rect 5408 148 5472 5172
rect -204 -5172 -140 -148
rect 5408 -5172 5472 -148
<< mimcap >>
rect -5452 5120 -452 5160
rect -5452 200 -5412 5120
rect -492 200 -452 5120
rect -5452 160 -452 200
rect 160 5120 5160 5160
rect 160 200 200 5120
rect 5120 200 5160 5120
rect 160 160 5160 200
rect -5452 -200 -452 -160
rect -5452 -5120 -5412 -200
rect -492 -5120 -452 -200
rect -5452 -5160 -452 -5120
rect 160 -200 5160 -160
rect 160 -5120 200 -200
rect 5120 -5120 5160 -200
rect 160 -5160 5160 -5120
<< mimcapcontact >>
rect -5412 200 -492 5120
rect 200 200 5120 5120
rect -5412 -5120 -492 -200
rect 200 -5120 5120 -200
<< metal4 >>
rect -3004 5121 -2900 5320
rect -224 5172 -120 5320
rect -5413 5120 -491 5121
rect -5413 200 -5412 5120
rect -492 200 -491 5120
rect -5413 199 -491 200
rect -3004 -199 -2900 199
rect -224 148 -204 5172
rect -140 148 -120 5172
rect 2608 5121 2712 5320
rect 5388 5172 5492 5320
rect 199 5120 5121 5121
rect 199 200 200 5120
rect 5120 200 5121 5120
rect 199 199 5121 200
rect -224 -148 -120 148
rect -5413 -200 -491 -199
rect -5413 -5120 -5412 -200
rect -492 -5120 -491 -200
rect -5413 -5121 -491 -5120
rect -3004 -5320 -2900 -5121
rect -224 -5172 -204 -148
rect -140 -5172 -120 -148
rect 2608 -199 2712 199
rect 5388 148 5408 5172
rect 5472 148 5492 5172
rect 5388 -148 5492 148
rect 199 -200 5121 -199
rect 199 -5120 200 -200
rect 5120 -5120 5121 -200
rect 199 -5121 5121 -5120
rect -224 -5320 -120 -5172
rect 2608 -5320 2712 -5121
rect 5388 -5172 5408 -148
rect 5472 -5172 5492 -148
rect 5388 -5320 5492 -5172
<< properties >>
string FIXED_BBOX 120 120 5200 5200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 25.0 val 1.269k carea 2.00 cperi 0.19 class capacitor nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
