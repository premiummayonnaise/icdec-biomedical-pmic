magic
tech sky130A
magscale 1 2
timestamp 1769402310
<< error_p >>
rect -34 381 34 387
rect -34 347 -22 381
rect -34 341 34 347
<< nmos >>
rect -125 -371 125 309
<< ndiff >>
rect -183 297 -125 309
rect -183 -359 -171 297
rect -137 -359 -125 297
rect -183 -371 -125 -359
rect 125 297 183 309
rect 125 -359 137 297
rect 171 -359 183 297
rect 125 -371 183 -359
<< ndiffc >>
rect -171 -359 -137 297
rect 137 -359 171 297
<< poly >>
rect -38 381 38 397
rect -38 364 -22 381
rect -125 347 -22 364
rect 22 364 38 381
rect 22 347 125 364
rect -125 309 125 347
rect -125 -397 125 -371
<< polycont >>
rect -22 347 22 381
<< locali >>
rect -38 347 -22 381
rect 22 347 38 381
rect -171 297 -137 313
rect -171 -375 -137 -359
rect 137 297 171 313
rect 137 -375 171 -359
<< viali >>
rect -22 347 22 381
rect -171 -359 -137 297
rect 137 -359 171 297
<< metal1 >>
rect -34 381 34 387
rect -34 347 -22 381
rect 22 347 34 381
rect -34 341 34 347
rect -177 297 -131 309
rect -177 -359 -171 297
rect -137 -359 -131 297
rect -177 -371 -131 -359
rect 131 297 177 309
rect 131 -359 137 297
rect 171 -359 177 297
rect 131 -371 177 -359
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.4 l 1.25 m 1 nf 1 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
