magic
tech sky130A
magscale 1 2
timestamp 1769616064
<< error_p >>
rect -521 254 -463 260
rect -193 254 -135 260
rect 135 254 193 260
rect 463 254 521 260
rect -521 220 -509 254
rect -193 220 -181 254
rect 135 220 147 254
rect 463 220 475 254
rect -521 214 -463 220
rect -193 214 -135 220
rect 135 214 193 220
rect 463 214 521 220
<< pwell >>
rect -795 -440 795 440
<< mvnmos >>
rect -567 -244 -417 182
rect -239 -244 -89 182
rect 89 -244 239 182
rect 417 -244 567 182
<< mvndiff >>
rect -625 170 -567 182
rect -625 -232 -613 170
rect -579 -232 -567 170
rect -625 -244 -567 -232
rect -417 170 -359 182
rect -417 -232 -405 170
rect -371 -232 -359 170
rect -417 -244 -359 -232
rect -297 170 -239 182
rect -297 -232 -285 170
rect -251 -232 -239 170
rect -297 -244 -239 -232
rect -89 170 -31 182
rect -89 -232 -77 170
rect -43 -232 -31 170
rect -89 -244 -31 -232
rect 31 170 89 182
rect 31 -232 43 170
rect 77 -232 89 170
rect 31 -244 89 -232
rect 239 170 297 182
rect 239 -232 251 170
rect 285 -232 297 170
rect 239 -244 297 -232
rect 359 170 417 182
rect 359 -232 371 170
rect 405 -232 417 170
rect 359 -244 417 -232
rect 567 170 625 182
rect 567 -232 579 170
rect 613 -232 625 170
rect 567 -244 625 -232
<< mvndiffc >>
rect -613 -232 -579 170
rect -405 -232 -371 170
rect -285 -232 -251 170
rect -77 -232 -43 170
rect 43 -232 77 170
rect 251 -232 285 170
rect 371 -232 405 170
rect 579 -232 613 170
<< mvpsubdiff >>
rect -759 346 759 404
rect -759 296 -701 346
rect -759 -296 -747 296
rect -713 -296 -701 296
rect 701 296 759 346
rect -759 -346 -701 -296
rect 701 -296 713 296
rect 747 -296 759 296
rect 701 -346 759 -296
rect -759 -404 759 -346
<< mvpsubdiffcont >>
rect -747 -296 -713 296
rect 713 -296 747 296
<< poly >>
rect -525 254 -459 270
rect -525 237 -509 254
rect -567 220 -509 237
rect -475 237 -459 254
rect -197 254 -131 270
rect -197 237 -181 254
rect -475 220 -417 237
rect -567 182 -417 220
rect -239 220 -181 237
rect -147 237 -131 254
rect 131 254 197 270
rect 131 237 147 254
rect -147 220 -89 237
rect -239 182 -89 220
rect 89 220 147 237
rect 181 237 197 254
rect 459 254 525 270
rect 459 237 475 254
rect 181 220 239 237
rect 89 182 239 220
rect 417 220 475 237
rect 509 237 525 254
rect 509 220 567 237
rect 417 182 567 220
rect -567 -270 -417 -244
rect -239 -270 -89 -244
rect 89 -270 239 -244
rect 417 -270 567 -244
<< polycont >>
rect -509 220 -475 254
rect -181 220 -147 254
rect 147 220 181 254
rect 475 220 509 254
<< locali >>
rect -747 296 -713 312
rect 713 296 747 312
rect -525 220 -509 254
rect -475 220 -459 254
rect -197 220 -181 254
rect -147 220 -131 254
rect 131 220 147 254
rect 181 220 197 254
rect 459 220 475 254
rect 509 220 525 254
rect -613 170 -579 186
rect -613 -248 -579 -232
rect -405 170 -371 186
rect -405 -248 -371 -232
rect -285 170 -251 186
rect -285 -248 -251 -232
rect -77 170 -43 186
rect -77 -248 -43 -232
rect 43 170 77 186
rect 43 -248 77 -232
rect 251 170 285 186
rect 251 -248 285 -232
rect 371 170 405 186
rect 371 -248 405 -232
rect 579 170 613 186
rect 579 -248 613 -232
rect -747 -312 -713 -296
rect 713 -312 747 -296
<< viali >>
rect -509 220 -475 254
rect -181 220 -147 254
rect 147 220 181 254
rect 475 220 509 254
rect -613 -232 -579 170
rect -405 -232 -371 170
rect -285 -232 -251 170
rect -77 -232 -43 170
rect 43 -232 77 170
rect 251 -232 285 170
rect 371 -232 405 170
rect 579 -232 613 170
<< metal1 >>
rect -521 254 -463 260
rect -521 220 -509 254
rect -475 220 -463 254
rect -521 214 -463 220
rect -193 254 -135 260
rect -193 220 -181 254
rect -147 220 -135 254
rect -193 214 -135 220
rect 135 254 193 260
rect 135 220 147 254
rect 181 220 193 254
rect 135 214 193 220
rect 463 254 521 260
rect 463 220 475 254
rect 509 220 521 254
rect 463 214 521 220
rect -619 170 -573 182
rect -619 -232 -613 170
rect -579 -232 -573 170
rect -619 -244 -573 -232
rect -411 170 -365 182
rect -411 -232 -405 170
rect -371 -232 -365 170
rect -411 -244 -365 -232
rect -291 170 -245 182
rect -291 -232 -285 170
rect -251 -232 -245 170
rect -291 -244 -245 -232
rect -83 170 -37 182
rect -83 -232 -77 170
rect -43 -232 -37 170
rect -83 -244 -37 -232
rect 37 170 83 182
rect 37 -232 43 170
rect 77 -232 83 170
rect 37 -244 83 -232
rect 245 170 291 182
rect 245 -232 251 170
rect 285 -232 291 170
rect 245 -244 291 -232
rect 365 170 411 182
rect 365 -232 371 170
rect 405 -232 411 170
rect 365 -244 411 -232
rect 573 170 619 182
rect 573 -232 579 170
rect 613 -232 619 170
rect 573 -244 619 -232
<< properties >>
string FIXED_BBOX -730 -375 730 375
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.125 l 0.75 m 1 nf 4 diffcov 100 polycov 20 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
