magic
tech sky130A
magscale 1 2
timestamp 1769397192
<< pwell >>
rect -783 -460 783 460
<< nmos >>
rect -587 -250 -337 250
rect -279 -250 -29 250
rect 29 -250 279 250
rect 337 -250 587 250
<< ndiff >>
rect -645 238 -587 250
rect -645 -238 -633 238
rect -599 -238 -587 238
rect -645 -250 -587 -238
rect -337 238 -279 250
rect -337 -238 -325 238
rect -291 -238 -279 238
rect -337 -250 -279 -238
rect -29 238 29 250
rect -29 -238 -17 238
rect 17 -238 29 238
rect -29 -250 29 -238
rect 279 238 337 250
rect 279 -238 291 238
rect 325 -238 337 238
rect 279 -250 337 -238
rect 587 238 645 250
rect 587 -238 599 238
rect 633 -238 645 238
rect 587 -250 645 -238
<< ndiffc >>
rect -633 -238 -599 238
rect -325 -238 -291 238
rect -17 -238 17 238
rect 291 -238 325 238
rect 599 -238 633 238
<< psubdiff >>
rect -747 390 -651 424
rect 651 390 747 424
rect -747 328 -713 390
rect 713 328 747 390
rect -747 -390 -713 -328
rect 713 -390 747 -328
rect -747 -424 -651 -390
rect 651 -424 747 -390
<< psubdiffcont >>
rect -651 390 651 424
rect -747 -328 -713 328
rect 713 -328 747 328
rect -651 -424 651 -390
<< poly >>
rect -587 322 -337 338
rect -587 288 -571 322
rect -353 288 -337 322
rect -587 250 -337 288
rect -279 322 -29 338
rect -279 288 -263 322
rect -45 288 -29 322
rect -279 250 -29 288
rect 29 322 279 338
rect 29 288 45 322
rect 263 288 279 322
rect 29 250 279 288
rect 337 322 587 338
rect 337 288 353 322
rect 571 288 587 322
rect 337 250 587 288
rect -587 -288 -337 -250
rect -587 -322 -571 -288
rect -353 -322 -337 -288
rect -587 -338 -337 -322
rect -279 -288 -29 -250
rect -279 -322 -263 -288
rect -45 -322 -29 -288
rect -279 -338 -29 -322
rect 29 -288 279 -250
rect 29 -322 45 -288
rect 263 -322 279 -288
rect 29 -338 279 -322
rect 337 -288 587 -250
rect 337 -322 353 -288
rect 571 -322 587 -288
rect 337 -338 587 -322
<< polycont >>
rect -571 288 -353 322
rect -263 288 -45 322
rect 45 288 263 322
rect 353 288 571 322
rect -571 -322 -353 -288
rect -263 -322 -45 -288
rect 45 -322 263 -288
rect 353 -322 571 -288
<< locali >>
rect -747 390 -651 424
rect 651 390 747 424
rect -747 328 -713 390
rect 713 328 747 390
rect -587 288 -571 322
rect -353 288 -337 322
rect -279 288 -263 322
rect -45 288 -29 322
rect 29 288 45 322
rect 263 288 279 322
rect 337 288 353 322
rect 571 288 587 322
rect -633 238 -599 254
rect -633 -254 -599 -238
rect -325 238 -291 254
rect -325 -254 -291 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 291 238 325 254
rect 291 -254 325 -238
rect 599 238 633 254
rect 599 -254 633 -238
rect -587 -322 -571 -288
rect -353 -322 -337 -288
rect -279 -322 -263 -288
rect -45 -322 -29 -288
rect 29 -322 45 -288
rect 263 -322 279 -288
rect 337 -322 353 -288
rect 571 -322 587 -288
rect -747 -390 -713 -328
rect 713 -390 747 -328
rect -747 -424 -651 -390
rect 651 -424 747 -390
<< viali >>
rect -571 288 -353 322
rect -263 288 -45 322
rect 45 288 263 322
rect 353 288 571 322
rect -633 -238 -599 238
rect -325 -238 -291 238
rect -17 -238 17 238
rect 291 -238 325 238
rect 599 -238 633 238
rect -571 -322 -353 -288
rect -263 -322 -45 -288
rect 45 -322 263 -288
rect 353 -322 571 -288
<< metal1 >>
rect -583 322 -341 328
rect -583 288 -571 322
rect -353 288 -341 322
rect -583 282 -341 288
rect -275 322 -33 328
rect -275 288 -263 322
rect -45 288 -33 322
rect -275 282 -33 288
rect 33 322 275 328
rect 33 288 45 322
rect 263 288 275 322
rect 33 282 275 288
rect 341 322 583 328
rect 341 288 353 322
rect 571 288 583 322
rect 341 282 583 288
rect -639 238 -593 250
rect -639 -238 -633 238
rect -599 -238 -593 238
rect -639 -250 -593 -238
rect -331 238 -285 250
rect -331 -238 -325 238
rect -291 -238 -285 238
rect -331 -250 -285 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 285 238 331 250
rect 285 -238 291 238
rect 325 -238 331 238
rect 285 -250 331 -238
rect 593 238 639 250
rect 593 -238 599 238
rect 633 -238 639 238
rect 593 -250 639 -238
rect -583 -288 -341 -282
rect -583 -322 -571 -288
rect -353 -322 -341 -288
rect -583 -328 -341 -322
rect -275 -288 -33 -282
rect -275 -322 -263 -288
rect -45 -322 -33 -288
rect -275 -328 -33 -322
rect 33 -288 275 -282
rect 33 -322 45 -288
rect 263 -322 275 -288
rect 33 -328 275 -322
rect 341 -288 583 -282
rect 341 -322 353 -288
rect 571 -322 583 -288
rect 341 -328 583 -322
<< properties >>
string FIXED_BBOX -730 -407 730 407
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
