magic
tech sky130A
magscale 1 2
timestamp 1769076474
<< mvnmos >>
rect -50 -385 50 447
<< mvndiff >>
rect -108 435 -50 447
rect -108 -373 -96 435
rect -62 -373 -50 435
rect -108 -385 -50 -373
rect 50 435 108 447
rect 50 -373 62 435
rect 96 -373 108 435
rect 50 -385 108 -373
<< mvndiffc >>
rect -96 -373 -62 435
rect 62 -373 96 435
<< poly >>
rect -50 447 50 473
rect -50 -423 50 -385
rect -50 -457 -34 -423
rect 34 -457 50 -423
rect -50 -473 50 -457
<< polycont >>
rect -34 -457 34 -423
<< locali >>
rect -96 435 -62 451
rect -96 -389 -62 -373
rect 62 435 96 451
rect 62 -389 96 -373
rect -50 -457 -34 -423
rect 34 -457 50 -423
<< viali >>
rect -96 -373 -62 435
rect 62 -373 96 435
rect -34 -457 34 -423
<< metal1 >>
rect -102 435 -56 447
rect -102 -373 -96 435
rect -62 -373 -56 435
rect -102 -385 -56 -373
rect 56 435 102 447
rect 56 -373 62 435
rect 96 -373 102 435
rect 56 -385 102 -373
rect -46 -423 46 -417
rect -46 -457 -34 -423
rect 34 -457 46 -423
rect -46 -463 46 -457
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.16 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
