magic
tech sky130A
magscale 1 2
timestamp 1769959185
<< pwell >>
rect 800 900 11500 6000
<< psubdiff >>
rect 800 5980 11500 6000
rect 800 5820 1020 5980
rect 11280 5820 11500 5980
rect 800 5800 11500 5820
rect 800 5780 1000 5800
rect 800 1120 820 5780
rect 980 1120 1000 5780
rect 11300 5760 11500 5800
rect 1200 5500 3500 5600
rect 1200 3700 1300 5500
rect 3400 5480 3500 5500
rect 3400 3720 3420 5480
rect 3480 3720 3500 5480
rect 3400 3700 3500 3720
rect 1200 3600 3500 3700
rect 3600 5500 5900 5600
rect 3600 5480 3700 5500
rect 3600 3720 3620 5480
rect 3680 3720 3700 5480
rect 3600 3700 3700 3720
rect 5800 3700 5900 5500
rect 3600 3600 5900 3700
rect 6400 5500 8700 5600
rect 6400 3700 6500 5500
rect 8600 5480 8700 5500
rect 8600 3720 8620 5480
rect 8680 3720 8700 5480
rect 8600 3700 8700 3720
rect 6400 3600 8700 3700
rect 8800 5500 11100 5600
rect 8800 5480 8900 5500
rect 8800 3720 8820 5480
rect 8880 3720 8900 5480
rect 8800 3700 8900 3720
rect 11000 3700 11100 5500
rect 8800 3600 11100 3700
rect 1200 3200 3500 3300
rect 1200 1400 1300 3200
rect 3400 3180 3500 3200
rect 3400 1420 3420 3180
rect 3480 1420 3500 3180
rect 3400 1400 3500 1420
rect 1200 1300 3500 1400
rect 3600 3200 5900 3300
rect 3600 3180 3700 3200
rect 3600 1420 3620 3180
rect 3680 1420 3700 3180
rect 3600 1400 3700 1420
rect 5800 1400 5900 3200
rect 3600 1300 5900 1400
rect 6400 3200 8700 3300
rect 6400 1400 6500 3200
rect 8600 3180 8700 3200
rect 8600 1420 8620 3180
rect 8680 1420 8700 3180
rect 8600 1400 8700 1420
rect 6400 1300 8700 1400
rect 8800 3200 11100 3300
rect 8800 3180 8900 3200
rect 8800 1420 8820 3180
rect 8880 1420 8900 3180
rect 8800 1400 8900 1420
rect 11000 1400 11100 3200
rect 8800 1300 11100 1400
rect 800 1100 1000 1120
rect 11300 1100 11320 5760
rect 11480 1100 11500 5760
rect 800 1080 11500 1100
rect 800 920 1020 1080
rect 11280 920 11500 1080
rect 800 900 11500 920
<< psubdiffcont >>
rect 1020 5820 11280 5980
rect 820 1120 980 5780
rect 3420 3720 3480 5480
rect 3620 3720 3680 5480
rect 8620 3720 8680 5480
rect 8820 3720 8880 5480
rect 3420 1420 3480 3180
rect 3620 1420 3680 3180
rect 8620 1420 8680 3180
rect 8820 1420 8880 3180
rect 11320 1100 11480 5760
rect 1020 920 11280 1080
<< locali >>
rect 800 5980 11500 6000
rect 800 5820 1020 5980
rect 11280 5820 11500 5980
rect 800 5780 11500 5820
rect 800 1120 820 5780
rect 980 5760 11500 5780
rect 980 5600 11320 5760
rect 980 1300 1200 5600
rect 1440 3600 1720 5420
rect 1960 3900 2120 5600
rect 2240 3840 2460 5380
rect 2580 3900 2740 5600
rect 3500 5500 3600 5600
rect 3400 5480 3700 5500
rect 1780 3600 2940 3840
rect 2980 3600 3260 5400
rect 3400 3720 3420 5480
rect 3480 3720 3620 5480
rect 3680 3720 3700 5480
rect 3840 3840 4120 5420
rect 4360 3900 4520 5600
rect 4980 3900 5140 5600
rect 3400 3700 3700 3720
rect 4180 3600 5340 3840
rect 5380 3820 5660 5400
rect 5900 3600 6400 5400
rect 6640 3820 6920 5400
rect 7160 3900 7320 5600
rect 7780 3900 7940 5600
rect 8700 5500 8800 5600
rect 8600 5480 8900 5500
rect 6980 3600 8140 3840
rect 8180 3820 8460 5400
rect 8600 3720 8620 5480
rect 8680 3720 8820 5480
rect 8880 3720 8900 5480
rect 8600 3700 8900 3720
rect 9040 3600 9320 5400
rect 9560 3900 9720 5600
rect 9840 3840 10060 5380
rect 10180 3900 10340 5600
rect 9360 3600 10520 3840
rect 10580 3600 10860 5400
rect 1400 3300 10900 3600
rect 1780 3080 2940 3300
rect 3400 3180 3700 3200
rect 1440 1500 1720 3080
rect 1960 1300 2120 3020
rect 2580 1300 2740 3020
rect 2980 1500 3260 3080
rect 3400 1420 3420 3180
rect 3480 1420 3620 3180
rect 3680 1420 3700 3180
rect 3840 1500 4120 3300
rect 4180 3080 5340 3300
rect 3400 1400 3700 1420
rect 3500 1300 3600 1400
rect 4360 1300 4520 3020
rect 4640 1500 4860 3080
rect 4980 1300 5140 3020
rect 5380 1500 5660 3300
rect 5900 2200 6400 3300
rect 5900 2060 5920 2200
rect 6060 2060 6240 2200
rect 6380 2060 6400 2200
rect 5900 2020 6400 2060
rect 5900 1880 5920 2020
rect 6060 1880 6240 2020
rect 6380 1880 6400 2020
rect 5900 1840 6400 1880
rect 5900 1700 5920 1840
rect 6060 1700 6240 1840
rect 6380 1700 6400 1840
rect 5900 1660 6400 1700
rect 5900 1520 5920 1660
rect 6060 1520 6240 1660
rect 6380 1520 6400 1660
rect 5900 1500 6400 1520
rect 6640 1500 6920 3300
rect 6980 3080 8140 3300
rect 7160 1300 7320 3020
rect 7440 1500 7660 3080
rect 7780 1300 7940 3020
rect 8180 1500 8460 3300
rect 8600 3180 8900 3200
rect 8600 1420 8620 3180
rect 8680 1420 8820 3180
rect 8880 1420 8900 3180
rect 9360 3080 10520 3300
rect 9040 1500 9320 3080
rect 8600 1400 8900 1420
rect 8700 1300 8800 1400
rect 9560 1300 9720 3020
rect 10180 1300 10340 3020
rect 10580 1500 10860 3080
rect 11100 1300 11320 5600
rect 980 1120 11320 1300
rect 800 1100 11320 1120
rect 11480 1100 11500 5760
rect 800 1080 11500 1100
rect 800 920 820 1080
rect 980 920 1020 1080
rect 11280 920 11500 1080
rect 800 900 11500 920
<< viali >>
rect 5920 2060 6060 2200
rect 6240 2060 6380 2200
rect 5920 1880 6060 2020
rect 6240 1880 6380 2020
rect 5920 1700 6060 1840
rect 6240 1700 6380 1840
rect 5920 1520 6060 1660
rect 6240 1520 6380 1660
rect 820 920 980 1080
<< metal1 >>
rect 5800 6380 6480 6400
rect 5800 6320 5820 6380
rect 5880 6320 5900 6380
rect 5960 6320 5980 6380
rect 6040 6320 6060 6380
rect 6120 6320 6160 6380
rect 6220 6320 6240 6380
rect 6300 6320 6320 6380
rect 6380 6320 6400 6380
rect 6460 6320 6480 6380
rect 5800 6260 6480 6320
rect 5800 6200 5820 6260
rect 5880 6200 5900 6260
rect 5960 6200 5980 6260
rect 6040 6200 6060 6260
rect 6120 6200 6160 6260
rect 6220 6200 6240 6260
rect 6300 6200 6320 6260
rect 6380 6200 6400 6260
rect 6460 6200 6480 6260
rect 5800 6180 6480 6200
rect 3800 5260 4160 5300
rect 3800 5200 3820 5260
rect 3880 5200 3900 5260
rect 3960 5200 4000 5260
rect 4060 5200 4080 5260
rect 4140 5200 4160 5260
rect 3800 5180 4160 5200
rect 3800 5120 3820 5180
rect 3880 5120 3900 5180
rect 3960 5120 4000 5180
rect 4060 5120 4080 5180
rect 4140 5120 4160 5180
rect 3800 5100 4160 5120
rect 3800 5040 3820 5100
rect 3880 5040 3900 5100
rect 3960 5040 4000 5100
rect 4060 5040 4080 5100
rect 4140 5040 4160 5100
rect 3800 5020 4160 5040
rect 3800 4960 3820 5020
rect 3880 4960 3900 5020
rect 3960 4960 4000 5020
rect 4060 4960 4080 5020
rect 4140 4960 4160 5020
rect 3800 4940 4160 4960
rect 3800 4880 3820 4940
rect 3880 4880 3900 4940
rect 3960 4880 4000 4940
rect 4060 4880 4080 4940
rect 4140 4880 4160 4940
rect 3800 4860 4160 4880
rect 3800 4800 3820 4860
rect 3880 4800 3900 4860
rect 3960 4800 4000 4860
rect 4060 4800 4080 4860
rect 4140 4800 4160 4860
rect 3800 4780 4160 4800
rect 3800 4720 3820 4780
rect 3880 4720 3900 4780
rect 3960 4720 4000 4780
rect 4060 4720 4080 4780
rect 4140 4720 4160 4780
rect 3800 4700 4160 4720
rect 4660 5260 4840 5300
rect 4720 5200 4780 5260
rect 4660 5180 4840 5200
rect 4720 5120 4780 5180
rect 4660 5100 4840 5120
rect 4720 5040 4780 5100
rect 4660 5020 4840 5040
rect 4720 4960 4780 5020
rect 4660 4940 4840 4960
rect 4720 4880 4780 4940
rect 4660 4860 4840 4880
rect 4720 4800 4780 4860
rect 4660 4780 4840 4800
rect 4720 4720 4780 4780
rect 4660 4700 4840 4720
rect 5340 5260 5700 5300
rect 5340 5200 5380 5260
rect 5440 5200 5460 5260
rect 5520 5200 5540 5260
rect 5600 5200 5620 5260
rect 5680 5200 5700 5260
rect 5340 5180 5700 5200
rect 5340 5120 5380 5180
rect 5440 5120 5460 5180
rect 5520 5120 5540 5180
rect 5600 5120 5620 5180
rect 5680 5120 5700 5180
rect 5340 5100 5700 5120
rect 5340 5040 5380 5100
rect 5440 5040 5460 5100
rect 5520 5040 5540 5100
rect 5600 5040 5620 5100
rect 5680 5040 5700 5100
rect 5340 5020 5700 5040
rect 5340 4960 5380 5020
rect 5440 4960 5460 5020
rect 5520 4960 5540 5020
rect 5600 4960 5620 5020
rect 5680 4960 5700 5020
rect 5340 4940 5700 4960
rect 5340 4880 5380 4940
rect 5440 4880 5460 4940
rect 5520 4880 5540 4940
rect 5600 4880 5620 4940
rect 5680 4880 5700 4940
rect 5340 4860 5700 4880
rect 5340 4800 5380 4860
rect 5440 4800 5460 4860
rect 5520 4800 5540 4860
rect 5600 4800 5620 4860
rect 5680 4800 5700 4860
rect 5340 4780 5700 4800
rect 5340 4720 5380 4780
rect 5440 4720 5460 4780
rect 5520 4720 5540 4780
rect 5600 4720 5620 4780
rect 5680 4720 5700 4780
rect 5340 4700 5700 4720
rect 5900 3600 6400 5400
rect 6600 5260 6960 5300
rect 6600 5200 6640 5260
rect 6700 5200 6720 5260
rect 6780 5200 6800 5260
rect 6860 5200 6880 5260
rect 6940 5200 6960 5260
rect 6600 5180 6960 5200
rect 6600 5120 6640 5180
rect 6700 5120 6720 5180
rect 6780 5120 6800 5180
rect 6860 5120 6880 5180
rect 6940 5120 6960 5180
rect 6600 5100 6960 5120
rect 6600 5040 6640 5100
rect 6700 5040 6720 5100
rect 6780 5040 6800 5100
rect 6860 5040 6880 5100
rect 6940 5040 6960 5100
rect 6600 5020 6960 5040
rect 6600 4960 6640 5020
rect 6700 4960 6720 5020
rect 6780 4960 6800 5020
rect 6860 4960 6880 5020
rect 6940 4960 6960 5020
rect 6600 4940 6960 4960
rect 6600 4880 6640 4940
rect 6700 4880 6720 4940
rect 6780 4880 6800 4940
rect 6860 4880 6880 4940
rect 6940 4880 6960 4940
rect 6600 4860 6960 4880
rect 6600 4800 6640 4860
rect 6700 4800 6720 4860
rect 6780 4800 6800 4860
rect 6860 4800 6880 4860
rect 6940 4800 6960 4860
rect 6600 4780 6960 4800
rect 6600 4720 6640 4780
rect 6700 4720 6720 4780
rect 6780 4720 6800 4780
rect 6860 4720 6880 4780
rect 6940 4720 6960 4780
rect 6600 4700 6960 4720
rect 7460 5260 7640 5300
rect 7520 5200 7580 5260
rect 7460 5180 7640 5200
rect 7520 5120 7580 5180
rect 7460 5100 7640 5120
rect 7520 5040 7580 5100
rect 7460 5020 7640 5040
rect 7520 4960 7580 5020
rect 7460 4940 7640 4960
rect 7520 4880 7580 4940
rect 7460 4860 7640 4880
rect 7520 4800 7580 4860
rect 7460 4780 7640 4800
rect 7520 4720 7580 4780
rect 7460 4700 7640 4720
rect 8140 5260 8500 5300
rect 8140 5200 8160 5260
rect 8220 5200 8240 5260
rect 8300 5200 8360 5260
rect 8420 5200 8440 5260
rect 8140 5180 8500 5200
rect 8140 5120 8160 5180
rect 8220 5120 8240 5180
rect 8300 5120 8360 5180
rect 8420 5120 8440 5180
rect 8140 5100 8500 5120
rect 8140 5040 8160 5100
rect 8220 5040 8240 5100
rect 8300 5040 8360 5100
rect 8420 5040 8440 5100
rect 8140 5020 8500 5040
rect 8140 4960 8160 5020
rect 8220 4960 8240 5020
rect 8300 4960 8360 5020
rect 8420 4960 8440 5020
rect 8140 4940 8500 4960
rect 8140 4880 8160 4940
rect 8220 4880 8240 4940
rect 8300 4880 8360 4940
rect 8420 4880 8440 4940
rect 8140 4860 8500 4880
rect 8140 4800 8160 4860
rect 8220 4800 8240 4860
rect 8300 4800 8360 4860
rect 8420 4800 8440 4860
rect 8140 4780 8500 4800
rect 8140 4720 8160 4780
rect 8220 4720 8240 4780
rect 8300 4720 8360 4780
rect 8420 4720 8440 4780
rect 8140 4700 8500 4720
rect 1400 3300 10900 3600
rect 5900 2200 6400 3300
rect 1400 1680 1760 2200
rect 1460 1620 1480 1680
rect 1540 1620 1620 1680
rect 1680 1620 1700 1680
rect 1400 1600 1760 1620
rect 2260 2160 2440 2200
rect 2320 2100 2380 2160
rect 2260 2080 2440 2100
rect 2320 2020 2380 2080
rect 2260 2000 2440 2020
rect 2320 1940 2380 2000
rect 2260 1920 2440 1940
rect 2320 1860 2380 1920
rect 2260 1840 2440 1860
rect 2320 1780 2380 1840
rect 2260 1760 2440 1780
rect 2320 1700 2380 1760
rect 2260 1680 2440 1700
rect 2320 1620 2380 1680
rect 2260 1600 2440 1620
rect 2940 1680 3300 2200
rect 2940 1620 2980 1680
rect 3040 1620 3060 1680
rect 3120 1620 3160 1680
rect 3220 1620 3240 1680
rect 2940 1600 3300 1620
rect 5900 2060 5920 2200
rect 6060 2060 6240 2200
rect 6380 2060 6400 2200
rect 5900 2020 6400 2060
rect 5900 1880 5920 2020
rect 6060 1880 6240 2020
rect 6380 1880 6400 2020
rect 5900 1840 6400 1880
rect 5900 1700 5920 1840
rect 6060 1700 6240 1840
rect 6380 1700 6400 1840
rect 5900 1660 6400 1700
rect 5900 1520 5920 1660
rect 6060 1520 6240 1660
rect 6380 1520 6400 1660
rect 9000 1680 9360 2200
rect 9000 1620 9020 1680
rect 9080 1620 9100 1680
rect 9160 1620 9180 1680
rect 9240 1620 9260 1680
rect 9320 1620 9360 1680
rect 9000 1600 9360 1620
rect 9860 2160 10040 2200
rect 9920 2100 9980 2160
rect 9860 2080 10040 2100
rect 9920 2020 9980 2080
rect 9860 2000 10040 2020
rect 9920 1940 9980 2000
rect 9860 1920 10040 1940
rect 9920 1860 9980 1920
rect 9860 1840 10040 1860
rect 9920 1780 9980 1840
rect 9860 1760 10040 1780
rect 9920 1700 9980 1760
rect 9860 1680 10040 1700
rect 9920 1620 9980 1680
rect 9860 1600 10040 1620
rect 10540 1680 10900 2200
rect 10540 1620 10580 1680
rect 10640 1620 10660 1680
rect 10720 1620 10740 1680
rect 10800 1620 10820 1680
rect 10880 1620 10900 1680
rect 10540 1600 10900 1620
rect 800 1080 1000 1100
rect 800 920 820 1080
rect 980 920 1000 1080
rect 800 900 1000 920
rect 5900 260 6400 1520
<< via1 >>
rect 5820 6320 5880 6380
rect 5900 6320 5960 6380
rect 5980 6320 6040 6380
rect 6060 6320 6120 6380
rect 6160 6320 6220 6380
rect 6240 6320 6300 6380
rect 6320 6320 6380 6380
rect 6400 6320 6460 6380
rect 5820 6200 5880 6260
rect 5900 6200 5960 6260
rect 5980 6200 6040 6260
rect 6060 6200 6120 6260
rect 6160 6200 6220 6260
rect 6240 6200 6300 6260
rect 6320 6200 6380 6260
rect 6400 6200 6460 6260
rect 3820 5200 3880 5260
rect 3900 5200 3960 5260
rect 4000 5200 4060 5260
rect 4080 5200 4140 5260
rect 3820 5120 3880 5180
rect 3900 5120 3960 5180
rect 4000 5120 4060 5180
rect 4080 5120 4140 5180
rect 3820 5040 3880 5100
rect 3900 5040 3960 5100
rect 4000 5040 4060 5100
rect 4080 5040 4140 5100
rect 3820 4960 3880 5020
rect 3900 4960 3960 5020
rect 4000 4960 4060 5020
rect 4080 4960 4140 5020
rect 3820 4880 3880 4940
rect 3900 4880 3960 4940
rect 4000 4880 4060 4940
rect 4080 4880 4140 4940
rect 3820 4800 3880 4860
rect 3900 4800 3960 4860
rect 4000 4800 4060 4860
rect 4080 4800 4140 4860
rect 3820 4720 3880 4780
rect 3900 4720 3960 4780
rect 4000 4720 4060 4780
rect 4080 4720 4140 4780
rect 4660 5200 4720 5260
rect 4780 5200 4840 5260
rect 4660 5120 4720 5180
rect 4780 5120 4840 5180
rect 4660 5040 4720 5100
rect 4780 5040 4840 5100
rect 4660 4960 4720 5020
rect 4780 4960 4840 5020
rect 4660 4880 4720 4940
rect 4780 4880 4840 4940
rect 4660 4800 4720 4860
rect 4780 4800 4840 4860
rect 4660 4720 4720 4780
rect 4780 4720 4840 4780
rect 5380 5200 5440 5260
rect 5460 5200 5520 5260
rect 5540 5200 5600 5260
rect 5620 5200 5680 5260
rect 5380 5120 5440 5180
rect 5460 5120 5520 5180
rect 5540 5120 5600 5180
rect 5620 5120 5680 5180
rect 5380 5040 5440 5100
rect 5460 5040 5520 5100
rect 5540 5040 5600 5100
rect 5620 5040 5680 5100
rect 5380 4960 5440 5020
rect 5460 4960 5520 5020
rect 5540 4960 5600 5020
rect 5620 4960 5680 5020
rect 5380 4880 5440 4940
rect 5460 4880 5520 4940
rect 5540 4880 5600 4940
rect 5620 4880 5680 4940
rect 5380 4800 5440 4860
rect 5460 4800 5520 4860
rect 5540 4800 5600 4860
rect 5620 4800 5680 4860
rect 5380 4720 5440 4780
rect 5460 4720 5520 4780
rect 5540 4720 5600 4780
rect 5620 4720 5680 4780
rect 6640 5200 6700 5260
rect 6720 5200 6780 5260
rect 6800 5200 6860 5260
rect 6880 5200 6940 5260
rect 6640 5120 6700 5180
rect 6720 5120 6780 5180
rect 6800 5120 6860 5180
rect 6880 5120 6940 5180
rect 6640 5040 6700 5100
rect 6720 5040 6780 5100
rect 6800 5040 6860 5100
rect 6880 5040 6940 5100
rect 6640 4960 6700 5020
rect 6720 4960 6780 5020
rect 6800 4960 6860 5020
rect 6880 4960 6940 5020
rect 6640 4880 6700 4940
rect 6720 4880 6780 4940
rect 6800 4880 6860 4940
rect 6880 4880 6940 4940
rect 6640 4800 6700 4860
rect 6720 4800 6780 4860
rect 6800 4800 6860 4860
rect 6880 4800 6940 4860
rect 6640 4720 6700 4780
rect 6720 4720 6780 4780
rect 6800 4720 6860 4780
rect 6880 4720 6940 4780
rect 7460 5200 7520 5260
rect 7580 5200 7640 5260
rect 7460 5120 7520 5180
rect 7580 5120 7640 5180
rect 7460 5040 7520 5100
rect 7580 5040 7640 5100
rect 7460 4960 7520 5020
rect 7580 4960 7640 5020
rect 7460 4880 7520 4940
rect 7580 4880 7640 4940
rect 7460 4800 7520 4860
rect 7580 4800 7640 4860
rect 7460 4720 7520 4780
rect 7580 4720 7640 4780
rect 8160 5200 8220 5260
rect 8240 5200 8300 5260
rect 8360 5200 8420 5260
rect 8440 5200 8500 5260
rect 8160 5120 8220 5180
rect 8240 5120 8300 5180
rect 8360 5120 8420 5180
rect 8440 5120 8500 5180
rect 8160 5040 8220 5100
rect 8240 5040 8300 5100
rect 8360 5040 8420 5100
rect 8440 5040 8500 5100
rect 8160 4960 8220 5020
rect 8240 4960 8300 5020
rect 8360 4960 8420 5020
rect 8440 4960 8500 5020
rect 8160 4880 8220 4940
rect 8240 4880 8300 4940
rect 8360 4880 8420 4940
rect 8440 4880 8500 4940
rect 8160 4800 8220 4860
rect 8240 4800 8300 4860
rect 8360 4800 8420 4860
rect 8440 4800 8500 4860
rect 8160 4720 8220 4780
rect 8240 4720 8300 4780
rect 8360 4720 8420 4780
rect 8440 4720 8500 4780
rect 1400 1620 1460 1680
rect 1480 1620 1540 1680
rect 1620 1620 1680 1680
rect 1700 1620 1760 1680
rect 2260 2100 2320 2160
rect 2380 2100 2440 2160
rect 2260 2020 2320 2080
rect 2380 2020 2440 2080
rect 2260 1940 2320 2000
rect 2380 1940 2440 2000
rect 2260 1860 2320 1920
rect 2380 1860 2440 1920
rect 2260 1780 2320 1840
rect 2380 1780 2440 1840
rect 2260 1700 2320 1760
rect 2380 1700 2440 1760
rect 2260 1620 2320 1680
rect 2380 1620 2440 1680
rect 2980 1620 3040 1680
rect 3060 1620 3120 1680
rect 3160 1620 3220 1680
rect 3240 1620 3300 1680
rect 9020 1620 9080 1680
rect 9100 1620 9160 1680
rect 9180 1620 9240 1680
rect 9260 1620 9320 1680
rect 9860 2100 9920 2160
rect 9980 2100 10040 2160
rect 9860 2020 9920 2080
rect 9980 2020 10040 2080
rect 9860 1940 9920 2000
rect 9980 1940 10040 2000
rect 9860 1860 9920 1920
rect 9980 1860 10040 1920
rect 9860 1780 9920 1840
rect 9980 1780 10040 1840
rect 9860 1700 9920 1760
rect 9980 1700 10040 1760
rect 9860 1620 9920 1680
rect 9980 1620 10040 1680
rect 10580 1620 10640 1680
rect 10660 1620 10720 1680
rect 10740 1620 10800 1680
rect 10820 1620 10880 1680
<< metal2 >>
rect 5800 6380 6480 6400
rect 5800 6320 5820 6380
rect 5880 6320 5900 6380
rect 5960 6320 5980 6380
rect 6040 6320 6060 6380
rect 6120 6320 6160 6380
rect 6220 6320 6240 6380
rect 6300 6320 6320 6380
rect 6380 6320 6400 6380
rect 6460 6320 6480 6380
rect 5800 6260 6480 6320
rect 5800 6200 5820 6260
rect 5880 6200 5900 6260
rect 5960 6200 5980 6260
rect 6040 6200 6060 6260
rect 6120 6200 6160 6260
rect 6220 6200 6240 6260
rect 6300 6200 6320 6260
rect 6380 6200 6400 6260
rect 6460 6200 6480 6260
rect 5800 5300 6480 6200
rect 800 5260 11500 5300
rect 800 5200 3820 5260
rect 3880 5200 3900 5260
rect 3960 5200 4000 5260
rect 4060 5200 4080 5260
rect 4140 5200 4660 5260
rect 4720 5200 4780 5260
rect 4840 5200 5380 5260
rect 5440 5200 5460 5260
rect 5520 5200 5540 5260
rect 5600 5200 5620 5260
rect 5680 5200 6640 5260
rect 6700 5200 6720 5260
rect 6780 5200 6800 5260
rect 6860 5200 6880 5260
rect 6940 5200 7460 5260
rect 7520 5200 7580 5260
rect 7640 5200 8160 5260
rect 8220 5200 8240 5260
rect 8300 5200 8360 5260
rect 8420 5200 8440 5260
rect 8500 5200 11500 5260
rect 800 5180 11500 5200
rect 800 5120 3820 5180
rect 3880 5120 3900 5180
rect 3960 5120 4000 5180
rect 4060 5120 4080 5180
rect 4140 5120 4660 5180
rect 4720 5120 4780 5180
rect 4840 5120 5380 5180
rect 5440 5120 5460 5180
rect 5520 5120 5540 5180
rect 5600 5120 5620 5180
rect 5680 5120 6640 5180
rect 6700 5120 6720 5180
rect 6780 5120 6800 5180
rect 6860 5120 6880 5180
rect 6940 5120 7460 5180
rect 7520 5120 7580 5180
rect 7640 5120 8160 5180
rect 8220 5120 8240 5180
rect 8300 5120 8360 5180
rect 8420 5120 8440 5180
rect 8500 5120 11500 5180
rect 800 5100 11500 5120
rect 800 5040 3820 5100
rect 3880 5040 3900 5100
rect 3960 5040 4000 5100
rect 4060 5040 4080 5100
rect 4140 5040 4660 5100
rect 4720 5040 4780 5100
rect 4840 5040 5380 5100
rect 5440 5040 5460 5100
rect 5520 5040 5540 5100
rect 5600 5040 5620 5100
rect 5680 5040 6640 5100
rect 6700 5040 6720 5100
rect 6780 5040 6800 5100
rect 6860 5040 6880 5100
rect 6940 5040 7460 5100
rect 7520 5040 7580 5100
rect 7640 5040 8160 5100
rect 8220 5040 8240 5100
rect 8300 5040 8360 5100
rect 8420 5040 8440 5100
rect 8500 5040 11500 5100
rect 800 5020 11500 5040
rect 800 4960 3820 5020
rect 3880 4960 3900 5020
rect 3960 4960 4000 5020
rect 4060 4960 4080 5020
rect 4140 4960 4660 5020
rect 4720 4960 4780 5020
rect 4840 4960 5380 5020
rect 5440 4960 5460 5020
rect 5520 4960 5540 5020
rect 5600 4960 5620 5020
rect 5680 4960 6640 5020
rect 6700 4960 6720 5020
rect 6780 4960 6800 5020
rect 6860 4960 6880 5020
rect 6940 4960 7460 5020
rect 7520 4960 7580 5020
rect 7640 4960 8160 5020
rect 8220 4960 8240 5020
rect 8300 4960 8360 5020
rect 8420 4960 8440 5020
rect 8500 4960 11500 5020
rect 800 4940 11500 4960
rect 800 4880 3820 4940
rect 3880 4880 3900 4940
rect 3960 4880 4000 4940
rect 4060 4880 4080 4940
rect 4140 4880 4660 4940
rect 4720 4880 4780 4940
rect 4840 4880 5380 4940
rect 5440 4880 5460 4940
rect 5520 4880 5540 4940
rect 5600 4880 5620 4940
rect 5680 4880 6640 4940
rect 6700 4880 6720 4940
rect 6780 4880 6800 4940
rect 6860 4880 6880 4940
rect 6940 4880 7460 4940
rect 7520 4880 7580 4940
rect 7640 4880 8160 4940
rect 8220 4880 8240 4940
rect 8300 4880 8360 4940
rect 8420 4880 8440 4940
rect 8500 4880 11500 4940
rect 800 4860 11500 4880
rect 800 4800 3820 4860
rect 3880 4800 3900 4860
rect 3960 4800 4000 4860
rect 4060 4800 4080 4860
rect 4140 4800 4660 4860
rect 4720 4800 4780 4860
rect 4840 4800 5380 4860
rect 5440 4800 5460 4860
rect 5520 4800 5540 4860
rect 5600 4800 5620 4860
rect 5680 4800 6640 4860
rect 6700 4800 6720 4860
rect 6780 4800 6800 4860
rect 6860 4800 6880 4860
rect 6940 4800 7460 4860
rect 7520 4800 7580 4860
rect 7640 4800 8160 4860
rect 8220 4800 8240 4860
rect 8300 4800 8360 4860
rect 8420 4800 8440 4860
rect 8500 4800 11500 4860
rect 800 4780 11500 4800
rect 800 4720 3820 4780
rect 3880 4720 3900 4780
rect 3960 4720 4000 4780
rect 4060 4720 4080 4780
rect 4140 4720 4660 4780
rect 4720 4720 4780 4780
rect 4840 4720 5380 4780
rect 5440 4720 5460 4780
rect 5520 4720 5540 4780
rect 5600 4720 5620 4780
rect 5680 4720 6640 4780
rect 6700 4720 6720 4780
rect 6780 4720 6800 4780
rect 6860 4720 6880 4780
rect 6940 4720 7460 4780
rect 7520 4720 7580 4780
rect 7640 4720 8160 4780
rect 8220 4720 8240 4780
rect 8300 4720 8360 4780
rect 8420 4720 8440 4780
rect 8500 4720 11500 4780
rect 800 4700 11500 4720
rect 5800 2200 6500 4700
rect 800 2160 11500 2200
rect 800 2100 2260 2160
rect 2320 2100 2380 2160
rect 2440 2100 9860 2160
rect 9920 2100 9980 2160
rect 10040 2100 11500 2160
rect 800 2080 11500 2100
rect 800 2020 2260 2080
rect 2320 2020 2380 2080
rect 2440 2020 9860 2080
rect 9920 2020 9980 2080
rect 10040 2020 11500 2080
rect 800 2000 11500 2020
rect 800 1940 2260 2000
rect 2320 1940 2380 2000
rect 2440 1940 9860 2000
rect 9920 1940 9980 2000
rect 10040 1940 11500 2000
rect 800 1920 11500 1940
rect 800 1860 2260 1920
rect 2320 1860 2380 1920
rect 2440 1860 9860 1920
rect 9920 1860 9980 1920
rect 10040 1860 11500 1920
rect 800 1840 11500 1860
rect 800 1780 2260 1840
rect 2320 1780 2380 1840
rect 2440 1780 9860 1840
rect 9920 1780 9980 1840
rect 10040 1780 11500 1840
rect 800 1760 11500 1780
rect 800 1700 2260 1760
rect 2320 1700 2380 1760
rect 2440 1700 9860 1760
rect 9920 1700 9980 1760
rect 10040 1700 11500 1760
rect 800 1680 11500 1700
rect 800 1620 1400 1680
rect 1460 1620 1480 1680
rect 1540 1620 1620 1680
rect 1680 1620 1700 1680
rect 1760 1620 2260 1680
rect 2320 1620 2380 1680
rect 2440 1620 2980 1680
rect 3040 1620 3060 1680
rect 3120 1620 3160 1680
rect 3220 1620 3240 1680
rect 3300 1620 9020 1680
rect 9080 1620 9100 1680
rect 9160 1620 9180 1680
rect 9240 1620 9260 1680
rect 9320 1620 9860 1680
rect 9920 1620 9980 1680
rect 10040 1620 10580 1680
rect 10640 1620 10660 1680
rect 10720 1620 10740 1680
rect 10800 1620 10820 1680
rect 10880 1620 11500 1680
rect 800 1600 11500 1620
use sky130_fd_pr__nfet_g5v0d10v5_986LJA  sky130_fd_pr__nfet_g5v0d10v5_986LJA_0 /foss/designs/icdec-biomedical-pmic/xschem/error-amplifier/schematics/sub-blocks
timestamp 1769958744
transform 1 0 9953 0 1 4607
box -953 -807 953 807
use sky130_fd_pr__nfet_g5v0d10v5_986LJA  sky130_fd_pr__nfet_g5v0d10v5_986LJA_1
timestamp 1769958744
transform 1 0 7553 0 1 4607
box -953 -807 953 807
use sky130_fd_pr__nfet_g5v0d10v5_986LJA  sky130_fd_pr__nfet_g5v0d10v5_986LJA_2
timestamp 1769958744
transform 1 0 4753 0 1 4607
box -953 -807 953 807
use sky130_fd_pr__nfet_g5v0d10v5_986LJA  sky130_fd_pr__nfet_g5v0d10v5_986LJA_3
timestamp 1769958744
transform 1 0 2353 0 1 4607
box -953 -807 953 807
use sky130_fd_pr__nfet_g5v0d10v5_R5DZJA  sky130_fd_pr__nfet_g5v0d10v5_R5DZJA_0 /foss/designs/icdec-biomedical-pmic/xschem/error-amplifier/schematics/sub-blocks
timestamp 1769958744
transform 1 0 2353 0 1 2307
box -953 -807 953 807
use sky130_fd_pr__nfet_g5v0d10v5_R5DZJA  sky130_fd_pr__nfet_g5v0d10v5_R5DZJA_1
timestamp 1769958744
transform 1 0 4753 0 1 2307
box -953 -807 953 807
use sky130_fd_pr__nfet_g5v0d10v5_R5DZJA  sky130_fd_pr__nfet_g5v0d10v5_R5DZJA_2
timestamp 1769958744
transform 1 0 7553 0 1 2307
box -953 -807 953 807
use sky130_fd_pr__nfet_g5v0d10v5_R5DZJA  sky130_fd_pr__nfet_g5v0d10v5_R5DZJA_3
timestamp 1769958744
transform 1 0 9953 0 1 2307
box -953 -807 953 807
<< labels >>
flabel metal1 6020 260 6220 460 0 FreeSans 256 0 0 0 IBIAS
port 0 nsew
flabel metal1 800 900 1000 1100 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 6040 6180 6240 6380 0 FreeSans 256 0 0 0 S
port 1 nsew
<< end >>
