magic
tech sky130A
magscale 1 2
timestamp 1769172933
<< mvnmos >>
rect -1623 -719 -1373 781
rect -1195 -719 -945 781
rect -767 -719 -517 781
rect -339 -719 -89 781
rect 89 -719 339 781
rect 517 -719 767 781
rect 945 -719 1195 781
rect 1373 -719 1623 781
<< mvndiff >>
rect -1681 769 -1623 781
rect -1681 -707 -1669 769
rect -1635 -707 -1623 769
rect -1681 -719 -1623 -707
rect -1373 769 -1315 781
rect -1373 -707 -1361 769
rect -1327 -707 -1315 769
rect -1373 -719 -1315 -707
rect -1253 769 -1195 781
rect -1253 -707 -1241 769
rect -1207 -707 -1195 769
rect -1253 -719 -1195 -707
rect -945 769 -887 781
rect -945 -707 -933 769
rect -899 -707 -887 769
rect -945 -719 -887 -707
rect -825 769 -767 781
rect -825 -707 -813 769
rect -779 -707 -767 769
rect -825 -719 -767 -707
rect -517 769 -459 781
rect -517 -707 -505 769
rect -471 -707 -459 769
rect -517 -719 -459 -707
rect -397 769 -339 781
rect -397 -707 -385 769
rect -351 -707 -339 769
rect -397 -719 -339 -707
rect -89 769 -31 781
rect -89 -707 -77 769
rect -43 -707 -31 769
rect -89 -719 -31 -707
rect 31 769 89 781
rect 31 -707 43 769
rect 77 -707 89 769
rect 31 -719 89 -707
rect 339 769 397 781
rect 339 -707 351 769
rect 385 -707 397 769
rect 339 -719 397 -707
rect 459 769 517 781
rect 459 -707 471 769
rect 505 -707 517 769
rect 459 -719 517 -707
rect 767 769 825 781
rect 767 -707 779 769
rect 813 -707 825 769
rect 767 -719 825 -707
rect 887 769 945 781
rect 887 -707 899 769
rect 933 -707 945 769
rect 887 -719 945 -707
rect 1195 769 1253 781
rect 1195 -707 1207 769
rect 1241 -707 1253 769
rect 1195 -719 1253 -707
rect 1315 769 1373 781
rect 1315 -707 1327 769
rect 1361 -707 1373 769
rect 1315 -719 1373 -707
rect 1623 769 1681 781
rect 1623 -707 1635 769
rect 1669 -707 1681 769
rect 1623 -719 1681 -707
<< mvndiffc >>
rect -1669 -707 -1635 769
rect -1361 -707 -1327 769
rect -1241 -707 -1207 769
rect -933 -707 -899 769
rect -813 -707 -779 769
rect -505 -707 -471 769
rect -385 -707 -351 769
rect -77 -707 -43 769
rect 43 -707 77 769
rect 351 -707 385 769
rect 471 -707 505 769
rect 779 -707 813 769
rect 899 -707 933 769
rect 1207 -707 1241 769
rect 1327 -707 1361 769
rect 1635 -707 1669 769
<< poly >>
rect -1623 781 -1373 807
rect -1195 781 -945 807
rect -767 781 -517 807
rect -339 781 -89 807
rect 89 781 339 807
rect 517 781 767 807
rect 945 781 1195 807
rect 1373 781 1623 807
rect -1623 -757 -1373 -719
rect -1623 -791 -1607 -757
rect -1389 -791 -1373 -757
rect -1623 -807 -1373 -791
rect -1195 -757 -945 -719
rect -1195 -791 -1179 -757
rect -961 -791 -945 -757
rect -1195 -807 -945 -791
rect -767 -757 -517 -719
rect -767 -791 -751 -757
rect -533 -791 -517 -757
rect -767 -807 -517 -791
rect -339 -757 -89 -719
rect -339 -791 -323 -757
rect -105 -791 -89 -757
rect -339 -807 -89 -791
rect 89 -757 339 -719
rect 89 -791 105 -757
rect 323 -791 339 -757
rect 89 -807 339 -791
rect 517 -757 767 -719
rect 517 -791 533 -757
rect 751 -791 767 -757
rect 517 -807 767 -791
rect 945 -757 1195 -719
rect 945 -791 961 -757
rect 1179 -791 1195 -757
rect 945 -807 1195 -791
rect 1373 -757 1623 -719
rect 1373 -791 1389 -757
rect 1607 -791 1623 -757
rect 1373 -807 1623 -791
<< polycont >>
rect -1607 -791 -1389 -757
rect -1179 -791 -961 -757
rect -751 -791 -533 -757
rect -323 -791 -105 -757
rect 105 -791 323 -757
rect 533 -791 751 -757
rect 961 -791 1179 -757
rect 1389 -791 1607 -757
<< locali >>
rect -1669 769 -1635 785
rect -1669 -723 -1635 -707
rect -1361 769 -1327 785
rect -1361 -723 -1327 -707
rect -1241 769 -1207 785
rect -1241 -723 -1207 -707
rect -933 769 -899 785
rect -933 -723 -899 -707
rect -813 769 -779 785
rect -813 -723 -779 -707
rect -505 769 -471 785
rect -505 -723 -471 -707
rect -385 769 -351 785
rect -385 -723 -351 -707
rect -77 769 -43 785
rect -77 -723 -43 -707
rect 43 769 77 785
rect 43 -723 77 -707
rect 351 769 385 785
rect 351 -723 385 -707
rect 471 769 505 785
rect 471 -723 505 -707
rect 779 769 813 785
rect 779 -723 813 -707
rect 899 769 933 785
rect 899 -723 933 -707
rect 1207 769 1241 785
rect 1207 -723 1241 -707
rect 1327 769 1361 785
rect 1327 -723 1361 -707
rect 1635 769 1669 785
rect 1635 -723 1669 -707
rect -1623 -791 -1607 -757
rect -1389 -791 -1373 -757
rect -1195 -791 -1179 -757
rect -961 -791 -945 -757
rect -767 -791 -751 -757
rect -533 -791 -517 -757
rect -339 -791 -323 -757
rect -105 -791 -89 -757
rect 89 -791 105 -757
rect 323 -791 339 -757
rect 517 -791 533 -757
rect 751 -791 767 -757
rect 945 -791 961 -757
rect 1179 -791 1195 -757
rect 1373 -791 1389 -757
rect 1607 -791 1623 -757
<< viali >>
rect -1669 -707 -1635 769
rect -1361 -707 -1327 769
rect -1241 -707 -1207 769
rect -933 -707 -899 769
rect -813 -707 -779 769
rect -505 -707 -471 769
rect -385 -707 -351 769
rect -77 -707 -43 769
rect 43 -707 77 769
rect 351 -707 385 769
rect 471 -707 505 769
rect 779 -707 813 769
rect 899 -707 933 769
rect 1207 -707 1241 769
rect 1327 -707 1361 769
rect 1635 -707 1669 769
rect -1607 -791 -1389 -757
rect -1179 -791 -961 -757
rect -751 -791 -533 -757
rect -323 -791 -105 -757
rect 105 -791 323 -757
rect 533 -791 751 -757
rect 961 -791 1179 -757
rect 1389 -791 1607 -757
<< metal1 >>
rect -1675 769 -1629 781
rect -1675 -707 -1669 769
rect -1635 -707 -1629 769
rect -1675 -719 -1629 -707
rect -1367 769 -1321 781
rect -1367 -707 -1361 769
rect -1327 -707 -1321 769
rect -1367 -719 -1321 -707
rect -1247 769 -1201 781
rect -1247 -707 -1241 769
rect -1207 -707 -1201 769
rect -1247 -719 -1201 -707
rect -939 769 -893 781
rect -939 -707 -933 769
rect -899 -707 -893 769
rect -939 -719 -893 -707
rect -819 769 -773 781
rect -819 -707 -813 769
rect -779 -707 -773 769
rect -819 -719 -773 -707
rect -511 769 -465 781
rect -511 -707 -505 769
rect -471 -707 -465 769
rect -511 -719 -465 -707
rect -391 769 -345 781
rect -391 -707 -385 769
rect -351 -707 -345 769
rect -391 -719 -345 -707
rect -83 769 -37 781
rect -83 -707 -77 769
rect -43 -707 -37 769
rect -83 -719 -37 -707
rect 37 769 83 781
rect 37 -707 43 769
rect 77 -707 83 769
rect 37 -719 83 -707
rect 345 769 391 781
rect 345 -707 351 769
rect 385 -707 391 769
rect 345 -719 391 -707
rect 465 769 511 781
rect 465 -707 471 769
rect 505 -707 511 769
rect 465 -719 511 -707
rect 773 769 819 781
rect 773 -707 779 769
rect 813 -707 819 769
rect 773 -719 819 -707
rect 893 769 939 781
rect 893 -707 899 769
rect 933 -707 939 769
rect 893 -719 939 -707
rect 1201 769 1247 781
rect 1201 -707 1207 769
rect 1241 -707 1247 769
rect 1201 -719 1247 -707
rect 1321 769 1367 781
rect 1321 -707 1327 769
rect 1361 -707 1367 769
rect 1321 -719 1367 -707
rect 1629 769 1675 781
rect 1629 -707 1635 769
rect 1669 -707 1675 769
rect 1629 -719 1675 -707
rect -1619 -757 -1377 -751
rect -1619 -791 -1607 -757
rect -1389 -791 -1377 -757
rect -1619 -797 -1377 -791
rect -1191 -757 -949 -751
rect -1191 -791 -1179 -757
rect -961 -791 -949 -757
rect -1191 -797 -949 -791
rect -763 -757 -521 -751
rect -763 -791 -751 -757
rect -533 -791 -521 -757
rect -763 -797 -521 -791
rect -335 -757 -93 -751
rect -335 -791 -323 -757
rect -105 -791 -93 -757
rect -335 -797 -93 -791
rect 93 -757 335 -751
rect 93 -791 105 -757
rect 323 -791 335 -757
rect 93 -797 335 -791
rect 521 -757 763 -751
rect 521 -791 533 -757
rect 751 -791 763 -757
rect 521 -797 763 -791
rect 949 -757 1191 -751
rect 949 -791 961 -757
rect 1179 -791 1191 -757
rect 949 -797 1191 -791
rect 1377 -757 1619 -751
rect 1377 -791 1389 -757
rect 1607 -791 1619 -757
rect 1377 -797 1619 -791
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
