magic
tech sky130A
magscale 1 2
timestamp 1770023980
<< error_p >>
rect -1112 791 -1044 797
rect -804 791 -736 797
rect -496 791 -428 797
rect -188 791 -120 797
rect 120 791 188 797
rect 428 791 496 797
rect 736 791 804 797
rect 1044 791 1112 797
rect -1112 757 -1100 791
rect -804 757 -792 791
rect -496 757 -484 791
rect -188 757 -176 791
rect 120 757 132 791
rect 428 757 440 791
rect 736 757 748 791
rect 1044 757 1056 791
rect -1112 751 -1044 757
rect -804 751 -736 757
rect -496 751 -428 757
rect -188 751 -120 757
rect 120 751 188 757
rect 428 751 496 757
rect 736 751 804 757
rect 1044 751 1112 757
<< mvnmos >>
rect -1203 -781 -953 719
rect -895 -781 -645 719
rect -587 -781 -337 719
rect -279 -781 -29 719
rect 29 -781 279 719
rect 337 -781 587 719
rect 645 -781 895 719
rect 953 -781 1203 719
<< mvndiff >>
rect -1261 707 -1203 719
rect -1261 -769 -1249 707
rect -1215 -769 -1203 707
rect -1261 -781 -1203 -769
rect -953 707 -895 719
rect -953 -769 -941 707
rect -907 -769 -895 707
rect -953 -781 -895 -769
rect -645 707 -587 719
rect -645 -769 -633 707
rect -599 -769 -587 707
rect -645 -781 -587 -769
rect -337 707 -279 719
rect -337 -769 -325 707
rect -291 -769 -279 707
rect -337 -781 -279 -769
rect -29 707 29 719
rect -29 -769 -17 707
rect 17 -769 29 707
rect -29 -781 29 -769
rect 279 707 337 719
rect 279 -769 291 707
rect 325 -769 337 707
rect 279 -781 337 -769
rect 587 707 645 719
rect 587 -769 599 707
rect 633 -769 645 707
rect 587 -781 645 -769
rect 895 707 953 719
rect 895 -769 907 707
rect 941 -769 953 707
rect 895 -781 953 -769
rect 1203 707 1261 719
rect 1203 -769 1215 707
rect 1249 -769 1261 707
rect 1203 -781 1261 -769
<< mvndiffc >>
rect -1249 -769 -1215 707
rect -941 -769 -907 707
rect -633 -769 -599 707
rect -325 -769 -291 707
rect -17 -769 17 707
rect 291 -769 325 707
rect 599 -769 633 707
rect 907 -769 941 707
rect 1215 -769 1249 707
<< poly >>
rect -1116 791 -1040 807
rect -1116 774 -1100 791
rect -1203 757 -1100 774
rect -1056 774 -1040 791
rect -808 791 -732 807
rect -808 774 -792 791
rect -1056 757 -953 774
rect -1203 719 -953 757
rect -895 757 -792 774
rect -748 774 -732 791
rect -500 791 -424 807
rect -500 774 -484 791
rect -748 757 -645 774
rect -895 719 -645 757
rect -587 757 -484 774
rect -440 774 -424 791
rect -192 791 -116 807
rect -192 774 -176 791
rect -440 757 -337 774
rect -587 719 -337 757
rect -279 757 -176 774
rect -132 774 -116 791
rect 116 791 192 807
rect 116 774 132 791
rect -132 757 -29 774
rect -279 719 -29 757
rect 29 757 132 774
rect 176 774 192 791
rect 424 791 500 807
rect 424 774 440 791
rect 176 757 279 774
rect 29 719 279 757
rect 337 757 440 774
rect 484 774 500 791
rect 732 791 808 807
rect 732 774 748 791
rect 484 757 587 774
rect 337 719 587 757
rect 645 757 748 774
rect 792 774 808 791
rect 1040 791 1116 807
rect 1040 774 1056 791
rect 792 757 895 774
rect 645 719 895 757
rect 953 757 1056 774
rect 1100 774 1116 791
rect 1100 757 1203 774
rect 953 719 1203 757
rect -1203 -807 -953 -781
rect -895 -807 -645 -781
rect -587 -807 -337 -781
rect -279 -807 -29 -781
rect 29 -807 279 -781
rect 337 -807 587 -781
rect 645 -807 895 -781
rect 953 -807 1203 -781
<< polycont >>
rect -1100 757 -1056 791
rect -792 757 -748 791
rect -484 757 -440 791
rect -176 757 -132 791
rect 132 757 176 791
rect 440 757 484 791
rect 748 757 792 791
rect 1056 757 1100 791
<< locali >>
rect -1116 757 -1100 791
rect -1056 757 -1040 791
rect -808 757 -792 791
rect -748 757 -732 791
rect -500 757 -484 791
rect -440 757 -424 791
rect -192 757 -176 791
rect -132 757 -116 791
rect 116 757 132 791
rect 176 757 192 791
rect 424 757 440 791
rect 484 757 500 791
rect 732 757 748 791
rect 792 757 808 791
rect 1040 757 1056 791
rect 1100 757 1116 791
rect -1249 707 -1215 723
rect -1249 -785 -1215 -769
rect -941 707 -907 723
rect -941 -785 -907 -769
rect -633 707 -599 723
rect -633 -785 -599 -769
rect -325 707 -291 723
rect -325 -785 -291 -769
rect -17 707 17 723
rect -17 -785 17 -769
rect 291 707 325 723
rect 291 -785 325 -769
rect 599 707 633 723
rect 599 -785 633 -769
rect 907 707 941 723
rect 907 -785 941 -769
rect 1215 707 1249 723
rect 1215 -785 1249 -769
<< viali >>
rect -1100 757 -1056 791
rect -792 757 -748 791
rect -484 757 -440 791
rect -176 757 -132 791
rect 132 757 176 791
rect 440 757 484 791
rect 748 757 792 791
rect 1056 757 1100 791
rect -1249 -769 -1215 707
rect -941 -769 -907 707
rect -633 -769 -599 707
rect -325 -769 -291 707
rect -17 -769 17 707
rect 291 -769 325 707
rect 599 -769 633 707
rect 907 -769 941 707
rect 1215 -769 1249 707
<< metal1 >>
rect -1112 791 -1044 797
rect -1112 757 -1100 791
rect -1056 757 -1044 791
rect -1112 751 -1044 757
rect -804 791 -736 797
rect -804 757 -792 791
rect -748 757 -736 791
rect -804 751 -736 757
rect -496 791 -428 797
rect -496 757 -484 791
rect -440 757 -428 791
rect -496 751 -428 757
rect -188 791 -120 797
rect -188 757 -176 791
rect -132 757 -120 791
rect -188 751 -120 757
rect 120 791 188 797
rect 120 757 132 791
rect 176 757 188 791
rect 120 751 188 757
rect 428 791 496 797
rect 428 757 440 791
rect 484 757 496 791
rect 428 751 496 757
rect 736 791 804 797
rect 736 757 748 791
rect 792 757 804 791
rect 736 751 804 757
rect 1044 791 1112 797
rect 1044 757 1056 791
rect 1100 757 1112 791
rect 1044 751 1112 757
rect -1255 707 -1209 719
rect -1255 -769 -1249 707
rect -1215 -769 -1209 707
rect -1255 -781 -1209 -769
rect -947 707 -901 719
rect -947 -769 -941 707
rect -907 -769 -901 707
rect -947 -781 -901 -769
rect -639 707 -593 719
rect -639 -769 -633 707
rect -599 -769 -593 707
rect -639 -781 -593 -769
rect -331 707 -285 719
rect -331 -769 -325 707
rect -291 -769 -285 707
rect -331 -781 -285 -769
rect -23 707 23 719
rect -23 -769 -17 707
rect 17 200 23 707
rect 285 707 331 719
rect 17 0 200 200
rect 17 -200 23 0
rect 17 -400 200 -200
rect 17 -600 23 -400
rect 17 -769 200 -600
rect -23 -781 200 -769
rect 285 -769 291 707
rect 325 -769 331 707
rect 285 -781 331 -769
rect 593 707 639 719
rect 593 -769 599 707
rect 633 -769 639 707
rect 593 -781 639 -769
rect 901 707 947 719
rect 901 -769 907 707
rect 941 -769 947 707
rect 901 -781 947 -769
rect 1209 707 1255 719
rect 1209 -769 1215 707
rect 1249 -769 1255 707
rect 1209 -781 1255 -769
rect 0 -800 200 -781
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X0
timestamp 0
transform 1 0 -973 0 1 -7057
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X1
timestamp 0
transform 1 0 -332 0 1 -7122
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X2
timestamp 0
transform 1 0 309 0 1 -7187
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_X6YUYU  X3
timestamp 0
transform 1 0 950 0 1 -7252
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_XZ8YPJ  X4
timestamp 0
transform 1 0 1591 0 1 -7317
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X5
timestamp 0
transform 1 0 2232 0 1 -7382
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X6
timestamp 0
transform 1 0 2873 0 1 -7447
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_ZX75FA  X7
timestamp 0
transform 1 0 3514 0 1 -7512
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 a_n953_n781#
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 a_n587_n807#
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 a_645_n807#
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 {}
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 a_29_n807#
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 a_279_n781#
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 a_895_n781#
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 a_n1261_n781#
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 a_n29_n781#
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 a_n645_n781#
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 a_n279_n807#
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 a_n895_n807#
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 a_337_n807#
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 a_953_n807#
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 a_587_n781#
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 a_1203_n781#
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 a_n337_n781#
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 a_n1203_n807#
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 {}
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 VSUBS
port 20 nsew
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 8 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
