magic
tech sky130A
magscale 1 2
timestamp 1770123317
<< pwell >>
rect -825 -558 825 558
<< mvnmos >>
rect -595 -300 -445 300
rect -387 -300 -237 300
rect -179 -300 -29 300
rect 29 -300 179 300
rect 237 -300 387 300
rect 445 -300 595 300
<< mvndiff >>
rect -653 288 -595 300
rect -653 -288 -641 288
rect -607 -288 -595 288
rect -653 -300 -595 -288
rect -445 288 -387 300
rect -445 -288 -433 288
rect -399 -288 -387 288
rect -445 -300 -387 -288
rect -237 288 -179 300
rect -237 -288 -225 288
rect -191 -288 -179 288
rect -237 -300 -179 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 179 288 237 300
rect 179 -288 191 288
rect 225 -288 237 288
rect 179 -300 237 -288
rect 387 288 445 300
rect 387 -288 399 288
rect 433 -288 445 288
rect 387 -300 445 -288
rect 595 288 653 300
rect 595 -288 607 288
rect 641 -288 653 288
rect 595 -300 653 -288
<< mvndiffc >>
rect -641 -288 -607 288
rect -433 -288 -399 288
rect -225 -288 -191 288
rect -17 -288 17 288
rect 191 -288 225 288
rect 399 -288 433 288
rect 607 -288 641 288
<< mvpsubdiff >>
rect -789 510 789 522
rect -789 476 -681 510
rect 681 476 789 510
rect -789 464 789 476
rect -789 -464 -731 464
rect 731 -464 789 464
rect -789 -476 789 -464
rect -789 -510 -681 -476
rect 681 -510 789 -476
rect -789 -522 789 -510
<< mvpsubdiffcont >>
rect -681 476 681 510
rect -681 -510 681 -476
<< poly >>
rect -595 372 -445 388
rect -595 338 -579 372
rect -461 338 -445 372
rect -595 300 -445 338
rect -387 372 -237 388
rect -387 338 -371 372
rect -253 338 -237 372
rect -387 300 -237 338
rect -179 372 -29 388
rect -179 338 -163 372
rect -45 338 -29 372
rect -179 300 -29 338
rect 29 372 179 388
rect 29 338 45 372
rect 163 338 179 372
rect 29 300 179 338
rect 237 372 387 388
rect 237 338 253 372
rect 371 338 387 372
rect 237 300 387 338
rect 445 372 595 388
rect 445 338 461 372
rect 579 338 595 372
rect 445 300 595 338
rect -595 -338 -445 -300
rect -595 -372 -579 -338
rect -461 -372 -445 -338
rect -595 -388 -445 -372
rect -387 -338 -237 -300
rect -387 -372 -371 -338
rect -253 -372 -237 -338
rect -387 -388 -237 -372
rect -179 -338 -29 -300
rect -179 -372 -163 -338
rect -45 -372 -29 -338
rect -179 -388 -29 -372
rect 29 -338 179 -300
rect 29 -372 45 -338
rect 163 -372 179 -338
rect 29 -388 179 -372
rect 237 -338 387 -300
rect 237 -372 253 -338
rect 371 -372 387 -338
rect 237 -388 387 -372
rect 445 -338 595 -300
rect 445 -372 461 -338
rect 579 -372 595 -338
rect 445 -388 595 -372
<< polycont >>
rect -579 338 -461 372
rect -371 338 -253 372
rect -163 338 -45 372
rect 45 338 163 372
rect 253 338 371 372
rect 461 338 579 372
rect -579 -372 -461 -338
rect -371 -372 -253 -338
rect -163 -372 -45 -338
rect 45 -372 163 -338
rect 253 -372 371 -338
rect 461 -372 579 -338
<< locali >>
rect -777 476 -681 510
rect 681 476 777 510
rect -777 -476 -743 476
rect -595 338 -579 372
rect -461 338 -445 372
rect -387 338 -371 372
rect -253 338 -237 372
rect -179 338 -163 372
rect -45 338 -29 372
rect 29 338 45 372
rect 163 338 179 372
rect 237 338 253 372
rect 371 338 387 372
rect 445 338 461 372
rect 579 338 595 372
rect -641 288 -607 304
rect -641 -304 -607 -288
rect -433 288 -399 304
rect -433 -304 -399 -288
rect -225 288 -191 304
rect -225 -304 -191 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 191 288 225 304
rect 191 -304 225 -288
rect 399 288 433 304
rect 399 -304 433 -288
rect 607 288 641 304
rect 607 -304 641 -288
rect -595 -372 -579 -338
rect -461 -372 -445 -338
rect -387 -372 -371 -338
rect -253 -372 -237 -338
rect -179 -372 -163 -338
rect -45 -372 -29 -338
rect 29 -372 45 -338
rect 163 -372 179 -338
rect 237 -372 253 -338
rect 371 -372 387 -338
rect 445 -372 461 -338
rect 579 -372 595 -338
rect 743 -476 777 476
rect -777 -510 -681 -476
rect 681 -510 777 -476
<< viali >>
rect -579 338 -461 372
rect -371 338 -253 372
rect -163 338 -45 372
rect 45 338 163 372
rect 253 338 371 372
rect 461 338 579 372
rect -641 -288 -607 288
rect -433 -288 -399 288
rect -225 -288 -191 288
rect -17 -288 17 288
rect 191 -288 225 288
rect 399 -288 433 288
rect 607 -288 641 288
rect -579 -372 -461 -338
rect -371 -372 -253 -338
rect -163 -372 -45 -338
rect 45 -372 163 -338
rect 253 -372 371 -338
rect 461 -372 579 -338
<< metal1 >>
rect -591 372 -449 378
rect -591 338 -579 372
rect -461 338 -449 372
rect -591 332 -449 338
rect -383 372 -241 378
rect -383 338 -371 372
rect -253 338 -241 372
rect -383 332 -241 338
rect -175 372 -33 378
rect -175 338 -163 372
rect -45 338 -33 372
rect -175 332 -33 338
rect 33 372 175 378
rect 33 338 45 372
rect 163 338 175 372
rect 33 332 175 338
rect 241 372 383 378
rect 241 338 253 372
rect 371 338 383 372
rect 241 332 383 338
rect 449 372 591 378
rect 449 338 461 372
rect 579 338 591 372
rect 449 332 591 338
rect -647 288 -601 300
rect -647 -288 -641 288
rect -607 -288 -601 288
rect -647 -300 -601 -288
rect -439 288 -393 300
rect -439 -288 -433 288
rect -399 -288 -393 288
rect -439 -300 -393 -288
rect -231 288 -185 300
rect -231 -288 -225 288
rect -191 -288 -185 288
rect -231 -300 -185 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 185 288 231 300
rect 185 -288 191 288
rect 225 -288 231 288
rect 185 -300 231 -288
rect 393 288 439 300
rect 393 -288 399 288
rect 433 -288 439 288
rect 393 -300 439 -288
rect 601 288 647 300
rect 601 -288 607 288
rect 641 -288 647 288
rect 601 -300 647 -288
rect -591 -338 -449 -332
rect -591 -372 -579 -338
rect -461 -372 -449 -338
rect -591 -378 -449 -372
rect -383 -338 -241 -332
rect -383 -372 -371 -338
rect -253 -372 -241 -338
rect -383 -378 -241 -372
rect -175 -338 -33 -332
rect -175 -372 -163 -338
rect -45 -372 -33 -338
rect -175 -378 -33 -372
rect 33 -338 175 -332
rect 33 -372 45 -338
rect 163 -372 175 -338
rect 33 -378 175 -372
rect 241 -338 383 -332
rect 241 -372 253 -338
rect 371 -372 383 -338
rect 241 -378 383 -372
rect 449 -338 591 -332
rect 449 -372 461 -338
rect 579 -372 591 -338
rect 449 -378 591 -372
<< labels >>
rlabel mvpsubdiffcont 0 -493 0 -493 0 B
port 1 nsew
rlabel mvndiffc -624 0 -624 0 0 D0
port 2 nsew
rlabel polycont -520 355 -520 355 0 G0
port 3 nsew
rlabel mvndiffc -416 0 -416 0 0 S1
port 4 nsew
rlabel polycont -312 355 -312 355 0 G1
port 5 nsew
rlabel mvndiffc -208 0 -208 0 0 D2
port 6 nsew
rlabel polycont -104 355 -104 355 0 G2
port 7 nsew
rlabel mvndiffc 0 0 0 0 0 S3
port 8 nsew
rlabel polycont 104 355 104 355 0 G3
port 9 nsew
rlabel mvndiffc 208 0 208 0 0 D4
port 10 nsew
rlabel polycont 312 355 312 355 0 G4
port 11 nsew
rlabel mvndiffc 416 0 416 0 0 S5
port 12 nsew
rlabel polycont 520 355 520 355 0 G5
port 13 nsew
<< properties >>
string FIXED_BBOX -760 -493 760 493
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 0.75 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
