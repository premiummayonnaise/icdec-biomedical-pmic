magic
tech sky130A
magscale 1 2
timestamp 1769436194
<< pwell >>
rect -451 -18294 451 18294
<< psubdiff >>
rect -415 18224 -319 18258
rect 319 18224 415 18258
rect -415 18162 -381 18224
rect 381 18162 415 18224
rect -415 -18224 -381 -18162
rect 381 -18224 415 -18162
rect -415 -18258 -319 -18224
rect 319 -18258 415 -18224
<< psubdiffcont >>
rect -319 18224 319 18258
rect -415 -18162 -381 18162
rect 381 -18162 415 18162
rect -319 -18258 319 -18224
<< xpolycontact >>
rect -285 17696 285 18128
rect -285 14596 285 15028
rect -285 14060 285 14492
rect -285 10960 285 11392
rect -285 10424 285 10856
rect -285 7324 285 7756
rect -285 6788 285 7220
rect -285 3688 285 4120
rect -285 3152 285 3584
rect -285 52 285 484
rect -285 -484 285 -52
rect -285 -3584 285 -3152
rect -285 -4120 285 -3688
rect -285 -7220 285 -6788
rect -285 -7756 285 -7324
rect -285 -10856 285 -10424
rect -285 -11392 285 -10960
rect -285 -14492 285 -14060
rect -285 -15028 285 -14596
rect -285 -18128 285 -17696
<< ppolyres >>
rect -285 15028 285 17696
rect -285 11392 285 14060
rect -285 7756 285 10424
rect -285 4120 285 6788
rect -285 484 285 3152
rect -285 -3152 285 -484
rect -285 -6788 285 -4120
rect -285 -10424 285 -7756
rect -285 -14060 285 -11392
rect -285 -17696 285 -15028
<< locali >>
rect -415 18224 -319 18258
rect 319 18224 415 18258
rect -415 18162 -381 18224
rect 381 18162 415 18224
rect -415 -18224 -381 -18162
rect 381 -18224 415 -18162
rect -415 -18258 -319 -18224
rect 319 -18258 415 -18224
<< viali >>
rect -269 17713 269 18110
rect -269 14614 269 15011
rect -269 14077 269 14474
rect -269 10978 269 11375
rect -269 10441 269 10838
rect -269 7342 269 7739
rect -269 6805 269 7202
rect -269 3706 269 4103
rect -269 3169 269 3566
rect -269 70 269 467
rect -269 -467 269 -70
rect -269 -3566 269 -3169
rect -269 -4103 269 -3706
rect -269 -7202 269 -6805
rect -269 -7739 269 -7342
rect -269 -10838 269 -10441
rect -269 -11375 269 -10978
rect -269 -14474 269 -14077
rect -269 -15011 269 -14614
rect -269 -18110 269 -17713
<< metal1 >>
rect -281 18110 281 18116
rect -281 17713 -269 18110
rect 269 17713 281 18110
rect -281 17707 281 17713
rect -281 15011 281 15017
rect -281 14614 -269 15011
rect 269 14614 281 15011
rect -281 14608 281 14614
rect -281 14474 281 14480
rect -281 14077 -269 14474
rect 269 14077 281 14474
rect -281 14071 281 14077
rect -281 11375 281 11381
rect -281 10978 -269 11375
rect 269 10978 281 11375
rect -281 10972 281 10978
rect -281 10838 281 10844
rect -281 10441 -269 10838
rect 269 10441 281 10838
rect -281 10435 281 10441
rect -281 7739 281 7745
rect -281 7342 -269 7739
rect 269 7342 281 7739
rect -281 7336 281 7342
rect -281 7202 281 7208
rect -281 6805 -269 7202
rect 269 6805 281 7202
rect -281 6799 281 6805
rect -281 4103 281 4109
rect -281 3706 -269 4103
rect 269 3706 281 4103
rect -281 3700 281 3706
rect -281 3566 281 3572
rect -281 3169 -269 3566
rect 269 3169 281 3566
rect -281 3163 281 3169
rect -281 467 281 473
rect -281 70 -269 467
rect 269 70 281 467
rect -281 64 281 70
rect -281 -70 281 -64
rect -281 -467 -269 -70
rect 269 -467 281 -70
rect -281 -473 281 -467
rect -281 -3169 281 -3163
rect -281 -3566 -269 -3169
rect 269 -3566 281 -3169
rect -281 -3572 281 -3566
rect -281 -3706 281 -3700
rect -281 -4103 -269 -3706
rect 269 -4103 281 -3706
rect -281 -4109 281 -4103
rect -281 -6805 281 -6799
rect -281 -7202 -269 -6805
rect 269 -7202 281 -6805
rect -281 -7208 281 -7202
rect -281 -7342 281 -7336
rect -281 -7739 -269 -7342
rect 269 -7739 281 -7342
rect -281 -7745 281 -7739
rect -281 -10441 281 -10435
rect -281 -10838 -269 -10441
rect 269 -10838 281 -10441
rect -281 -10844 281 -10838
rect -281 -10978 281 -10972
rect -281 -11375 -269 -10978
rect 269 -11375 281 -10978
rect -281 -11381 281 -11375
rect -281 -14077 281 -14071
rect -281 -14474 -269 -14077
rect 269 -14474 281 -14077
rect -281 -14480 281 -14474
rect -281 -14614 281 -14608
rect -281 -15011 -269 -14614
rect 269 -15011 281 -14614
rect -281 -15017 281 -15011
rect -281 -17713 281 -17707
rect -281 -18110 -269 -17713
rect 269 -18110 281 -17713
rect -281 -18116 281 -18110
<< properties >>
string FIXED_BBOX -398 -18241 398 18241
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string parameters w 2.850 l 13.5 m 10 nx 1 wmin 2.850 lmin 0.50 class resistor rho 319.8 val 1.651k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 2.850 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
