* =============================================================
* tb_ac_pex.spice
* PEX-backed AC testbench for two-stage-miller (sky130A)
* =============================================================

.GLOBAL GND

* --- Models / Corner ---
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice ss

* --- Include extracted PEX netlist ---
.include "two-stage-miller_pex.spice"

* =============================================================
* Testbench sources (TOP LEVEL — NOT a subckt)
* =============================================================

* Differential input
V2 VN  VSS ac -1m dc 1.25
V3 VP  VSS ac  1m dc 1.25

* Supplies
V5 VDD VSS 5
V7 VSS GND 0

* Bias
I4 VDD IBIAS 200u

* Output loading
C2 OUT  VSS 1p

* Common-mode path
V1 VCM VSS ac 1m DC 0.9
C1 OUT2 VSS 5p

* PSRR path
V4 VDDr VSS DC 5 AC 1
C3 OUT3 VSS 10p
R1 OUT3 VN 1k

* =============================================================
* DUT instantiations (PEX-backed)
* =============================================================

x1 VDD  OUT  VP  VN  IBIAS VSS two-stage-miller
x2 VDD  OUT2 VCM VCM IBIAS VSS two-stage-miller
x3 VDDr OUT3 VP  VN  IBIAS VSS two-stage-miller

* =============================================================
* Control block (MUST be top-level)
* =============================================================

.control
  .temp 27
  op
  ac dec 100 1 100MEG
  save all

  let vd = v(vp) - v(vn)
  let Av = db( v(OUT) / vd)
  let phase = 180*cph( v(OUT) )/pi

  meas ac f_0db when Av = 0
  meas ac phase_at_unity find phase when Av = 0

  let p_total = v(vdd) * i(Vdd)

  let Acm = db( v(OUT2)/vcm)
  let cmrr = Av - Acm
  let psrr = -20*log10(OUT3)

  print f_0db phase_at_unity
  plot psrr
  plot av
  plot acm
  plot cmrr
  plot phase
  plot p_total
.endc

.end
