magic
tech sky130A
magscale 1 2
timestamp 1770003475
<< pwell >>
rect -353 -1008 353 1008
<< mvnmos >>
rect -125 -750 125 750
<< mvndiff >>
rect -183 738 -125 750
rect -183 -738 -171 738
rect -137 -738 -125 738
rect -183 -750 -125 -738
rect 125 738 183 750
rect 125 -738 137 738
rect 171 -738 183 738
rect 125 -750 183 -738
<< mvndiffc >>
rect -171 -738 -137 738
rect 137 -738 171 738
<< mvpsubdiff >>
rect -317 960 317 972
rect -317 926 -209 960
rect 209 926 317 960
rect -317 914 317 926
rect -317 864 -259 914
rect -317 -864 -305 864
rect -271 -864 -259 864
rect 259 864 317 914
rect -317 -914 -259 -864
rect 259 -864 271 864
rect 305 -864 317 864
rect 259 -914 317 -864
rect -317 -926 317 -914
rect -317 -960 -209 -926
rect 209 -960 317 -926
rect -317 -972 317 -960
<< mvpsubdiffcont >>
rect -209 926 209 960
rect -305 -864 -271 864
rect 271 -864 305 864
rect -209 -960 209 -926
<< poly >>
rect -125 822 125 838
rect -125 788 -109 822
rect 109 788 125 822
rect -125 750 125 788
rect -125 -788 125 -750
rect -125 -822 -109 -788
rect 109 -822 125 -788
rect -125 -838 125 -822
<< polycont >>
rect -109 788 109 822
rect -109 -822 109 -788
<< locali >>
rect -305 926 -209 960
rect 209 926 305 960
rect -305 864 -271 926
rect 271 864 305 926
rect -125 788 -109 822
rect 109 788 125 822
rect -171 738 -137 754
rect -171 -754 -137 -738
rect 137 738 171 754
rect 137 -754 171 -738
rect -125 -822 -109 -788
rect 109 -822 125 -788
rect -305 -926 -271 -864
rect 271 -926 305 -864
rect -305 -960 -209 -926
rect 209 -960 305 -926
<< viali >>
rect -109 788 109 822
rect -171 -738 -137 738
rect 137 -738 171 738
rect -109 -822 109 -788
<< metal1 >>
rect -121 822 121 828
rect -121 788 -109 822
rect 109 788 121 822
rect -121 782 121 788
rect -177 738 -131 750
rect -177 -738 -171 738
rect -137 -738 -131 738
rect -177 -750 -131 -738
rect 131 738 177 750
rect 131 -738 137 738
rect 171 -738 177 738
rect 131 -750 177 -738
rect -121 -788 121 -782
rect -121 -822 -109 -788
rect 109 -822 121 -788
rect -121 -828 121 -822
<< properties >>
string FIXED_BBOX -288 -943 288 943
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
