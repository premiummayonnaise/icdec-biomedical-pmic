magic
tech sky130A
magscale 1 2
timestamp 1769135993
<< nwell >>
rect -1415 -414 1415 414
<< pmos >>
rect -1219 -195 -1069 195
rect -1011 -195 -861 195
rect -803 -195 -653 195
rect -595 -195 -445 195
rect -387 -195 -237 195
rect -179 -195 -29 195
rect 29 -195 179 195
rect 237 -195 387 195
rect 445 -195 595 195
rect 653 -195 803 195
rect 861 -195 1011 195
rect 1069 -195 1219 195
<< pdiff >>
rect -1277 183 -1219 195
rect -1277 -183 -1265 183
rect -1231 -183 -1219 183
rect -1277 -195 -1219 -183
rect -1069 183 -1011 195
rect -1069 -183 -1057 183
rect -1023 -183 -1011 183
rect -1069 -195 -1011 -183
rect -861 183 -803 195
rect -861 -183 -849 183
rect -815 -183 -803 183
rect -861 -195 -803 -183
rect -653 183 -595 195
rect -653 -183 -641 183
rect -607 -183 -595 183
rect -653 -195 -595 -183
rect -445 183 -387 195
rect -445 -183 -433 183
rect -399 -183 -387 183
rect -445 -195 -387 -183
rect -237 183 -179 195
rect -237 -183 -225 183
rect -191 -183 -179 183
rect -237 -195 -179 -183
rect -29 183 29 195
rect -29 -183 -17 183
rect 17 -183 29 183
rect -29 -195 29 -183
rect 179 183 237 195
rect 179 -183 191 183
rect 225 -183 237 183
rect 179 -195 237 -183
rect 387 183 445 195
rect 387 -183 399 183
rect 433 -183 445 183
rect 387 -195 445 -183
rect 595 183 653 195
rect 595 -183 607 183
rect 641 -183 653 183
rect 595 -195 653 -183
rect 803 183 861 195
rect 803 -183 815 183
rect 849 -183 861 183
rect 803 -195 861 -183
rect 1011 183 1069 195
rect 1011 -183 1023 183
rect 1057 -183 1069 183
rect 1011 -195 1069 -183
rect 1219 183 1277 195
rect 1219 -183 1231 183
rect 1265 -183 1277 183
rect 1219 -195 1277 -183
<< pdiffc >>
rect -1265 -183 -1231 183
rect -1057 -183 -1023 183
rect -849 -183 -815 183
rect -641 -183 -607 183
rect -433 -183 -399 183
rect -225 -183 -191 183
rect -17 -183 17 183
rect 191 -183 225 183
rect 399 -183 433 183
rect 607 -183 641 183
rect 815 -183 849 183
rect 1023 -183 1057 183
rect 1231 -183 1265 183
<< nsubdiff >>
rect -1379 344 -1283 378
rect 1283 344 1379 378
rect -1379 282 -1345 344
rect 1345 282 1379 344
rect -1379 -344 -1345 -282
rect 1345 -344 1379 -282
rect -1379 -378 -1283 -344
rect 1283 -378 1379 -344
<< nsubdiffcont >>
rect -1283 344 1283 378
rect -1379 -282 -1345 282
rect 1345 -282 1379 282
rect -1283 -378 1283 -344
<< poly >>
rect -1219 276 -1069 292
rect -1219 242 -1203 276
rect -1085 242 -1069 276
rect -1219 195 -1069 242
rect -1011 276 -861 292
rect -1011 242 -995 276
rect -877 242 -861 276
rect -1011 195 -861 242
rect -803 276 -653 292
rect -803 242 -787 276
rect -669 242 -653 276
rect -803 195 -653 242
rect -595 276 -445 292
rect -595 242 -579 276
rect -461 242 -445 276
rect -595 195 -445 242
rect -387 276 -237 292
rect -387 242 -371 276
rect -253 242 -237 276
rect -387 195 -237 242
rect -179 276 -29 292
rect -179 242 -163 276
rect -45 242 -29 276
rect -179 195 -29 242
rect 29 276 179 292
rect 29 242 45 276
rect 163 242 179 276
rect 29 195 179 242
rect 237 276 387 292
rect 237 242 253 276
rect 371 242 387 276
rect 237 195 387 242
rect 445 276 595 292
rect 445 242 461 276
rect 579 242 595 276
rect 445 195 595 242
rect 653 276 803 292
rect 653 242 669 276
rect 787 242 803 276
rect 653 195 803 242
rect 861 276 1011 292
rect 861 242 877 276
rect 995 242 1011 276
rect 861 195 1011 242
rect 1069 276 1219 292
rect 1069 242 1085 276
rect 1203 242 1219 276
rect 1069 195 1219 242
rect -1219 -242 -1069 -195
rect -1219 -276 -1203 -242
rect -1085 -276 -1069 -242
rect -1219 -292 -1069 -276
rect -1011 -242 -861 -195
rect -1011 -276 -995 -242
rect -877 -276 -861 -242
rect -1011 -292 -861 -276
rect -803 -242 -653 -195
rect -803 -276 -787 -242
rect -669 -276 -653 -242
rect -803 -292 -653 -276
rect -595 -242 -445 -195
rect -595 -276 -579 -242
rect -461 -276 -445 -242
rect -595 -292 -445 -276
rect -387 -242 -237 -195
rect -387 -276 -371 -242
rect -253 -276 -237 -242
rect -387 -292 -237 -276
rect -179 -242 -29 -195
rect -179 -276 -163 -242
rect -45 -276 -29 -242
rect -179 -292 -29 -276
rect 29 -242 179 -195
rect 29 -276 45 -242
rect 163 -276 179 -242
rect 29 -292 179 -276
rect 237 -242 387 -195
rect 237 -276 253 -242
rect 371 -276 387 -242
rect 237 -292 387 -276
rect 445 -242 595 -195
rect 445 -276 461 -242
rect 579 -276 595 -242
rect 445 -292 595 -276
rect 653 -242 803 -195
rect 653 -276 669 -242
rect 787 -276 803 -242
rect 653 -292 803 -276
rect 861 -242 1011 -195
rect 861 -276 877 -242
rect 995 -276 1011 -242
rect 861 -292 1011 -276
rect 1069 -242 1219 -195
rect 1069 -276 1085 -242
rect 1203 -276 1219 -242
rect 1069 -292 1219 -276
<< polycont >>
rect -1203 242 -1085 276
rect -995 242 -877 276
rect -787 242 -669 276
rect -579 242 -461 276
rect -371 242 -253 276
rect -163 242 -45 276
rect 45 242 163 276
rect 253 242 371 276
rect 461 242 579 276
rect 669 242 787 276
rect 877 242 995 276
rect 1085 242 1203 276
rect -1203 -276 -1085 -242
rect -995 -276 -877 -242
rect -787 -276 -669 -242
rect -579 -276 -461 -242
rect -371 -276 -253 -242
rect -163 -276 -45 -242
rect 45 -276 163 -242
rect 253 -276 371 -242
rect 461 -276 579 -242
rect 669 -276 787 -242
rect 877 -276 995 -242
rect 1085 -276 1203 -242
<< locali >>
rect -1379 344 -1283 378
rect 1283 344 1379 378
rect -1379 282 -1345 344
rect 1345 282 1379 344
rect -1219 242 -1203 276
rect -1085 242 -1069 276
rect -1011 242 -995 276
rect -877 242 -861 276
rect -803 242 -787 276
rect -669 242 -653 276
rect -595 242 -579 276
rect -461 242 -445 276
rect -387 242 -371 276
rect -253 242 -237 276
rect -179 242 -163 276
rect -45 242 -29 276
rect 29 242 45 276
rect 163 242 179 276
rect 237 242 253 276
rect 371 242 387 276
rect 445 242 461 276
rect 579 242 595 276
rect 653 242 669 276
rect 787 242 803 276
rect 861 242 877 276
rect 995 242 1011 276
rect 1069 242 1085 276
rect 1203 242 1219 276
rect -1265 183 -1231 199
rect -1265 -199 -1231 -183
rect -1057 183 -1023 199
rect -1057 -199 -1023 -183
rect -849 183 -815 199
rect -849 -199 -815 -183
rect -641 183 -607 199
rect -641 -199 -607 -183
rect -433 183 -399 199
rect -433 -199 -399 -183
rect -225 183 -191 199
rect -225 -199 -191 -183
rect -17 183 17 199
rect -17 -199 17 -183
rect 191 183 225 199
rect 191 -199 225 -183
rect 399 183 433 199
rect 399 -199 433 -183
rect 607 183 641 199
rect 607 -199 641 -183
rect 815 183 849 199
rect 815 -199 849 -183
rect 1023 183 1057 199
rect 1023 -199 1057 -183
rect 1231 183 1265 199
rect 1231 -199 1265 -183
rect -1219 -276 -1203 -242
rect -1085 -276 -1069 -242
rect -1011 -276 -995 -242
rect -877 -276 -861 -242
rect -803 -276 -787 -242
rect -669 -276 -653 -242
rect -595 -276 -579 -242
rect -461 -276 -445 -242
rect -387 -276 -371 -242
rect -253 -276 -237 -242
rect -179 -276 -163 -242
rect -45 -276 -29 -242
rect 29 -276 45 -242
rect 163 -276 179 -242
rect 237 -276 253 -242
rect 371 -276 387 -242
rect 445 -276 461 -242
rect 579 -276 595 -242
rect 653 -276 669 -242
rect 787 -276 803 -242
rect 861 -276 877 -242
rect 995 -276 1011 -242
rect 1069 -276 1085 -242
rect 1203 -276 1219 -242
rect -1379 -344 -1345 -282
rect 1345 -344 1379 -282
rect -1379 -378 -1283 -344
rect 1283 -378 1379 -344
<< viali >>
rect -1203 242 -1085 276
rect -995 242 -877 276
rect -787 242 -669 276
rect -579 242 -461 276
rect -371 242 -253 276
rect -163 242 -45 276
rect 45 242 163 276
rect 253 242 371 276
rect 461 242 579 276
rect 669 242 787 276
rect 877 242 995 276
rect 1085 242 1203 276
rect -1265 -183 -1231 183
rect -1057 -183 -1023 183
rect -849 -183 -815 183
rect -641 -183 -607 183
rect -433 -183 -399 183
rect -225 -183 -191 183
rect -17 -183 17 183
rect 191 -183 225 183
rect 399 -183 433 183
rect 607 -183 641 183
rect 815 -183 849 183
rect 1023 -183 1057 183
rect 1231 -183 1265 183
rect -1203 -276 -1085 -242
rect -995 -276 -877 -242
rect -787 -276 -669 -242
rect -579 -276 -461 -242
rect -371 -276 -253 -242
rect -163 -276 -45 -242
rect 45 -276 163 -242
rect 253 -276 371 -242
rect 461 -276 579 -242
rect 669 -276 787 -242
rect 877 -276 995 -242
rect 1085 -276 1203 -242
<< metal1 >>
rect -1215 276 -1073 282
rect -1215 242 -1203 276
rect -1085 242 -1073 276
rect -1215 236 -1073 242
rect -1007 276 -865 282
rect -1007 242 -995 276
rect -877 242 -865 276
rect -1007 236 -865 242
rect -799 276 -657 282
rect -799 242 -787 276
rect -669 242 -657 276
rect -799 236 -657 242
rect -591 276 -449 282
rect -591 242 -579 276
rect -461 242 -449 276
rect -591 236 -449 242
rect -383 276 -241 282
rect -383 242 -371 276
rect -253 242 -241 276
rect -383 236 -241 242
rect -175 276 -33 282
rect -175 242 -163 276
rect -45 242 -33 276
rect -175 236 -33 242
rect 33 276 175 282
rect 33 242 45 276
rect 163 242 175 276
rect 33 236 175 242
rect 241 276 383 282
rect 241 242 253 276
rect 371 242 383 276
rect 241 236 383 242
rect 449 276 591 282
rect 449 242 461 276
rect 579 242 591 276
rect 449 236 591 242
rect 657 276 799 282
rect 657 242 669 276
rect 787 242 799 276
rect 657 236 799 242
rect 865 276 1007 282
rect 865 242 877 276
rect 995 242 1007 276
rect 865 236 1007 242
rect 1073 276 1215 282
rect 1073 242 1085 276
rect 1203 242 1215 276
rect 1073 236 1215 242
rect -1271 183 -1225 195
rect -1271 -183 -1265 183
rect -1231 -183 -1225 183
rect -1271 -195 -1225 -183
rect -1063 183 -1017 195
rect -1063 -183 -1057 183
rect -1023 -183 -1017 183
rect -1063 -195 -1017 -183
rect -855 183 -809 195
rect -855 -183 -849 183
rect -815 -183 -809 183
rect -855 -195 -809 -183
rect -647 183 -601 195
rect -647 -183 -641 183
rect -607 -183 -601 183
rect -647 -195 -601 -183
rect -439 183 -393 195
rect -439 -183 -433 183
rect -399 -183 -393 183
rect -439 -195 -393 -183
rect -231 183 -185 195
rect -231 -183 -225 183
rect -191 -183 -185 183
rect -231 -195 -185 -183
rect -23 183 23 195
rect -23 -183 -17 183
rect 17 -183 23 183
rect -23 -195 23 -183
rect 185 183 231 195
rect 185 -183 191 183
rect 225 -183 231 183
rect 185 -195 231 -183
rect 393 183 439 195
rect 393 -183 399 183
rect 433 -183 439 183
rect 393 -195 439 -183
rect 601 183 647 195
rect 601 -183 607 183
rect 641 -183 647 183
rect 601 -195 647 -183
rect 809 183 855 195
rect 809 -183 815 183
rect 849 -183 855 183
rect 809 -195 855 -183
rect 1017 183 1063 195
rect 1017 -183 1023 183
rect 1057 -183 1063 183
rect 1017 -195 1063 -183
rect 1225 183 1271 195
rect 1225 -183 1231 183
rect 1265 -183 1271 183
rect 1225 -195 1271 -183
rect -1215 -242 -1073 -236
rect -1215 -276 -1203 -242
rect -1085 -276 -1073 -242
rect -1215 -282 -1073 -276
rect -1007 -242 -865 -236
rect -1007 -276 -995 -242
rect -877 -276 -865 -242
rect -1007 -282 -865 -276
rect -799 -242 -657 -236
rect -799 -276 -787 -242
rect -669 -276 -657 -242
rect -799 -282 -657 -276
rect -591 -242 -449 -236
rect -591 -276 -579 -242
rect -461 -276 -449 -242
rect -591 -282 -449 -276
rect -383 -242 -241 -236
rect -383 -276 -371 -242
rect -253 -276 -241 -242
rect -383 -282 -241 -276
rect -175 -242 -33 -236
rect -175 -276 -163 -242
rect -45 -276 -33 -242
rect -175 -282 -33 -276
rect 33 -242 175 -236
rect 33 -276 45 -242
rect 163 -276 175 -242
rect 33 -282 175 -276
rect 241 -242 383 -236
rect 241 -276 253 -242
rect 371 -276 383 -242
rect 241 -282 383 -276
rect 449 -242 591 -236
rect 449 -276 461 -242
rect 579 -276 591 -242
rect 449 -282 591 -276
rect 657 -242 799 -236
rect 657 -276 669 -242
rect 787 -276 799 -242
rect 657 -282 799 -276
rect 865 -242 1007 -236
rect 865 -276 877 -242
rect 995 -276 1007 -242
rect 865 -282 1007 -276
rect 1073 -242 1215 -236
rect 1073 -276 1085 -242
rect 1203 -276 1215 -242
rect 1073 -282 1215 -276
<< properties >>
string FIXED_BBOX -1362 -361 1362 361
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.95 l 0.75 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
