magic
tech sky130A
magscale 1 2
timestamp 1770035380
<< error_p >>
rect -1214 512 -1156 518
rect -1056 512 -998 518
rect -898 512 -840 518
rect -740 512 -682 518
rect -582 512 -524 518
rect -424 512 -366 518
rect -266 512 -208 518
rect -108 512 -50 518
rect 50 512 108 518
rect 208 512 266 518
rect 366 512 424 518
rect 524 512 582 518
rect 682 512 740 518
rect 840 512 898 518
rect 998 512 1056 518
rect 1156 512 1214 518
rect -1214 478 -1202 512
rect -1056 478 -1044 512
rect -898 478 -886 512
rect -740 478 -728 512
rect -582 478 -570 512
rect -424 478 -412 512
rect -266 478 -254 512
rect -108 478 -96 512
rect 50 478 62 512
rect 208 478 220 512
rect 366 478 378 512
rect 524 478 536 512
rect 682 478 694 512
rect 840 478 852 512
rect 998 478 1010 512
rect 1156 478 1168 512
rect -1214 472 -1156 478
rect -1056 472 -998 478
rect -898 472 -840 478
rect -740 472 -682 478
rect -582 472 -524 478
rect -424 472 -366 478
rect -266 472 -208 478
rect -108 472 -50 478
rect 50 472 108 478
rect 208 472 266 478
rect 366 472 424 478
rect 524 472 582 478
rect 682 472 740 478
rect 840 472 898 478
rect 998 472 1056 478
rect 1156 472 1214 478
<< mvnmos >>
rect -1235 -502 -1135 440
rect -1077 -502 -977 440
rect -919 -502 -819 440
rect -761 -502 -661 440
rect -603 -502 -503 440
rect -445 -502 -345 440
rect -287 -502 -187 440
rect -129 -502 -29 440
rect 29 -502 129 440
rect 187 -502 287 440
rect 345 -502 445 440
rect 503 -502 603 440
rect 661 -502 761 440
rect 819 -502 919 440
rect 977 -502 1077 440
rect 1135 -502 1235 440
<< mvndiff >>
rect -1293 428 -1235 440
rect -1293 -490 -1281 428
rect -1247 -490 -1235 428
rect -1293 -502 -1235 -490
rect -1135 428 -1077 440
rect -1135 -490 -1123 428
rect -1089 -490 -1077 428
rect -1135 -502 -1077 -490
rect -977 428 -919 440
rect -977 -490 -965 428
rect -931 -490 -919 428
rect -977 -502 -919 -490
rect -819 428 -761 440
rect -819 -490 -807 428
rect -773 -490 -761 428
rect -819 -502 -761 -490
rect -661 428 -603 440
rect -661 -490 -649 428
rect -615 -490 -603 428
rect -661 -502 -603 -490
rect -503 428 -445 440
rect -503 -490 -491 428
rect -457 -490 -445 428
rect -503 -502 -445 -490
rect -345 428 -287 440
rect -345 -490 -333 428
rect -299 -490 -287 428
rect -345 -502 -287 -490
rect -187 428 -129 440
rect -187 -490 -175 428
rect -141 -490 -129 428
rect -187 -502 -129 -490
rect -29 428 29 440
rect -29 -490 -17 428
rect 17 -490 29 428
rect -29 -502 29 -490
rect 129 428 187 440
rect 129 -490 141 428
rect 175 -490 187 428
rect 129 -502 187 -490
rect 287 428 345 440
rect 287 -490 299 428
rect 333 -490 345 428
rect 287 -502 345 -490
rect 445 428 503 440
rect 445 -490 457 428
rect 491 -490 503 428
rect 445 -502 503 -490
rect 603 428 661 440
rect 603 -490 615 428
rect 649 -490 661 428
rect 603 -502 661 -490
rect 761 428 819 440
rect 761 -490 773 428
rect 807 -490 819 428
rect 761 -502 819 -490
rect 919 428 977 440
rect 919 -490 931 428
rect 965 -490 977 428
rect 919 -502 977 -490
rect 1077 428 1135 440
rect 1077 -490 1089 428
rect 1123 -490 1135 428
rect 1077 -502 1135 -490
rect 1235 428 1293 440
rect 1235 -490 1247 428
rect 1281 -490 1293 428
rect 1235 -502 1293 -490
<< mvndiffc >>
rect -1281 -490 -1247 428
rect -1123 -490 -1089 428
rect -965 -490 -931 428
rect -807 -490 -773 428
rect -649 -490 -615 428
rect -491 -490 -457 428
rect -333 -490 -299 428
rect -175 -490 -141 428
rect -17 -490 17 428
rect 141 -490 175 428
rect 299 -490 333 428
rect 457 -490 491 428
rect 615 -490 649 428
rect 773 -490 807 428
rect 931 -490 965 428
rect 1089 -490 1123 428
rect 1247 -490 1281 428
<< poly >>
rect -1218 512 -1152 528
rect -1218 495 -1202 512
rect -1235 478 -1202 495
rect -1168 495 -1152 512
rect -1060 512 -994 528
rect -1060 495 -1044 512
rect -1168 478 -1135 495
rect -1235 440 -1135 478
rect -1077 478 -1044 495
rect -1010 495 -994 512
rect -902 512 -836 528
rect -902 495 -886 512
rect -1010 478 -977 495
rect -1077 440 -977 478
rect -919 478 -886 495
rect -852 495 -836 512
rect -744 512 -678 528
rect -744 495 -728 512
rect -852 478 -819 495
rect -919 440 -819 478
rect -761 478 -728 495
rect -694 495 -678 512
rect -586 512 -520 528
rect -586 495 -570 512
rect -694 478 -661 495
rect -761 440 -661 478
rect -603 478 -570 495
rect -536 495 -520 512
rect -428 512 -362 528
rect -428 495 -412 512
rect -536 478 -503 495
rect -603 440 -503 478
rect -445 478 -412 495
rect -378 495 -362 512
rect -270 512 -204 528
rect -270 495 -254 512
rect -378 478 -345 495
rect -445 440 -345 478
rect -287 478 -254 495
rect -220 495 -204 512
rect -112 512 -46 528
rect -112 495 -96 512
rect -220 478 -187 495
rect -287 440 -187 478
rect -129 478 -96 495
rect -62 495 -46 512
rect 46 512 112 528
rect 46 495 62 512
rect -62 478 -29 495
rect -129 440 -29 478
rect 29 478 62 495
rect 96 495 112 512
rect 204 512 270 528
rect 204 495 220 512
rect 96 478 129 495
rect 29 440 129 478
rect 187 478 220 495
rect 254 495 270 512
rect 362 512 428 528
rect 362 495 378 512
rect 254 478 287 495
rect 187 440 287 478
rect 345 478 378 495
rect 412 495 428 512
rect 520 512 586 528
rect 520 495 536 512
rect 412 478 445 495
rect 345 440 445 478
rect 503 478 536 495
rect 570 495 586 512
rect 678 512 744 528
rect 678 495 694 512
rect 570 478 603 495
rect 503 440 603 478
rect 661 478 694 495
rect 728 495 744 512
rect 836 512 902 528
rect 836 495 852 512
rect 728 478 761 495
rect 661 440 761 478
rect 819 478 852 495
rect 886 495 902 512
rect 994 512 1060 528
rect 994 495 1010 512
rect 886 478 919 495
rect 819 440 919 478
rect 977 478 1010 495
rect 1044 495 1060 512
rect 1152 512 1218 528
rect 1152 495 1168 512
rect 1044 478 1077 495
rect 977 440 1077 478
rect 1135 478 1168 495
rect 1202 495 1218 512
rect 1202 478 1235 495
rect 1135 440 1235 478
rect -1235 -528 -1135 -502
rect -1077 -528 -977 -502
rect -919 -528 -819 -502
rect -761 -528 -661 -502
rect -603 -528 -503 -502
rect -445 -528 -345 -502
rect -287 -528 -187 -502
rect -129 -528 -29 -502
rect 29 -528 129 -502
rect 187 -528 287 -502
rect 345 -528 445 -502
rect 503 -528 603 -502
rect 661 -528 761 -502
rect 819 -528 919 -502
rect 977 -528 1077 -502
rect 1135 -528 1235 -502
<< polycont >>
rect -1202 478 -1168 512
rect -1044 478 -1010 512
rect -886 478 -852 512
rect -728 478 -694 512
rect -570 478 -536 512
rect -412 478 -378 512
rect -254 478 -220 512
rect -96 478 -62 512
rect 62 478 96 512
rect 220 478 254 512
rect 378 478 412 512
rect 536 478 570 512
rect 694 478 728 512
rect 852 478 886 512
rect 1010 478 1044 512
rect 1168 478 1202 512
<< locali >>
rect -1218 478 -1202 512
rect -1168 478 -1152 512
rect -1060 478 -1044 512
rect -1010 478 -994 512
rect -902 478 -886 512
rect -852 478 -836 512
rect -744 478 -728 512
rect -694 478 -678 512
rect -586 478 -570 512
rect -536 478 -520 512
rect -428 478 -412 512
rect -378 478 -362 512
rect -270 478 -254 512
rect -220 478 -204 512
rect -112 478 -96 512
rect -62 478 -46 512
rect 46 478 62 512
rect 96 478 112 512
rect 204 478 220 512
rect 254 478 270 512
rect 362 478 378 512
rect 412 478 428 512
rect 520 478 536 512
rect 570 478 586 512
rect 678 478 694 512
rect 728 478 744 512
rect 836 478 852 512
rect 886 478 902 512
rect 994 478 1010 512
rect 1044 478 1060 512
rect 1152 478 1168 512
rect 1202 478 1218 512
rect -1281 428 -1247 444
rect -1281 -506 -1247 -490
rect -1123 428 -1089 444
rect -1123 -506 -1089 -490
rect -965 428 -931 444
rect -965 -506 -931 -490
rect -807 428 -773 444
rect -807 -506 -773 -490
rect -649 428 -615 444
rect -649 -506 -615 -490
rect -491 428 -457 444
rect -491 -506 -457 -490
rect -333 428 -299 444
rect -333 -506 -299 -490
rect -175 428 -141 444
rect -175 -506 -141 -490
rect -17 428 17 444
rect -17 -506 17 -490
rect 141 428 175 444
rect 141 -506 175 -490
rect 299 428 333 444
rect 299 -506 333 -490
rect 457 428 491 444
rect 457 -506 491 -490
rect 615 428 649 444
rect 615 -506 649 -490
rect 773 428 807 444
rect 773 -506 807 -490
rect 931 428 965 444
rect 931 -506 965 -490
rect 1089 428 1123 444
rect 1089 -506 1123 -490
rect 1247 428 1281 444
rect 1247 -506 1281 -490
<< viali >>
rect -1202 478 -1168 512
rect -1044 478 -1010 512
rect -886 478 -852 512
rect -728 478 -694 512
rect -570 478 -536 512
rect -412 478 -378 512
rect -254 478 -220 512
rect -96 478 -62 512
rect 62 478 96 512
rect 220 478 254 512
rect 378 478 412 512
rect 536 478 570 512
rect 694 478 728 512
rect 852 478 886 512
rect 1010 478 1044 512
rect 1168 478 1202 512
rect -1281 -490 -1247 428
rect -1123 -490 -1089 428
rect -965 -490 -931 428
rect -807 -490 -773 428
rect -649 -490 -615 428
rect -491 -490 -457 428
rect -333 -490 -299 428
rect -175 -490 -141 428
rect -17 -490 17 428
rect 141 -490 175 428
rect 299 -490 333 428
rect 457 -490 491 428
rect 615 -490 649 428
rect 773 -490 807 428
rect 931 -490 965 428
rect 1089 -490 1123 428
rect 1247 -490 1281 428
<< metal1 >>
rect -1214 512 -1156 518
rect -1214 478 -1202 512
rect -1168 478 -1156 512
rect -1214 472 -1156 478
rect -1056 512 -998 518
rect -1056 478 -1044 512
rect -1010 478 -998 512
rect -1056 472 -998 478
rect -898 512 -840 518
rect -898 478 -886 512
rect -852 478 -840 512
rect -898 472 -840 478
rect -740 512 -682 518
rect -740 478 -728 512
rect -694 478 -682 512
rect -740 472 -682 478
rect -582 512 -524 518
rect -582 478 -570 512
rect -536 478 -524 512
rect -582 472 -524 478
rect -424 512 -366 518
rect -424 478 -412 512
rect -378 478 -366 512
rect -424 472 -366 478
rect -266 512 -208 518
rect -266 478 -254 512
rect -220 478 -208 512
rect -266 472 -208 478
rect -108 512 -50 518
rect -108 478 -96 512
rect -62 478 -50 512
rect -108 472 -50 478
rect 50 512 108 518
rect 50 478 62 512
rect 96 478 108 512
rect 50 472 108 478
rect 208 512 266 518
rect 208 478 220 512
rect 254 478 266 512
rect 208 472 266 478
rect 366 512 424 518
rect 366 478 378 512
rect 412 478 424 512
rect 366 472 424 478
rect 524 512 582 518
rect 524 478 536 512
rect 570 478 582 512
rect 524 472 582 478
rect 682 512 740 518
rect 682 478 694 512
rect 728 478 740 512
rect 682 472 740 478
rect 840 512 898 518
rect 840 478 852 512
rect 886 478 898 512
rect 840 472 898 478
rect 998 512 1056 518
rect 998 478 1010 512
rect 1044 478 1056 512
rect 998 472 1056 478
rect 1156 512 1214 518
rect 1156 478 1168 512
rect 1202 478 1214 512
rect 1156 472 1214 478
rect -1287 428 -1241 440
rect -1287 -490 -1281 428
rect -1247 -490 -1241 428
rect -1287 -502 -1241 -490
rect -1129 428 -1083 440
rect -1129 -490 -1123 428
rect -1089 -490 -1083 428
rect -1129 -502 -1083 -490
rect -971 428 -925 440
rect -971 -490 -965 428
rect -931 -490 -925 428
rect -971 -502 -925 -490
rect -813 428 -767 440
rect -813 -490 -807 428
rect -773 -490 -767 428
rect -813 -502 -767 -490
rect -655 428 -609 440
rect -655 -490 -649 428
rect -615 -490 -609 428
rect -655 -502 -609 -490
rect -497 428 -451 440
rect -497 -490 -491 428
rect -457 -490 -451 428
rect -497 -502 -451 -490
rect -339 428 -293 440
rect -339 -490 -333 428
rect -299 -490 -293 428
rect -339 -502 -293 -490
rect -181 428 -135 440
rect -181 -490 -175 428
rect -141 -490 -135 428
rect -181 -502 -135 -490
rect -23 428 23 440
rect -23 -490 -17 428
rect 17 200 23 428
rect 135 428 181 440
rect 135 200 141 428
rect 17 0 141 200
rect 17 -200 23 0
rect 135 -200 141 0
rect 17 -400 141 -200
rect 17 -490 23 -400
rect -23 -502 23 -490
rect 135 -490 141 -400
rect 175 200 181 428
rect 293 428 339 440
rect 175 0 200 200
rect 175 -200 181 0
rect 175 -400 200 -200
rect 175 -490 181 -400
rect 135 -502 181 -490
rect 293 -490 299 428
rect 333 -490 339 428
rect 293 -502 339 -490
rect 451 428 497 440
rect 451 -490 457 428
rect 491 -490 497 428
rect 451 -502 497 -490
rect 609 428 655 440
rect 609 -490 615 428
rect 649 -490 655 428
rect 609 -502 655 -490
rect 767 428 813 440
rect 767 -490 773 428
rect 807 -490 813 428
rect 767 -502 813 -490
rect 925 428 971 440
rect 925 -490 931 428
rect 965 -490 971 428
rect 925 -502 971 -490
rect 1083 428 1129 440
rect 1083 -490 1089 428
rect 1123 -490 1129 428
rect 1083 -502 1129 -490
rect 1241 428 1287 440
rect 1241 -490 1247 428
rect 1281 -490 1287 428
rect 1241 -502 1287 -490
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
rect 0 -8800 200 -8600
rect 0 -9200 200 -9000
rect 0 -9600 200 -9400
rect 0 -10000 200 -9800
rect 0 -10400 200 -10200
rect 0 -10800 200 -10600
rect 0 -11200 200 -11000
rect 0 -11600 200 -11400
rect 0 -12000 200 -11800
rect 0 -12400 200 -12200
rect 0 -12800 200 -12600
rect 0 -13200 200 -13000
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X0
timestamp 0
transform 1 0 -1080 0 1 -12536
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X1
timestamp 0
transform 1 0 -589 0 1 -12601
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X2
timestamp 0
transform 1 0 -98 0 1 -12666
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X3
timestamp 0
transform 1 0 393 0 1 -12731
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X4
timestamp 0
transform 1 0 884 0 1 -12796
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X5
timestamp 0
transform 1 0 1375 0 1 -12861
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X6
timestamp 0
transform 1 0 1866 0 1 -12926
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X7
timestamp 0
transform 1 0 2357 0 1 -12991
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X8
timestamp 0
transform 1 0 2848 0 1 -13056
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_CJYKFD  X9
timestamp 0
transform 1 0 3339 0 1 -13121
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_JAZF34  X10
timestamp 0
transform 1 0 3830 0 1 -13186
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X11
timestamp 0
transform 1 0 4321 0 1 -13251
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X12
timestamp 0
transform 1 0 4812 0 1 -13316
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X13
timestamp 0
transform 1 0 5303 0 1 -13381
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X14
timestamp 0
transform 1 0 5794 0 1 -13446
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_HGUXL5  X15
timestamp 0
transform 1 0 6285 0 1 -13511
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 a_n819_n502#
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 a_n1135_n502#
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 a_129_n502#
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 {}
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 a_n503_n502#
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 a_n1293_n502#
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 a_29_n528#
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 a_n129_n528#
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 a_n661_n502#
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 a_187_n528#
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 a_819_n528#
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 a_n287_n528#
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 a_n1077_n528#
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 a_445_n502#
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 a_345_n528#
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 a_n919_n528#
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 a_977_n528#
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 a_n445_n528#
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 {}
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 a_1077_n502#
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 256 0 0 0 a_n1235_n528#
port 21 nsew
flabel metal1 0 -8800 200 -8600 0 FreeSans 256 0 0 0 a_603_n502#
port 22 nsew
flabel metal1 0 -9200 200 -9000 0 FreeSans 256 0 0 0 a_503_n528#
port 23 nsew
flabel metal1 0 -9600 200 -9400 0 FreeSans 256 0 0 0 a_n603_n528#
port 24 nsew
flabel metal1 0 -10000 200 -9800 0 FreeSans 256 0 0 0 a_1235_n502#
port 25 nsew
flabel metal1 0 -10400 200 -10200 0 FreeSans 256 0 0 0 a_1135_n528#
port 26 nsew
flabel metal1 0 -10800 200 -10600 0 FreeSans 256 0 0 0 {}
port 27 nsew
flabel metal1 0 -11200 200 -11000 0 FreeSans 256 0 0 0 a_661_n528#
port 28 nsew
flabel metal1 0 -11600 200 -11400 0 FreeSans 256 0 0 0 a_761_n502#
port 29 nsew
flabel metal1 0 -12000 200 -11800 0 FreeSans 256 0 0 0 a_n29_n502#
port 30 nsew
flabel metal1 0 -12400 200 -12200 0 FreeSans 256 0 0 0 a_n761_n528#
port 31 nsew
flabel metal1 0 -12800 200 -12600 0 FreeSans 256 0 0 0 a_n187_n502#
port 32 nsew
flabel metal1 0 -13200 200 -13000 0 FreeSans 256 0 0 0 VSUBS
port 33 nsew
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.7125 l 0.5 m 1 nf 16 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
