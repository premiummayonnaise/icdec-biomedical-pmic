magic
tech sky130A
magscale 1 2
timestamp 1769411983
<< error_p >>
rect -2559 1098 2559 1102
rect -2559 -1030 -2529 1098
rect -2493 1032 2493 1036
rect -2493 -964 -2463 1032
rect 2463 -964 2493 1032
rect 2529 -1030 2559 1098
<< nwell >>
rect -2529 -1064 2529 1098
<< mvpmos >>
rect -2435 -964 -2185 1036
rect -2127 -964 -1877 1036
rect -1819 -964 -1569 1036
rect -1511 -964 -1261 1036
rect -1203 -964 -953 1036
rect -895 -964 -645 1036
rect -587 -964 -337 1036
rect -279 -964 -29 1036
rect 29 -964 279 1036
rect 337 -964 587 1036
rect 645 -964 895 1036
rect 953 -964 1203 1036
rect 1261 -964 1511 1036
rect 1569 -964 1819 1036
rect 1877 -964 2127 1036
rect 2185 -964 2435 1036
<< mvpdiff >>
rect -2493 1024 -2435 1036
rect -2493 -952 -2481 1024
rect -2447 -952 -2435 1024
rect -2493 -964 -2435 -952
rect -2185 1024 -2127 1036
rect -2185 -952 -2173 1024
rect -2139 -952 -2127 1024
rect -2185 -964 -2127 -952
rect -1877 1024 -1819 1036
rect -1877 -952 -1865 1024
rect -1831 -952 -1819 1024
rect -1877 -964 -1819 -952
rect -1569 1024 -1511 1036
rect -1569 -952 -1557 1024
rect -1523 -952 -1511 1024
rect -1569 -964 -1511 -952
rect -1261 1024 -1203 1036
rect -1261 -952 -1249 1024
rect -1215 -952 -1203 1024
rect -1261 -964 -1203 -952
rect -953 1024 -895 1036
rect -953 -952 -941 1024
rect -907 -952 -895 1024
rect -953 -964 -895 -952
rect -645 1024 -587 1036
rect -645 -952 -633 1024
rect -599 -952 -587 1024
rect -645 -964 -587 -952
rect -337 1024 -279 1036
rect -337 -952 -325 1024
rect -291 -952 -279 1024
rect -337 -964 -279 -952
rect -29 1024 29 1036
rect -29 -952 -17 1024
rect 17 -952 29 1024
rect -29 -964 29 -952
rect 279 1024 337 1036
rect 279 -952 291 1024
rect 325 -952 337 1024
rect 279 -964 337 -952
rect 587 1024 645 1036
rect 587 -952 599 1024
rect 633 -952 645 1024
rect 587 -964 645 -952
rect 895 1024 953 1036
rect 895 -952 907 1024
rect 941 -952 953 1024
rect 895 -964 953 -952
rect 1203 1024 1261 1036
rect 1203 -952 1215 1024
rect 1249 -952 1261 1024
rect 1203 -964 1261 -952
rect 1511 1024 1569 1036
rect 1511 -952 1523 1024
rect 1557 -952 1569 1024
rect 1511 -964 1569 -952
rect 1819 1024 1877 1036
rect 1819 -952 1831 1024
rect 1865 -952 1877 1024
rect 1819 -964 1877 -952
rect 2127 1024 2185 1036
rect 2127 -952 2139 1024
rect 2173 -952 2185 1024
rect 2127 -964 2185 -952
rect 2435 1024 2493 1036
rect 2435 -952 2447 1024
rect 2481 -952 2493 1024
rect 2435 -964 2493 -952
<< mvpdiffc >>
rect -2481 -952 -2447 1024
rect -2173 -952 -2139 1024
rect -1865 -952 -1831 1024
rect -1557 -952 -1523 1024
rect -1249 -952 -1215 1024
rect -941 -952 -907 1024
rect -633 -952 -599 1024
rect -325 -952 -291 1024
rect -17 -952 17 1024
rect 291 -952 325 1024
rect 599 -952 633 1024
rect 907 -952 941 1024
rect 1215 -952 1249 1024
rect 1523 -952 1557 1024
rect 1831 -952 1865 1024
rect 2139 -952 2173 1024
rect 2447 -952 2481 1024
<< poly >>
rect -2435 1036 -2185 1062
rect -2127 1036 -1877 1062
rect -1819 1036 -1569 1062
rect -1511 1036 -1261 1062
rect -1203 1036 -953 1062
rect -895 1036 -645 1062
rect -587 1036 -337 1062
rect -279 1036 -29 1062
rect 29 1036 279 1062
rect 337 1036 587 1062
rect 645 1036 895 1062
rect 953 1036 1203 1062
rect 1261 1036 1511 1062
rect 1569 1036 1819 1062
rect 1877 1036 2127 1062
rect 2185 1036 2435 1062
rect -2435 -1011 -2185 -964
rect -2435 -1045 -2419 -1011
rect -2201 -1045 -2185 -1011
rect -2435 -1061 -2185 -1045
rect -2127 -1011 -1877 -964
rect -2127 -1045 -2111 -1011
rect -1893 -1045 -1877 -1011
rect -2127 -1061 -1877 -1045
rect -1819 -1011 -1569 -964
rect -1819 -1045 -1803 -1011
rect -1585 -1045 -1569 -1011
rect -1819 -1061 -1569 -1045
rect -1511 -1011 -1261 -964
rect -1511 -1045 -1495 -1011
rect -1277 -1045 -1261 -1011
rect -1511 -1061 -1261 -1045
rect -1203 -1011 -953 -964
rect -1203 -1045 -1187 -1011
rect -969 -1045 -953 -1011
rect -1203 -1061 -953 -1045
rect -895 -1011 -645 -964
rect -895 -1045 -879 -1011
rect -661 -1045 -645 -1011
rect -895 -1061 -645 -1045
rect -587 -1011 -337 -964
rect -587 -1045 -571 -1011
rect -353 -1045 -337 -1011
rect -587 -1061 -337 -1045
rect -279 -1011 -29 -964
rect -279 -1045 -263 -1011
rect -45 -1045 -29 -1011
rect -279 -1061 -29 -1045
rect 29 -1011 279 -964
rect 29 -1045 45 -1011
rect 263 -1045 279 -1011
rect 29 -1061 279 -1045
rect 337 -1011 587 -964
rect 337 -1045 353 -1011
rect 571 -1045 587 -1011
rect 337 -1061 587 -1045
rect 645 -1011 895 -964
rect 645 -1045 661 -1011
rect 879 -1045 895 -1011
rect 645 -1061 895 -1045
rect 953 -1011 1203 -964
rect 953 -1045 969 -1011
rect 1187 -1045 1203 -1011
rect 953 -1061 1203 -1045
rect 1261 -1011 1511 -964
rect 1261 -1045 1277 -1011
rect 1495 -1045 1511 -1011
rect 1261 -1061 1511 -1045
rect 1569 -1011 1819 -964
rect 1569 -1045 1585 -1011
rect 1803 -1045 1819 -1011
rect 1569 -1061 1819 -1045
rect 1877 -1011 2127 -964
rect 1877 -1045 1893 -1011
rect 2111 -1045 2127 -1011
rect 1877 -1061 2127 -1045
rect 2185 -1011 2435 -964
rect 2185 -1045 2201 -1011
rect 2419 -1045 2435 -1011
rect 2185 -1061 2435 -1045
<< polycont >>
rect -2419 -1045 -2201 -1011
rect -2111 -1045 -1893 -1011
rect -1803 -1045 -1585 -1011
rect -1495 -1045 -1277 -1011
rect -1187 -1045 -969 -1011
rect -879 -1045 -661 -1011
rect -571 -1045 -353 -1011
rect -263 -1045 -45 -1011
rect 45 -1045 263 -1011
rect 353 -1045 571 -1011
rect 661 -1045 879 -1011
rect 969 -1045 1187 -1011
rect 1277 -1045 1495 -1011
rect 1585 -1045 1803 -1011
rect 1893 -1045 2111 -1011
rect 2201 -1045 2419 -1011
<< locali >>
rect -2481 1024 -2447 1040
rect -2481 -968 -2447 -952
rect -2173 1024 -2139 1040
rect -2173 -968 -2139 -952
rect -1865 1024 -1831 1040
rect -1865 -968 -1831 -952
rect -1557 1024 -1523 1040
rect -1557 -968 -1523 -952
rect -1249 1024 -1215 1040
rect -1249 -968 -1215 -952
rect -941 1024 -907 1040
rect -941 -968 -907 -952
rect -633 1024 -599 1040
rect -633 -968 -599 -952
rect -325 1024 -291 1040
rect -325 -968 -291 -952
rect -17 1024 17 1040
rect -17 -968 17 -952
rect 291 1024 325 1040
rect 291 -968 325 -952
rect 599 1024 633 1040
rect 599 -968 633 -952
rect 907 1024 941 1040
rect 907 -968 941 -952
rect 1215 1024 1249 1040
rect 1215 -968 1249 -952
rect 1523 1024 1557 1040
rect 1523 -968 1557 -952
rect 1831 1024 1865 1040
rect 1831 -968 1865 -952
rect 2139 1024 2173 1040
rect 2139 -968 2173 -952
rect 2447 1024 2481 1040
rect 2447 -968 2481 -952
rect -2435 -1045 -2419 -1011
rect -2201 -1045 -2185 -1011
rect -2127 -1045 -2111 -1011
rect -1893 -1045 -1877 -1011
rect -1819 -1045 -1803 -1011
rect -1585 -1045 -1569 -1011
rect -1511 -1045 -1495 -1011
rect -1277 -1045 -1261 -1011
rect -1203 -1045 -1187 -1011
rect -969 -1045 -953 -1011
rect -895 -1045 -879 -1011
rect -661 -1045 -645 -1011
rect -587 -1045 -571 -1011
rect -353 -1045 -337 -1011
rect -279 -1045 -263 -1011
rect -45 -1045 -29 -1011
rect 29 -1045 45 -1011
rect 263 -1045 279 -1011
rect 337 -1045 353 -1011
rect 571 -1045 587 -1011
rect 645 -1045 661 -1011
rect 879 -1045 895 -1011
rect 953 -1045 969 -1011
rect 1187 -1045 1203 -1011
rect 1261 -1045 1277 -1011
rect 1495 -1045 1511 -1011
rect 1569 -1045 1585 -1011
rect 1803 -1045 1819 -1011
rect 1877 -1045 1893 -1011
rect 2111 -1045 2127 -1011
rect 2185 -1045 2201 -1011
rect 2419 -1045 2435 -1011
<< viali >>
rect -2481 -952 -2447 1024
rect -2173 -952 -2139 1024
rect -1865 -952 -1831 1024
rect -1557 -952 -1523 1024
rect -1249 -952 -1215 1024
rect -941 -952 -907 1024
rect -633 -952 -599 1024
rect -325 -952 -291 1024
rect -17 -952 17 1024
rect 291 -952 325 1024
rect 599 -952 633 1024
rect 907 -952 941 1024
rect 1215 -952 1249 1024
rect 1523 -952 1557 1024
rect 1831 -952 1865 1024
rect 2139 -952 2173 1024
rect 2447 -952 2481 1024
rect -2419 -1045 -2201 -1011
rect -2111 -1045 -1893 -1011
rect -1803 -1045 -1585 -1011
rect -1495 -1045 -1277 -1011
rect -1187 -1045 -969 -1011
rect -879 -1045 -661 -1011
rect -571 -1045 -353 -1011
rect -263 -1045 -45 -1011
rect 45 -1045 263 -1011
rect 353 -1045 571 -1011
rect 661 -1045 879 -1011
rect 969 -1045 1187 -1011
rect 1277 -1045 1495 -1011
rect 1585 -1045 1803 -1011
rect 1893 -1045 2111 -1011
rect 2201 -1045 2419 -1011
<< metal1 >>
rect -2487 1024 -2441 1036
rect -2487 -952 -2481 1024
rect -2447 -952 -2441 1024
rect -2487 -964 -2441 -952
rect -2179 1024 -2133 1036
rect -2179 -952 -2173 1024
rect -2139 -952 -2133 1024
rect -2179 -964 -2133 -952
rect -1871 1024 -1825 1036
rect -1871 -952 -1865 1024
rect -1831 -952 -1825 1024
rect -1871 -964 -1825 -952
rect -1563 1024 -1517 1036
rect -1563 -952 -1557 1024
rect -1523 -952 -1517 1024
rect -1563 -964 -1517 -952
rect -1255 1024 -1209 1036
rect -1255 -952 -1249 1024
rect -1215 -952 -1209 1024
rect -1255 -964 -1209 -952
rect -947 1024 -901 1036
rect -947 -952 -941 1024
rect -907 -952 -901 1024
rect -947 -964 -901 -952
rect -639 1024 -593 1036
rect -639 -952 -633 1024
rect -599 -952 -593 1024
rect -639 -964 -593 -952
rect -331 1024 -285 1036
rect -331 -952 -325 1024
rect -291 -952 -285 1024
rect -331 -964 -285 -952
rect -23 1024 23 1036
rect -23 -952 -17 1024
rect 17 -952 23 1024
rect -23 -964 23 -952
rect 285 1024 331 1036
rect 285 -952 291 1024
rect 325 -952 331 1024
rect 285 -964 331 -952
rect 593 1024 639 1036
rect 593 -952 599 1024
rect 633 -952 639 1024
rect 593 -964 639 -952
rect 901 1024 947 1036
rect 901 -952 907 1024
rect 941 -952 947 1024
rect 901 -964 947 -952
rect 1209 1024 1255 1036
rect 1209 -952 1215 1024
rect 1249 -952 1255 1024
rect 1209 -964 1255 -952
rect 1517 1024 1563 1036
rect 1517 -952 1523 1024
rect 1557 -952 1563 1024
rect 1517 -964 1563 -952
rect 1825 1024 1871 1036
rect 1825 -952 1831 1024
rect 1865 -952 1871 1024
rect 1825 -964 1871 -952
rect 2133 1024 2179 1036
rect 2133 -952 2139 1024
rect 2173 -952 2179 1024
rect 2133 -964 2179 -952
rect 2441 1024 2487 1036
rect 2441 -952 2447 1024
rect 2481 -952 2487 1024
rect 2441 -964 2487 -952
rect -2431 -1011 -2189 -1005
rect -2431 -1045 -2419 -1011
rect -2201 -1045 -2189 -1011
rect -2431 -1051 -2189 -1045
rect -2123 -1011 -1881 -1005
rect -2123 -1045 -2111 -1011
rect -1893 -1045 -1881 -1011
rect -2123 -1051 -1881 -1045
rect -1815 -1011 -1573 -1005
rect -1815 -1045 -1803 -1011
rect -1585 -1045 -1573 -1011
rect -1815 -1051 -1573 -1045
rect -1507 -1011 -1265 -1005
rect -1507 -1045 -1495 -1011
rect -1277 -1045 -1265 -1011
rect -1507 -1051 -1265 -1045
rect -1199 -1011 -957 -1005
rect -1199 -1045 -1187 -1011
rect -969 -1045 -957 -1011
rect -1199 -1051 -957 -1045
rect -891 -1011 -649 -1005
rect -891 -1045 -879 -1011
rect -661 -1045 -649 -1011
rect -891 -1051 -649 -1045
rect -583 -1011 -341 -1005
rect -583 -1045 -571 -1011
rect -353 -1045 -341 -1011
rect -583 -1051 -341 -1045
rect -275 -1011 -33 -1005
rect -275 -1045 -263 -1011
rect -45 -1045 -33 -1011
rect -275 -1051 -33 -1045
rect 33 -1011 275 -1005
rect 33 -1045 45 -1011
rect 263 -1045 275 -1011
rect 33 -1051 275 -1045
rect 341 -1011 583 -1005
rect 341 -1045 353 -1011
rect 571 -1045 583 -1011
rect 341 -1051 583 -1045
rect 649 -1011 891 -1005
rect 649 -1045 661 -1011
rect 879 -1045 891 -1011
rect 649 -1051 891 -1045
rect 957 -1011 1199 -1005
rect 957 -1045 969 -1011
rect 1187 -1045 1199 -1011
rect 957 -1051 1199 -1045
rect 1265 -1011 1507 -1005
rect 1265 -1045 1277 -1011
rect 1495 -1045 1507 -1011
rect 1265 -1051 1507 -1045
rect 1573 -1011 1815 -1005
rect 1573 -1045 1585 -1011
rect 1803 -1045 1815 -1011
rect 1573 -1051 1815 -1045
rect 1881 -1011 2123 -1005
rect 1881 -1045 1893 -1011
rect 2111 -1045 2123 -1011
rect 1881 -1051 2123 -1045
rect 2189 -1011 2431 -1005
rect 2189 -1045 2201 -1011
rect 2419 -1045 2431 -1011
rect 2189 -1051 2431 -1045
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 1.25 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
