magic
tech sky130A
magscale 1 2
timestamp 1769397192
<< metal3 >>
rect -2186 8492 2186 8520
rect -2186 4468 2102 8492
rect 2166 4468 2186 8492
rect -2186 4440 2186 4468
rect -2186 4172 2186 4200
rect -2186 148 2102 4172
rect 2166 148 2186 4172
rect -2186 120 2186 148
rect -2186 -148 2186 -120
rect -2186 -4172 2102 -148
rect 2166 -4172 2186 -148
rect -2186 -4200 2186 -4172
rect -2186 -4468 2186 -4440
rect -2186 -8492 2102 -4468
rect 2166 -8492 2186 -4468
rect -2186 -8520 2186 -8492
<< via3 >>
rect 2102 4468 2166 8492
rect 2102 148 2166 4172
rect 2102 -4172 2166 -148
rect 2102 -8492 2166 -4468
<< mimcap >>
rect -2146 8440 1854 8480
rect -2146 4520 -2106 8440
rect 1814 4520 1854 8440
rect -2146 4480 1854 4520
rect -2146 4120 1854 4160
rect -2146 200 -2106 4120
rect 1814 200 1854 4120
rect -2146 160 1854 200
rect -2146 -200 1854 -160
rect -2146 -4120 -2106 -200
rect 1814 -4120 1854 -200
rect -2146 -4160 1854 -4120
rect -2146 -4520 1854 -4480
rect -2146 -8440 -2106 -4520
rect 1814 -8440 1854 -4520
rect -2146 -8480 1854 -8440
<< mimcapcontact >>
rect -2106 4520 1814 8440
rect -2106 200 1814 4120
rect -2106 -4120 1814 -200
rect -2106 -8440 1814 -4520
<< metal4 >>
rect -198 8441 -94 8640
rect 2082 8492 2186 8640
rect -2107 8440 1815 8441
rect -2107 4520 -2106 8440
rect 1814 4520 1815 8440
rect -2107 4519 1815 4520
rect -198 4121 -94 4519
rect 2082 4468 2102 8492
rect 2166 4468 2186 8492
rect 2082 4172 2186 4468
rect -2107 4120 1815 4121
rect -2107 200 -2106 4120
rect 1814 200 1815 4120
rect -2107 199 1815 200
rect -198 -199 -94 199
rect 2082 148 2102 4172
rect 2166 148 2186 4172
rect 2082 -148 2186 148
rect -2107 -200 1815 -199
rect -2107 -4120 -2106 -200
rect 1814 -4120 1815 -200
rect -2107 -4121 1815 -4120
rect -198 -4519 -94 -4121
rect 2082 -4172 2102 -148
rect 2166 -4172 2186 -148
rect 2082 -4468 2186 -4172
rect -2107 -4520 1815 -4519
rect -2107 -8440 -2106 -4520
rect 1814 -8440 1815 -4520
rect -2107 -8441 1815 -8440
rect -198 -8640 -94 -8441
rect 2082 -8492 2102 -4468
rect 2166 -8492 2186 -4468
rect 2082 -8640 2186 -8492
<< properties >>
string FIXED_BBOX -2186 4440 1894 8520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20.0 l 20.0 val 815.2 carea 2.00 cperi 0.19 class capacitor nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
