magic
tech sky130A
magscale 1 2
timestamp 1769952370
<< mvnmos >>
rect -287 -501 -187 439
rect -129 -501 -29 439
rect 29 -501 129 439
rect 187 -501 287 439
<< mvndiff >>
rect -345 427 -287 439
rect -345 -489 -333 427
rect -299 -489 -287 427
rect -345 -501 -287 -489
rect -187 427 -129 439
rect -187 -489 -175 427
rect -141 -489 -129 427
rect -187 -501 -129 -489
rect -29 427 29 439
rect -29 -489 -17 427
rect 17 -489 29 427
rect -29 -501 29 -489
rect 129 427 187 439
rect 129 -489 141 427
rect 175 -489 187 427
rect 129 -501 187 -489
rect 287 427 345 439
rect 287 -489 299 427
rect 333 -489 345 427
rect 287 -501 345 -489
<< mvndiffc >>
rect -333 -489 -299 427
rect -175 -489 -141 427
rect -17 -489 17 427
rect 141 -489 175 427
rect 299 -489 333 427
<< poly >>
rect -287 511 -187 527
rect -287 477 -271 511
rect -203 477 -187 511
rect -287 439 -187 477
rect -129 511 -29 527
rect -129 477 -113 511
rect -45 477 -29 511
rect -129 439 -29 477
rect 29 511 129 527
rect 29 477 45 511
rect 113 477 129 511
rect 29 439 129 477
rect 187 511 287 527
rect 187 477 203 511
rect 271 477 287 511
rect 187 439 287 477
rect -287 -527 -187 -501
rect -129 -527 -29 -501
rect 29 -527 129 -501
rect 187 -527 287 -501
<< polycont >>
rect -271 477 -203 511
rect -113 477 -45 511
rect 45 477 113 511
rect 203 477 271 511
<< locali >>
rect -287 477 -271 511
rect -203 477 -187 511
rect -129 477 -113 511
rect -45 477 -29 511
rect 29 477 45 511
rect 113 477 129 511
rect 187 477 203 511
rect 271 477 287 511
rect -333 427 -299 443
rect -333 -505 -299 -489
rect -175 427 -141 443
rect -175 -505 -141 -489
rect -17 427 17 443
rect -17 -505 17 -489
rect 141 427 175 443
rect 141 -505 175 -489
rect 299 427 333 443
rect 299 -505 333 -489
<< viali >>
rect -271 477 -203 511
rect -113 477 -45 511
rect 45 477 113 511
rect 203 477 271 511
rect -333 -489 -299 427
rect -175 -489 -141 427
rect -17 -489 17 427
rect 141 -489 175 427
rect 299 -489 333 427
<< metal1 >>
rect -283 511 -191 517
rect -283 477 -271 511
rect -203 477 -191 511
rect -283 471 -191 477
rect -125 511 -33 517
rect -125 477 -113 511
rect -45 477 -33 511
rect -125 471 -33 477
rect 33 511 125 517
rect 33 477 45 511
rect 113 477 125 511
rect 33 471 125 477
rect 191 511 283 517
rect 191 477 203 511
rect 271 477 283 511
rect 191 471 283 477
rect -339 427 -293 439
rect -339 -489 -333 427
rect -299 -489 -293 427
rect -339 -501 -293 -489
rect -181 427 -135 439
rect -181 -489 -175 427
rect -141 -489 -135 427
rect -181 -501 -135 -489
rect -23 427 23 439
rect -23 -489 -17 427
rect 17 -489 23 427
rect -23 -501 23 -489
rect 135 427 181 439
rect 135 -489 141 427
rect 175 -489 181 427
rect 135 -501 181 -489
rect 293 427 339 439
rect 293 -489 299 427
rect 333 -489 339 427
rect 293 -501 339 -489
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.7 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
