magic
tech sky130A
magscale 1 2
timestamp 1769075133
<< pwell >>
rect -407 -558 407 558
<< mvnmos >>
rect -179 -300 -29 300
rect 29 -300 179 300
<< mvndiff >>
rect -237 288 -179 300
rect -237 -288 -225 288
rect -191 -288 -179 288
rect -237 -300 -179 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 179 288 237 300
rect 179 -288 191 288
rect 225 -288 237 288
rect 179 -300 237 -288
<< mvndiffc >>
rect -225 -288 -191 288
rect -17 -288 17 288
rect 191 -288 225 288
<< mvpsubdiff >>
rect -371 510 371 522
rect -371 476 -263 510
rect 263 476 371 510
rect -371 464 371 476
rect -371 414 -313 464
rect -371 -414 -359 414
rect -325 -414 -313 414
rect 313 414 371 464
rect -371 -464 -313 -414
rect 313 -414 325 414
rect 359 -414 371 414
rect 313 -464 371 -414
rect -371 -476 371 -464
rect -371 -510 -263 -476
rect 263 -510 371 -476
rect -371 -522 371 -510
<< mvpsubdiffcont >>
rect -263 476 263 510
rect -359 -414 -325 414
rect 325 -414 359 414
rect -263 -510 263 -476
<< poly >>
rect -179 372 -29 388
rect -179 338 -163 372
rect -45 338 -29 372
rect -179 300 -29 338
rect 29 372 179 388
rect 29 338 45 372
rect 163 338 179 372
rect 29 300 179 338
rect -179 -338 -29 -300
rect -179 -372 -163 -338
rect -45 -372 -29 -338
rect -179 -388 -29 -372
rect 29 -338 179 -300
rect 29 -372 45 -338
rect 163 -372 179 -338
rect 29 -388 179 -372
<< polycont >>
rect -163 338 -45 372
rect 45 338 163 372
rect -163 -372 -45 -338
rect 45 -372 163 -338
<< locali >>
rect -359 476 -263 510
rect 263 476 359 510
rect -359 414 -325 476
rect 325 414 359 476
rect -179 338 -163 372
rect -45 338 -29 372
rect 29 338 45 372
rect 163 338 179 372
rect -225 288 -191 304
rect -225 -304 -191 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 191 288 225 304
rect 191 -304 225 -288
rect -179 -372 -163 -338
rect -45 -372 -29 -338
rect 29 -372 45 -338
rect 163 -372 179 -338
rect -359 -476 -325 -414
rect 325 -476 359 -414
rect -359 -510 -263 -476
rect 263 -510 359 -476
<< viali >>
rect -163 338 -45 372
rect 45 338 163 372
rect -225 -288 -191 288
rect -17 -288 17 288
rect 191 -288 225 288
rect -163 -372 -45 -338
rect 45 -372 163 -338
<< metal1 >>
rect -175 372 -33 378
rect -175 338 -163 372
rect -45 338 -33 372
rect -175 332 -33 338
rect 33 372 175 378
rect 33 338 45 372
rect 163 338 175 372
rect 33 332 175 338
rect -231 288 -185 300
rect -231 -288 -225 288
rect -191 -288 -185 288
rect -231 -300 -185 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 185 288 231 300
rect 185 -288 191 288
rect 225 -288 231 288
rect 185 -300 231 -288
rect -175 -338 -33 -332
rect -175 -372 -163 -338
rect -45 -372 -33 -338
rect -175 -378 -33 -372
rect 33 -338 175 -332
rect 33 -372 45 -338
rect 163 -372 175 -338
rect 33 -378 175 -372
<< properties >>
string FIXED_BBOX -342 -493 342 493
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 0.75 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
