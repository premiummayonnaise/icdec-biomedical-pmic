magic
tech sky130A
magscale 1 2
timestamp 1769616064
<< error_s >>
rect 3956 -50 3980 -46
<< nwell >>
rect 2540 -180 4220 -120
<< pwell >>
rect 2540 -2660 4220 -180
<< locali >>
rect 2540 760 4220 1020
rect 2740 120 2790 650
rect 3050 160 3100 760
rect 3660 160 3710 760
rect 3980 120 4030 650
rect 2740 70 4030 120
rect 2600 -2390 2660 -340
rect 2740 -990 2790 70
rect 3980 -50 4030 70
rect 3940 -80 4030 -50
rect 3940 -990 3990 -80
rect 2730 -1040 3990 -990
rect 2730 -1720 2790 -1210
rect 3280 -1640 3330 -1040
rect 3400 -1640 3450 -1040
rect 3280 -1710 3460 -1690
rect 3280 -1720 3290 -1710
rect 2730 -1750 3290 -1720
rect 3330 -1750 3410 -1710
rect 3450 -1720 3460 -1710
rect 3940 -1720 4000 -1210
rect 3450 -1750 4000 -1720
rect 2730 -1770 4000 -1750
rect 2890 -1910 3860 -1850
rect 2740 -2390 2800 -1970
rect 3060 -2290 3110 -1910
rect 3940 -2390 4000 -1960
rect 4060 -2390 4120 -320
rect 2600 -2400 4120 -2390
rect 2540 -2660 4220 -2400
<< viali >>
rect 3290 -1750 3330 -1710
rect 3410 -1750 3450 -1710
<< metal1 >>
rect 2540 760 4220 1020
rect 0 -400 200 -200
rect 3330 -400 3420 650
rect 0 -800 200 -600
rect 2840 -980 2910 -860
rect 0 -1200 200 -1000
rect 2840 -1180 2910 -1060
rect 0 -1600 200 -1400
rect 2980 -1820 3090 -410
rect 3170 -910 3240 -850
rect 3310 -1080 3420 -400
rect 3500 -910 3570 -850
rect 3170 -1190 3240 -1130
rect 3310 -1160 3320 -1080
rect 3410 -1160 3420 -1080
rect 3310 -1170 3420 -1160
rect 3500 -1190 3570 -1130
rect 3280 -1700 3460 -1680
rect 3280 -1710 3340 -1700
rect 3280 -1750 3290 -1710
rect 3330 -1750 3340 -1710
rect 3280 -1760 3340 -1750
rect 3400 -1710 3460 -1700
rect 3400 -1750 3410 -1710
rect 3450 -1750 3460 -1710
rect 3400 -1760 3460 -1750
rect 3280 -1770 3460 -1760
rect 3640 -1820 3750 -410
rect 3830 -980 3900 -860
rect 3830 -1180 3900 -1060
rect 2980 -1890 3750 -1820
rect 3630 -2290 3690 -1890
rect 2540 -2660 4220 -2400
<< via1 >>
rect 3320 -1160 3410 -1080
rect 3340 -1760 3400 -1700
<< metal2 >>
rect 3310 -1080 3420 -1070
rect 3310 -1160 3320 -1080
rect 3410 -1160 3420 -1080
rect 3310 -1680 3420 -1160
rect 3280 -1700 3460 -1680
rect 3280 -1760 3340 -1700
rect 3400 -1760 3460 -1700
rect 3280 -1770 3460 -1760
rect 3290 -2850 3460 -1810
<< metal3 >>
rect 2460 -980 4240 -920
rect 2460 -1120 4240 -1060
use sky130_fd_pr__nfet_g5v0d10v5_JD4JK9  sky130_fd_pr__nfet_g5v0d10v5_JD4JK9_0
timestamp 1769616064
transform 1 0 3369 0 1 -646
box -795 -440 795 440
use sky130_fd_pr__nfet_g5v0d10v5_UPKHYG  sky130_fd_pr__nfet_g5v0d10v5_UPKHYG_0
timestamp 1769616064
transform 1 0 2933 0 1 -2095
box -353 -385 353 385
use sky130_fd_pr__nfet_g5v0d10v5_UPKHYG  sky130_fd_pr__nfet_g5v0d10v5_UPKHYG_1
timestamp 1769616064
transform 1 0 3813 0 1 -2095
box -353 -385 353 385
use sky130_fd_pr__nfet_g5v0d10v5_ZPYJK9  sky130_fd_pr__nfet_g5v0d10v5_ZPYJK9_0
timestamp 1769616064
transform 1 0 3365 0 1 -1400
box -795 -440 795 440
use sky130_fd_pr__pfet_g5v0d10v5_CHVBE6  XM5
timestamp 1769616064
transform 1 0 3385 0 1 365
box -845 -505 845 505
<< labels >>
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 IBIAS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VN
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VP
port 4 nsew
flabel metal1 2600 800 2800 1000 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 2600 -2600 2800 -2400 0 FreeSans 256 0 0 0 VSS
port 5 nsew
<< end >>
