magic
tech sky130A
magscale 1 2
timestamp 1770370310
<< error_s >>
rect 2649 -116034 2666 -113738
rect 2703 -116083 2720 -113787
rect 5435 -114838 5493 -114686
rect 5476 -116129 5493 -114838
rect 5494 -114838 5559 -114802
rect 5494 -114896 5645 -114838
rect 5494 -116129 5588 -114896
rect 5494 -116195 5559 -116129
rect 7073 -116224 7120 -114849
rect 7127 -116278 7174 -114903
rect 8670 -116289 8717 -114903
rect 8724 -116343 8771 -114849
rect 11467 -116354 11514 -114421
rect 14318 -114439 14376 -114323
rect 11521 -116408 11568 -114475
rect 14252 -116419 14376 -114439
rect 14452 -116253 14463 -114323
rect 19514 -114635 19572 -114483
rect 14252 -116455 14365 -116419
rect 14318 -116473 14365 -116455
rect 19555 -116484 19572 -114635
rect 19573 -114635 19638 -114599
rect 19573 -114693 19724 -114635
rect 19573 -116484 19667 -114693
rect 19573 -116550 19638 -116484
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__cap_mim_m3_1_R7S84X  XC1
timestamp 1770370310
transform 1 0 25121 0 1 -132695
box -2686 -21280 2686 21280
use sky130_fd_pr__pfet_g5v0d10v5_SFZ6J8  XM1
timestamp 1770370310
transform 1 0 1271 0 1 -114863
box -1461 -1237 1461 1237
use sky130_fd_pr__pfet_g5v0d10v5_SFZ6J8  XM2
timestamp 1770370310
transform 1 0 4098 0 1 -114958
box -1461 -1237 1461 1237
use sky130_fd_pr__nfet_g5v0d10v5_5BVNGQ  XM3
timestamp 1770370310
transform 1 0 6325 0 1 -115531
box -831 -729 831 729
use sky130_fd_pr__nfet_g5v0d10v5_5BVNGQ  XM4
timestamp 1770370310
transform 1 0 7922 0 1 -115596
box -831 -729 831 729
use sky130_fd_pr__nfet_g5v0d10v5_4AXLQQ  XM5
timestamp 1770370310
transform 1 0 10119 0 1 -115382
box -1431 -1008 1431 1008
use sky130_fd_pr__nfet_g5v0d10v5_4AXLQQ  XM6
timestamp 1770370310
transform 1 0 12916 0 1 -115447
box -1431 -1008 1431 1008
use sky130_fd_pr__pfet_g5v0d10v5_HWRH7L  XM7
timestamp 1770370310
transform 1 0 16945 0 1 -115253
box -2693 -1297 2693 1297
use sky130_fd_pr__nfet_g5v0d10v5_4AXLQQ  XM8
timestamp 1770370310
transform 1 0 21004 0 1 -115607
box -1431 -1008 1431 1008
use sky130_fd_pr__pfet_g5v0d10v5_X45ZZ5  XM9
timestamp 1770370310
transform 1 0 28417 0 1 -153273
box -705 -797 705 797
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VP
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VN
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 IBIAS
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VSS
port 5 nsew
<< end >>
