magic
tech sky130A
magscale 1 2
timestamp 1769076474
<< pwell >>
rect -515 -466 515 466
<< mvnmos >>
rect -287 -208 -187 208
rect -129 -208 -29 208
rect 29 -208 129 208
rect 187 -208 287 208
<< mvndiff >>
rect -345 196 -287 208
rect -345 -196 -333 196
rect -299 -196 -287 196
rect -345 -208 -287 -196
rect -187 196 -129 208
rect -187 -196 -175 196
rect -141 -196 -129 196
rect -187 -208 -129 -196
rect -29 196 29 208
rect -29 -196 -17 196
rect 17 -196 29 196
rect -29 -208 29 -196
rect 129 196 187 208
rect 129 -196 141 196
rect 175 -196 187 196
rect 129 -208 187 -196
rect 287 196 345 208
rect 287 -196 299 196
rect 333 -196 345 196
rect 287 -208 345 -196
<< mvndiffc >>
rect -333 -196 -299 196
rect -175 -196 -141 196
rect -17 -196 17 196
rect 141 -196 175 196
rect 299 -196 333 196
<< mvpsubdiff >>
rect -479 418 479 430
rect -479 384 -371 418
rect 371 384 479 418
rect -479 372 479 384
rect -479 322 -421 372
rect -479 -322 -467 322
rect -433 -322 -421 322
rect 421 322 479 372
rect -479 -372 -421 -322
rect 421 -322 433 322
rect 467 -322 479 322
rect 421 -372 479 -322
rect -479 -384 479 -372
rect -479 -418 -371 -384
rect 371 -418 479 -384
rect -479 -430 479 -418
<< mvpsubdiffcont >>
rect -371 384 371 418
rect -467 -322 -433 322
rect 433 -322 467 322
rect -371 -418 371 -384
<< poly >>
rect -287 280 -187 296
rect -287 246 -271 280
rect -203 246 -187 280
rect -287 208 -187 246
rect -129 280 -29 296
rect -129 246 -113 280
rect -45 246 -29 280
rect -129 208 -29 246
rect 29 280 129 296
rect 29 246 45 280
rect 113 246 129 280
rect 29 208 129 246
rect 187 280 287 296
rect 187 246 203 280
rect 271 246 287 280
rect 187 208 287 246
rect -287 -246 -187 -208
rect -287 -280 -271 -246
rect -203 -280 -187 -246
rect -287 -296 -187 -280
rect -129 -246 -29 -208
rect -129 -280 -113 -246
rect -45 -280 -29 -246
rect -129 -296 -29 -280
rect 29 -246 129 -208
rect 29 -280 45 -246
rect 113 -280 129 -246
rect 29 -296 129 -280
rect 187 -246 287 -208
rect 187 -280 203 -246
rect 271 -280 287 -246
rect 187 -296 287 -280
<< polycont >>
rect -271 246 -203 280
rect -113 246 -45 280
rect 45 246 113 280
rect 203 246 271 280
rect -271 -280 -203 -246
rect -113 -280 -45 -246
rect 45 -280 113 -246
rect 203 -280 271 -246
<< locali >>
rect -467 384 -371 418
rect 371 384 467 418
rect -467 322 -433 384
rect 433 322 467 384
rect -287 246 -271 280
rect -203 246 -187 280
rect -129 246 -113 280
rect -45 246 -29 280
rect 29 246 45 280
rect 113 246 129 280
rect 187 246 203 280
rect 271 246 287 280
rect -333 196 -299 212
rect -333 -212 -299 -196
rect -175 196 -141 212
rect -175 -212 -141 -196
rect -17 196 17 212
rect -17 -212 17 -196
rect 141 196 175 212
rect 141 -212 175 -196
rect 299 196 333 212
rect 299 -212 333 -196
rect -287 -280 -271 -246
rect -203 -280 -187 -246
rect -129 -280 -113 -246
rect -45 -280 -29 -246
rect 29 -280 45 -246
rect 113 -280 129 -246
rect 187 -280 203 -246
rect 271 -280 287 -246
rect -467 -384 -433 -322
rect 433 -384 467 -322
rect -467 -418 -371 -384
rect 371 -418 467 -384
<< viali >>
rect -271 246 -203 280
rect -113 246 -45 280
rect 45 246 113 280
rect 203 246 271 280
rect -333 -196 -299 196
rect -175 -196 -141 196
rect -17 -196 17 196
rect 141 -196 175 196
rect 299 -196 333 196
rect -271 -280 -203 -246
rect -113 -280 -45 -246
rect 45 -280 113 -246
rect 203 -280 271 -246
<< metal1 >>
rect -283 280 -191 286
rect -283 246 -271 280
rect -203 246 -191 280
rect -283 240 -191 246
rect -125 280 -33 286
rect -125 246 -113 280
rect -45 246 -33 280
rect -125 240 -33 246
rect 33 280 125 286
rect 33 246 45 280
rect 113 246 125 280
rect 33 240 125 246
rect 191 280 283 286
rect 191 246 203 280
rect 271 246 283 280
rect 191 240 283 246
rect -339 196 -293 208
rect -339 -196 -333 196
rect -299 -196 -293 196
rect -339 -208 -293 -196
rect -181 196 -135 208
rect -181 -196 -175 196
rect -141 -196 -135 196
rect -181 -208 -135 -196
rect -23 196 23 208
rect -23 -196 -17 196
rect 17 -196 23 196
rect -23 -208 23 -196
rect 135 196 181 208
rect 135 -196 141 196
rect 175 -196 181 196
rect 135 -208 181 -196
rect 293 196 339 208
rect 293 -196 299 196
rect 333 -196 339 196
rect 293 -208 339 -196
rect -283 -246 -191 -240
rect -283 -280 -271 -246
rect -203 -280 -191 -246
rect -283 -286 -191 -280
rect -125 -246 -33 -240
rect -125 -280 -113 -246
rect -45 -280 -33 -246
rect -125 -286 -33 -280
rect 33 -246 125 -240
rect 33 -280 45 -246
rect 113 -280 125 -246
rect 33 -286 125 -280
rect 191 -246 283 -240
rect 191 -280 203 -246
rect 271 -280 283 -246
rect 191 -286 283 -280
<< properties >>
string FIXED_BBOX -450 -401 450 401
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.08 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
