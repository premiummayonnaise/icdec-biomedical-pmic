* NGSPICE file created from diff-pair.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_X57ESK a_n187_n506# a_n345_n506# a_129_n506#
+ a_287_n506# a_29_n532# a_n129_n532# a_187_n532# a_n287_n532# a_n29_n506# VSUBS
X0 a_n187_n506# a_n287_n532# a_n345_n506# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=1.3775 ps=10.08 w=4.75 l=0.5
X1 a_287_n506# a_187_n532# a_129_n506# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.3775 pd=10.08 as=0.68875 ps=5.04 w=4.75 l=0.5
X2 a_129_n506# a_29_n532# a_n29_n506# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=0.68875 ps=5.04 w=4.75 l=0.5
X3 a_n29_n506# a_n129_n532# a_n187_n506# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=0.68875 ps=5.04 w=4.75 l=0.5
C0 a_n29_n506# a_29_n532# 0.05102f
C1 a_129_n506# a_287_n506# 0.34129f
C2 a_n29_n506# a_129_n506# 0.34129f
C3 a_n29_n506# a_n187_n506# 0.34129f
C4 a_129_n506# a_29_n532# 0.05102f
C5 a_n29_n506# a_n129_n532# 0.05102f
C6 a_n129_n532# a_29_n532# 0.05942f
C7 a_287_n506# a_187_n532# 0.05102f
C8 a_n287_n532# a_n187_n506# 0.05102f
C9 a_n287_n532# a_n129_n532# 0.05942f
C10 a_n187_n506# a_n129_n532# 0.05102f
C11 a_n287_n532# a_n345_n506# 0.05102f
C12 a_187_n532# a_29_n532# 0.05942f
C13 a_n187_n506# a_n345_n506# 0.34129f
C14 a_129_n506# a_187_n532# 0.05102f
C15 a_287_n506# VSUBS 0.36723f
C16 a_129_n506# VSUBS 0.08691f
C17 a_n29_n506# VSUBS 0.08691f
C18 a_n187_n506# VSUBS 0.08691f
C19 a_n345_n506# VSUBS 0.36723f
C20 a_187_n532# VSUBS 0.25901f
C21 a_29_n532# VSUBS 0.2242f
C22 a_n129_n532# VSUBS 0.2242f
C23 a_n287_n532# VSUBS 0.25901f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SNDLS5 a_n29_n444# a_n187_n444# a_n345_n444#
+ a_29_n532# a_n129_n532# a_187_n532# a_129_n444# a_n287_n532# a_287_n444# VSUBS
X0 a_129_n444# a_29_n532# a_n29_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=0.68875 ps=5.04 w=4.75 l=0.5
X1 a_n29_n444# a_n129_n532# a_n187_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=0.68875 ps=5.04 w=4.75 l=0.5
X2 a_n187_n444# a_n287_n532# a_n345_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=1.3775 ps=10.08 w=4.75 l=0.5
X3 a_287_n444# a_187_n532# a_129_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.3775 pd=10.08 as=0.68875 ps=5.04 w=4.75 l=0.5
C0 a_n345_n444# a_n187_n444# 0.34523f
C1 a_n187_n444# a_n29_n444# 0.34523f
C2 a_n129_n532# a_n287_n532# 0.05942f
C3 a_129_n444# a_187_n532# 0.05102f
C4 a_n129_n532# a_n187_n444# 0.05102f
C5 a_187_n532# a_29_n532# 0.05942f
C6 a_187_n532# a_n29_n444# 0.00651f
C7 a_187_n532# a_287_n444# 0.05885f
C8 a_n187_n444# a_n287_n532# 0.05102f
C9 a_129_n444# a_29_n532# 0.05102f
C10 a_129_n444# a_n29_n444# 0.34523f
C11 a_n345_n444# a_n29_n444# 0.03881f
C12 a_129_n444# a_287_n444# 0.34523f
C13 a_29_n532# a_n29_n444# 0.05885f
C14 a_29_n532# a_287_n444# 0.00651f
C15 a_287_n444# a_n29_n444# 0.03881f
C16 a_n129_n532# a_n345_n444# 0.00651f
C17 a_29_n532# a_n129_n532# 0.05942f
C18 a_n129_n532# a_n29_n444# 0.05885f
C19 a_n345_n444# a_n287_n532# 0.05885f
C20 a_n287_n532# a_n29_n444# 0.00651f
C21 a_287_n444# VSUBS 0.4557f
C22 a_129_n444# VSUBS 0.08691f
C23 a_n29_n444# VSUBS 0.1204f
C24 a_n187_n444# VSUBS 0.08691f
C25 a_n345_n444# VSUBS 0.4557f
C26 a_187_n532# VSUBS 0.25901f
C27 a_29_n532# VSUBS 0.2242f
C28 a_n129_n532# VSUBS 0.2242f
C29 a_n287_n532# VSUBS 0.25901f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH a_n29_n444# a_n187_n444# a_n345_n444#
+ a_29_n532# a_n129_n532# a_187_n532# a_129_n444# a_n287_n532# a_287_n444# VSUBS
X0 a_129_n444# a_29_n532# a_n29_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=0.68875 ps=5.04 w=4.75 l=0.5
X1 a_n29_n444# a_n129_n532# a_n187_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=0.68875 ps=5.04 w=4.75 l=0.5
X2 a_n187_n444# a_n287_n532# a_n345_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=1.3775 ps=10.08 w=4.75 l=0.5
X3 a_287_n444# a_187_n532# a_129_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.3775 pd=10.08 as=0.68875 ps=5.04 w=4.75 l=0.5
C0 a_n129_n532# a_29_n532# 0.05942f
C1 a_n29_n444# a_n187_n444# 0.34129f
C2 a_29_n532# a_187_n532# 0.05942f
C3 a_n345_n444# a_n287_n532# 0.05102f
C4 a_n29_n444# a_129_n444# 0.34129f
C5 a_n287_n532# a_n129_n532# 0.05942f
C6 a_29_n532# a_129_n444# 0.05102f
C7 a_n287_n532# a_n187_n444# 0.05102f
C8 a_29_n532# a_n29_n444# 0.05102f
C9 a_n345_n444# a_n187_n444# 0.34129f
C10 a_n129_n532# a_n187_n444# 0.05102f
C11 a_287_n444# a_187_n532# 0.05102f
C12 a_129_n444# a_187_n532# 0.05102f
C13 a_n129_n532# a_n29_n444# 0.05102f
C14 a_287_n444# a_129_n444# 0.34129f
C15 a_287_n444# VSUBS 0.36723f
C16 a_129_n444# VSUBS 0.08691f
C17 a_n29_n444# VSUBS 0.08691f
C18 a_n187_n444# VSUBS 0.08691f
C19 a_n345_n444# VSUBS 0.36723f
C20 a_187_n532# VSUBS 0.25901f
C21 a_29_n532# VSUBS 0.2242f
C22 a_n129_n532# VSUBS 0.2242f
C23 a_n287_n532# VSUBS 0.25901f
.ends

.subckt diff-pair VP VN S D2 D1 VSS
Xsky130_fd_pr__nfet_g5v0d10v5_X57ESK_0 D1 D1 D1 D1 VP VP D1 D1 S VSS sky130_fd_pr__nfet_g5v0d10v5_X57ESK
Xsky130_fd_pr__nfet_g5v0d10v5_SNDLS5_0 S D2 D2 VN VN D2 D2 D2 D2 VSS sky130_fd_pr__nfet_g5v0d10v5_SNDLS5
Xsky130_fd_pr__nfet_g5v0d10v5_X57ESK_1 D1 D1 D1 D1 VP VP D1 D1 S VSS sky130_fd_pr__nfet_g5v0d10v5_X57ESK
Xsky130_fd_pr__nfet_g5v0d10v5_X57ESK_2 D1 D1 D1 D1 VP VP D1 D1 S VSS sky130_fd_pr__nfet_g5v0d10v5_X57ESK
Xsky130_fd_pr__nfet_g5v0d10v5_X57ESK_3 D1 D1 D1 D1 VP VP D1 D1 S VSS sky130_fd_pr__nfet_g5v0d10v5_X57ESK
Xsky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_0 S D2 D2 VN VN D2 D2 D2 D2 VSS sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH
Xsky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_1 S D2 D2 VN VN D2 D2 D2 D2 VSS sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH
Xsky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_2 S D2 D2 VN VN D2 D2 D2 D2 VSS sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH
C0 S a_6410_210# 0.01107f
C1 a_3710_2090# VP 0.00281f
C2 a_5210_200# D1 0.12337f
C3 a_4420_2100# D1 0.01332f
C4 VP a_4420_200# 0.01038f
C5 S a_2920_2100# 0.01618f
C6 a_1720_200# D2 0.13361f
C7 a_5210_2100# VP 0.03078f
C8 VP a_2510_2100# 0.04468f
C9 a_5620_200# D2 0.12979f
C10 a_3710_2090# D1 0.01306f
C11 a_6410_2100# VP 0.00358f
C12 a_2920_200# a_2920_2100# 0.00109f
C13 VP D1 2.1751f
C14 VN S 6.91268f
C15 a_4420_200# D1 0.11957f
C16 S a_2510_200# 0.01284f
C17 S a_1720_2100# 0.01132f
C18 a_5210_2100# D1 0.02102f
C19 a_2510_2100# D1 0.12736f
C20 a_3720_200# D2 0.01484f
C21 a_4420_2100# a_2920_2100# 0.00461f
C22 a_5620_2100# VP 0.045f
C23 VN a_2920_200# 0.00181f
C24 a_6410_2100# D1 0.13685f
C25 a_1720_200# S 0.0118f
C26 a_2510_200# a_2920_200# 0.04663f
C27 VP a_6410_210# 0.01049f
C28 a_5620_2100# a_5210_2100# 0.04663f
C29 S a_5620_200# 0.01261f
C30 a_3710_2090# a_2920_2100# 0.01133f
C31 VN a_5210_200# 0.00173f
C32 VP a_2920_2100# 0.03133f
C33 a_5620_2100# a_6410_2100# 0.02082f
C34 a_4420_2100# VN 0.01013f
C35 a_5620_2100# D1 0.1257f
C36 a_6410_2100# a_6410_210# 0.00108f
C37 D1 a_6410_210# 0.01737f
C38 a_2510_2100# a_2920_2100# 0.04663f
C39 a_3710_2090# VN 0.0109f
C40 VP VN 1.71011f
C41 S D2 3.74033f
C42 S a_3720_200# 0.13056f
C43 D1 a_2920_2100# 0.02172f
C44 VN a_4420_200# 0
C45 VP a_2510_200# 0.01092f
C46 VP a_1720_2100# 0.00351f
C47 a_5210_2100# VN 0.01013f
C48 a_5620_200# a_5210_200# 0.04571f
C49 VN a_2510_2100# 0.01013f
C50 a_2510_2100# a_2510_200# 0.00109f
C51 a_2920_200# D2 0.02516f
C52 a_2510_2100# a_1720_2100# 0.02082f
C53 a_3720_200# a_2920_200# 0.02054f
C54 a_6410_2100# VN 0.01013f
C55 a_1720_200# VP 0.01092f
C56 VN D1 1.44046f
C57 a_2510_200# D1 0.02386f
C58 D1 a_1720_2100# 0.13423f
C59 VP a_5620_200# 0.0101f
C60 a_5210_200# D2 0.02436f
C61 a_4420_2100# D2 0.13065f
C62 a_5620_2100# VN 0.01013f
C63 a_1720_200# D1 0.01752f
C64 VN a_6410_210# 0.04315f
C65 a_3710_2090# D2 0.1323f
C66 a_3710_2090# a_3720_200# 0
C67 a_5620_200# D1 0.02396f
C68 VP D2 1.7381f
C69 VP a_3720_200# 0.0112f
C70 S a_2920_200# 0.01404f
C71 VN a_2920_2100# 0.01013f
C72 a_4420_200# D2 0.01395f
C73 a_3720_200# a_4420_200# 0.01595f
C74 a_5210_2100# D2 0.128f
C75 a_2510_2100# D2 0.02128f
C76 a_5620_2100# a_5620_200# 0.00107f
C77 S a_5210_200# 0.01411f
C78 a_6410_2100# D2 0.01857f
C79 a_4420_2100# S 0.13132f
C80 D1 D2 10.72437f
C81 a_5620_200# a_6410_210# 0.01999f
C82 a_3720_200# D1 0.12743f
C83 VN a_2510_200# 0.00331f
C84 VN a_1720_2100# 0.01013f
C85 a_3710_2090# S 0.12441f
C86 VP S 7.19749f
C87 a_5620_2100# D2 0.02085f
C88 S a_4420_200# 0.12752f
C89 a_1720_200# VN 0.04439f
C90 D2 a_6410_210# 0.13273f
C91 a_5210_2100# S 0.01234f
C92 a_1720_200# a_2510_200# 0.02043f
C93 a_1720_200# a_1720_2100# 0.00109f
C94 S a_2510_2100# 0.01121f
C95 VN a_5620_200# 0.00316f
C96 VP a_2920_200# 0.0112f
C97 a_6410_2100# S 0.01089f
C98 a_2920_2100# D2 0.13272f
C99 S D1 3.32348f
C100 VP a_5210_200# 0.01039f
C101 a_4420_2100# a_3710_2090# 0.02486f
C102 a_4420_2100# VP 0.00273f
C103 a_5210_200# a_4420_200# 0.02082f
C104 a_2920_200# D1 0.12627f
C105 VN D2 2.00876f
C106 VN a_3720_200# 0
C107 a_5210_2100# a_5210_200# 0.00107f
C108 a_4420_2100# a_4420_200# 0.00107f
C109 a_5620_2100# S 0.01133f
C110 a_4420_2100# a_5210_2100# 0.02043f
C111 a_2510_200# D2 0.13428f
C112 a_1720_2100# D2 0.01861f
C113 a_6410_210# VSS 0.73929f $ **FLOATING
C114 a_5620_200# VSS 0.68028f $ **FLOATING
C115 a_5210_200# VSS 0.68003f $ **FLOATING
C116 a_4420_200# VSS 0.69659f $ **FLOATING
C117 a_3720_200# VSS 0.73656f $ **FLOATING
C118 a_2920_200# VSS 0.69319f $ **FLOATING
C119 a_2510_200# VSS 0.69291f $ **FLOATING
C120 a_1720_200# VSS 0.75406f $ **FLOATING
C121 a_6410_2100# VSS 0.75393f $ **FLOATING
C122 a_5620_2100# VSS 0.69351f $ **FLOATING
C123 a_5210_2100# VSS 0.69348f $ **FLOATING
C124 a_4420_2100# VSS 0.71053f $ **FLOATING
C125 a_3710_2090# VSS 0.71095f $ **FLOATING
C126 a_2920_2100# VSS 0.69357f $ **FLOATING
C127 a_2510_2100# VSS 0.69349f $ **FLOATING
C128 a_1720_2100# VSS 0.75462f $ **FLOATING
C129 D2 VSS 7.92398f
C130 VN VSS 5.76024f
C131 VP VSS 5.14956f
C132 D1 VSS 9.47276f
C133 S VSS 9.00222f
.ends

