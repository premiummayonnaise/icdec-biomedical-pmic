magic
tech sky130A
magscale 1 2
timestamp 1769437396
<< nwell >>
rect 10140 -73228 32340 -67028
<< pwell >>
rect -2900 -79100 800 -72600
rect -30800 -89700 9000 -83400
<< psubdiff >>
rect -2900 -72900 800 -72600
rect -2900 -78800 -2600 -72900
rect 500 -78800 800 -72900
rect -2900 -79100 800 -78800
rect -30800 -83480 9000 -83400
rect -30800 -83840 -30300 -83480
rect 8500 -83840 9000 -83480
rect -30800 -83900 9000 -83840
rect -30800 -89200 -30740 -83900
rect -30360 -89200 -30300 -83900
rect 8500 -89200 8560 -83900
rect 8940 -89200 9000 -83900
rect -30800 -89280 9000 -89200
rect -30800 -89640 -30300 -89280
rect 8500 -89640 9000 -89280
rect -30800 -89700 9000 -89640
<< nsubdiff >>
rect 10240 -67228 32240 -67128
rect 10240 -67528 10740 -67228
rect 31740 -67528 32240 -67228
rect 10240 -67628 32240 -67528
rect 10240 -72628 10340 -67628
rect 10640 -72628 10740 -67628
rect 31740 -72628 31840 -67628
rect 32140 -72628 32240 -67628
rect 10240 -72728 32240 -72628
rect 10240 -73028 10740 -72728
rect 31740 -73028 32240 -72728
rect 10240 -73128 32240 -73028
<< psubdiffcont >>
rect -30300 -83840 8500 -83480
rect -30740 -89200 -30360 -83900
rect 8560 -89200 8940 -83900
rect -30300 -89640 8500 -89280
<< nsubdiffcont >>
rect 10740 -67528 31740 -67228
rect 10340 -72628 10640 -67628
rect 31840 -72628 32140 -67628
rect 10740 -73028 31740 -72728
<< xpolycontact >>
rect -1600 -73500 -1530 -73068
rect -1600 -78600 -1530 -78168
rect -1400 -73500 -1330 -73068
rect -1400 -78600 -1330 -78168
rect -1200 -73500 -1130 -73068
rect -1200 -78600 -1130 -78168
rect -1000 -73500 -930 -73068
rect -1000 -78600 -930 -78168
rect -800 -73500 -730 -73068
rect -800 -78600 -730 -78168
rect -600 -73500 -530 -73068
rect -600 -78600 -530 -78168
rect -400 -73500 -330 -73068
rect -400 -78600 -330 -78168
rect -200 -73500 -130 -73068
rect -200 -78600 -130 -78168
<< ppolyres >>
rect -1600 -78168 -1530 -73500
rect -1400 -78168 -1330 -73500
rect -1200 -78168 -1130 -73500
rect -1000 -78168 -930 -73500
rect -800 -78168 -730 -73500
rect -600 -78168 -530 -73500
rect -400 -78168 -330 -73500
rect -200 -78168 -130 -73500
<< locali >>
rect 10240 -67228 32240 -67128
rect 10240 -67528 10740 -67228
rect 31740 -67528 32240 -67228
rect 10240 -67628 32240 -67528
rect -2900 -72900 800 -72600
rect -2900 -78800 -2600 -72900
rect 500 -78800 800 -72900
rect 10240 -72628 10340 -67628
rect 10640 -72628 10740 -67628
rect 31740 -72628 31840 -67628
rect 32140 -72628 32240 -67628
rect 10240 -72728 32240 -72628
rect 10240 -73028 10740 -72728
rect 31740 -73028 32240 -72728
rect 10240 -73128 32240 -73028
rect -2900 -79100 800 -78800
rect -30800 -83480 9000 -83400
rect -30800 -83840 -30300 -83480
rect 8500 -83840 9000 -83480
rect -30800 -83900 9000 -83840
rect -30800 -89200 -30740 -83900
rect -30360 -89200 -30300 -83900
rect 8500 -89200 8560 -83900
rect 8940 -89200 9000 -83900
rect -30800 -89280 9000 -89200
rect -30800 -89640 -30300 -89280
rect 8500 -89640 9000 -89280
rect -30800 -89700 9000 -89640
<< viali >>
rect -1584 -73483 -1546 -73086
rect -1384 -73483 -1346 -73086
rect -1184 -73483 -1146 -73086
rect -984 -73483 -946 -73086
rect -784 -73483 -746 -73086
rect -584 -73483 -546 -73086
rect -384 -73483 -346 -73086
rect -184 -73483 -146 -73086
rect -1584 -78582 -1546 -78185
rect -1384 -78582 -1346 -78185
rect -1184 -78582 -1146 -78185
rect -984 -78582 -946 -78185
rect -784 -78582 -746 -78185
rect -584 -78582 -546 -78185
rect -384 -78582 -346 -78185
rect -184 -78582 -146 -78185
<< metal1 >>
rect -1590 -73086 -1540 -73074
rect -1590 -73483 -1584 -73086
rect -1546 -73483 -1540 -73086
rect -1590 -73495 -1540 -73483
rect -1390 -73086 -1340 -73074
rect -1390 -73483 -1384 -73086
rect -1346 -73483 -1340 -73086
rect -1390 -73495 -1340 -73483
rect -1190 -73086 -1140 -73074
rect -1190 -73483 -1184 -73086
rect -1146 -73483 -1140 -73086
rect -1190 -73495 -1140 -73483
rect -990 -73086 -940 -73074
rect -990 -73483 -984 -73086
rect -946 -73483 -940 -73086
rect -990 -73495 -940 -73483
rect -790 -73086 -740 -73074
rect -790 -73483 -784 -73086
rect -746 -73483 -740 -73086
rect -790 -73495 -740 -73483
rect -590 -73086 -540 -73074
rect -590 -73483 -584 -73086
rect -546 -73483 -540 -73086
rect -590 -73495 -540 -73483
rect -390 -73086 -340 -73074
rect -390 -73483 -384 -73086
rect -346 -73483 -340 -73086
rect -390 -73495 -340 -73483
rect -190 -73086 -140 -73074
rect -190 -73483 -184 -73086
rect -146 -73483 -140 -73086
rect -190 -73495 -140 -73483
rect -1590 -78185 -1540 -78173
rect -1590 -78582 -1584 -78185
rect -1546 -78582 -1540 -78185
rect -1590 -78594 -1540 -78582
rect -1390 -78185 -1340 -78173
rect -1390 -78582 -1384 -78185
rect -1346 -78582 -1340 -78185
rect -1390 -78594 -1340 -78582
rect -1190 -78185 -1140 -78173
rect -1190 -78582 -1184 -78185
rect -1146 -78582 -1140 -78185
rect -1190 -78594 -1140 -78582
rect -990 -78185 -940 -78173
rect -990 -78582 -984 -78185
rect -946 -78582 -940 -78185
rect -990 -78594 -940 -78582
rect -790 -78185 -740 -78173
rect -790 -78582 -784 -78185
rect -746 -78582 -740 -78185
rect -790 -78594 -740 -78582
rect -590 -78185 -540 -78173
rect -590 -78582 -584 -78185
rect -546 -78582 -540 -78185
rect -590 -78594 -540 -78582
rect -390 -78185 -340 -78173
rect -390 -78582 -384 -78185
rect -346 -78582 -340 -78185
rect -390 -78594 -340 -78582
rect -190 -78185 -140 -78173
rect -190 -78582 -184 -78185
rect -146 -78582 -140 -78185
rect -190 -78594 -140 -78582
<< metal2 >>
rect -38000 -90000 -37000 -60000
rect -36000 -90000 -35000 -60000
rect -34000 -90000 -33000 -60000
<< metal4 >>
rect -25500 -72400 6100 -72000
rect -25500 -83000 -25100 -72400
rect -19900 -83000 -19500 -72400
rect -14300 -83000 -13900 -72400
rect -8600 -83000 -8200 -72400
<< metal5 >>
rect 10140 -66428 32340 -60228
rect 10140 -74238 32340 -74228
rect 10130 -80428 32340 -74238
rect 10130 -89622 32264 -80428
use err-amp  err-amp_0 /foss/designs/icdec-biomedical-pmic/xschem/error-amplifier/layout
timestamp 1769436194
transform 1 0 -31680 0 1 -67800
box -320 -4200 38300 7200
use sky130_fd_pr__pfet_g5v0d10v5_PYEB7S  sky130_fd_pr__pfet_g5v0d10v5_PYEB7S_0
timestamp 1769436194
transform 1 0 21171 0 1 -69995
box -8931 -1133 8931 1095
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_0
timestamp 1769436194
transform 1 0 -1765 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_1
timestamp 1769436194
transform 1 0 -1365 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_2
timestamp 1769436194
transform 1 0 -1565 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_3
timestamp 1769436194
transform 1 0 -765 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_4
timestamp 1769436194
transform 1 0 -565 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_5
timestamp 1769436194
transform 1 0 -1165 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_6
timestamp 1769436194
transform 1 0 -965 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_7
timestamp 1769436194
transform 1 0 -165 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  sky130_fd_pr__res_high_po_0p35_L4KQ4L_8
timestamp 1769436194
transform 1 0 -365 0 1 -75834
box -35 -2766 35 2766
use sky130_fd_pr__cap_mim_m3_1_RKP84X  XC2
timestamp 1769436194
transform 1 0 -19596 0 1 -77780
box -11104 -5320 11104 5320
use sky130_fd_pr__pfet_g5v0d10v5_6DTU7R  XM1
timestamp 1769436194
transform 1 0 -5739 0 1 -78103
box -861 -797 861 797
use sky130_fd_pr__nfet_g5v0d10v5_YZ2G8N  XM3
timestamp 1769436194
transform 1 0 -10839 0 1 -86543
box -17761 -2057 17761 2057
use sky130_fd_pr__res_high_po_2p85_HMPA8M  XR1
timestamp 1769436194
transform -1 0 -952 0 -1 -81268
box -3448 -1932 3448 1932
use sky130_fd_pr__res_high_po_0p35_L4KQ4L  XR2
timestamp 1769436194
transform 1 0 -1965 0 1 -75834
box -35 -2766 35 2766
<< end >>
