** sch_path: /foss/designs/icdec-biomedical-pmic/xschem/bandgap/bgr_ota/bgr-ota.sch
.subckt bgr-ota VDD OUT VP VN VSS
*.PININFO VSS:B VDD:B VP:I VN:I OUT:O
XM1 net1 VP net3 VSS sky130_fd_pr__nfet_01v8 L=0.3 W=2.5 nf=2 m=1
XM2 net2 VN net3 VSS sky130_fd_pr__nfet_01v8 L=0.3 W=2.5 nf=2 m=1
XM4 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=1.25 W=10.8 nf=4 m=1
XM5 net1 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=1.25 W=10.8 nf=4 m=1
XM6 net3 IB VSS VSS sky130_fd_pr__nfet_01v8 L=1.25 W=3.4 nf=1 m=1
XM3 IB net5 net4 net4 sky130_fd_pr__nfet_01v8 L=1.25 W=3.4 nf=1 m=1
XM7 IB IB VDD VDD sky130_fd_pr__pfet_01v8 L=1.25 W=10.8 nf=4 m=1
XM8 net5 IB VDD VDD sky130_fd_pr__pfet_01v8 L=1.25 W=10.8 nf=4 m=1
XM9 net5 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=1.25 W=3.4 nf=1 m=1
XM11 OUT net2 VDD VDD sky130_fd_pr__pfet_01v8 L=1.25 W=110 nf=32 m=1
XM12 OUT IB VSS VSS sky130_fd_pr__nfet_01v8 L=1.25 W=10 nf=4 m=1
XC1 OUT net2 sky130_fd_pr__cap_mim_m3_1 W=20 L=20 m=4
XM14 IB IB net5 net5 sky130_fd_pr__nfet_01v8 L=0.15 W=0.85 nf=1 m=1
XR1 net6 net4 VSS sky130_fd_pr__res_high_po_1p41 L=3.235 mult=1 m=1
XR2 net8 net6 VSS sky130_fd_pr__res_high_po_1p41 L=3.235 mult=1 m=1
XR3 net7 net8 VSS sky130_fd_pr__res_high_po_1p41 L=3.235 mult=1 m=1
XR4 net9 net7 VSS sky130_fd_pr__res_high_po_1p41 L=3.235 mult=1 m=1
XR5 VSS net9 VSS sky130_fd_pr__res_high_po_1p41 L=3.235 mult=1 m=1
.ends
