magic
tech sky130A
magscale 1 2
timestamp 1770112220
<< nwell >>
rect -2693 -1237 2693 1237
<< mvpmos >>
rect -2435 -940 -2185 940
rect -2127 -940 -1877 940
rect -1819 -940 -1569 940
rect -1511 -940 -1261 940
rect -1203 -940 -953 940
rect -895 -940 -645 940
rect -587 -940 -337 940
rect -279 -940 -29 940
rect 29 -940 279 940
rect 337 -940 587 940
rect 645 -940 895 940
rect 953 -940 1203 940
rect 1261 -940 1511 940
rect 1569 -940 1819 940
rect 1877 -940 2127 940
rect 2185 -940 2435 940
<< mvpdiff >>
rect -2493 928 -2435 940
rect -2493 -928 -2481 928
rect -2447 -928 -2435 928
rect -2493 -940 -2435 -928
rect -2185 928 -2127 940
rect -2185 -928 -2173 928
rect -2139 -928 -2127 928
rect -2185 -940 -2127 -928
rect -1877 928 -1819 940
rect -1877 -928 -1865 928
rect -1831 -928 -1819 928
rect -1877 -940 -1819 -928
rect -1569 928 -1511 940
rect -1569 -928 -1557 928
rect -1523 -928 -1511 928
rect -1569 -940 -1511 -928
rect -1261 928 -1203 940
rect -1261 -928 -1249 928
rect -1215 -928 -1203 928
rect -1261 -940 -1203 -928
rect -953 928 -895 940
rect -953 -928 -941 928
rect -907 -928 -895 928
rect -953 -940 -895 -928
rect -645 928 -587 940
rect -645 -928 -633 928
rect -599 -928 -587 928
rect -645 -940 -587 -928
rect -337 928 -279 940
rect -337 -928 -325 928
rect -291 -928 -279 928
rect -337 -940 -279 -928
rect -29 928 29 940
rect -29 -928 -17 928
rect 17 -928 29 928
rect -29 -940 29 -928
rect 279 928 337 940
rect 279 -928 291 928
rect 325 -928 337 928
rect 279 -940 337 -928
rect 587 928 645 940
rect 587 -928 599 928
rect 633 -928 645 928
rect 587 -940 645 -928
rect 895 928 953 940
rect 895 -928 907 928
rect 941 -928 953 928
rect 895 -940 953 -928
rect 1203 928 1261 940
rect 1203 -928 1215 928
rect 1249 -928 1261 928
rect 1203 -940 1261 -928
rect 1511 928 1569 940
rect 1511 -928 1523 928
rect 1557 -928 1569 928
rect 1511 -940 1569 -928
rect 1819 928 1877 940
rect 1819 -928 1831 928
rect 1865 -928 1877 928
rect 1819 -940 1877 -928
rect 2127 928 2185 940
rect 2127 -928 2139 928
rect 2173 -928 2185 928
rect 2127 -940 2185 -928
rect 2435 928 2493 940
rect 2435 -928 2447 928
rect 2481 -928 2493 928
rect 2435 -940 2493 -928
<< mvpdiffc >>
rect -2481 -928 -2447 928
rect -2173 -928 -2139 928
rect -1865 -928 -1831 928
rect -1557 -928 -1523 928
rect -1249 -928 -1215 928
rect -941 -928 -907 928
rect -633 -928 -599 928
rect -325 -928 -291 928
rect -17 -928 17 928
rect 291 -928 325 928
rect 599 -928 633 928
rect 907 -928 941 928
rect 1215 -928 1249 928
rect 1523 -928 1557 928
rect 1831 -928 1865 928
rect 2139 -928 2173 928
rect 2447 -928 2481 928
<< mvnsubdiff >>
rect -2627 1159 2627 1171
rect -2627 1125 -2519 1159
rect 2519 1125 2627 1159
rect -2627 1113 2627 1125
rect -2627 1063 -2569 1113
rect -2627 -1063 -2615 1063
rect -2581 -1063 -2569 1063
rect 2569 1063 2627 1113
rect -2627 -1113 -2569 -1063
rect 2569 -1063 2581 1063
rect 2615 -1063 2627 1063
rect 2569 -1113 2627 -1063
rect -2627 -1125 2627 -1113
rect -2627 -1159 -2519 -1125
rect 2519 -1159 2627 -1125
rect -2627 -1171 2627 -1159
<< mvnsubdiffcont >>
rect -2519 1125 2519 1159
rect -2615 -1063 -2581 1063
rect 2581 -1063 2615 1063
rect -2519 -1159 2519 -1125
<< poly >>
rect -2435 1021 -2185 1037
rect -2435 987 -2419 1021
rect -2201 987 -2185 1021
rect -2435 940 -2185 987
rect -2127 1021 -1877 1037
rect -2127 987 -2111 1021
rect -1893 987 -1877 1021
rect -2127 940 -1877 987
rect -1819 1021 -1569 1037
rect -1819 987 -1803 1021
rect -1585 987 -1569 1021
rect -1819 940 -1569 987
rect -1511 1021 -1261 1037
rect -1511 987 -1495 1021
rect -1277 987 -1261 1021
rect -1511 940 -1261 987
rect -1203 1021 -953 1037
rect -1203 987 -1187 1021
rect -969 987 -953 1021
rect -1203 940 -953 987
rect -895 1021 -645 1037
rect -895 987 -879 1021
rect -661 987 -645 1021
rect -895 940 -645 987
rect -587 1021 -337 1037
rect -587 987 -571 1021
rect -353 987 -337 1021
rect -587 940 -337 987
rect -279 1021 -29 1037
rect -279 987 -263 1021
rect -45 987 -29 1021
rect -279 940 -29 987
rect 29 1021 279 1037
rect 29 987 45 1021
rect 263 987 279 1021
rect 29 940 279 987
rect 337 1021 587 1037
rect 337 987 353 1021
rect 571 987 587 1021
rect 337 940 587 987
rect 645 1021 895 1037
rect 645 987 661 1021
rect 879 987 895 1021
rect 645 940 895 987
rect 953 1021 1203 1037
rect 953 987 969 1021
rect 1187 987 1203 1021
rect 953 940 1203 987
rect 1261 1021 1511 1037
rect 1261 987 1277 1021
rect 1495 987 1511 1021
rect 1261 940 1511 987
rect 1569 1021 1819 1037
rect 1569 987 1585 1021
rect 1803 987 1819 1021
rect 1569 940 1819 987
rect 1877 1021 2127 1037
rect 1877 987 1893 1021
rect 2111 987 2127 1021
rect 1877 940 2127 987
rect 2185 1021 2435 1037
rect 2185 987 2201 1021
rect 2419 987 2435 1021
rect 2185 940 2435 987
rect -2435 -987 -2185 -940
rect -2435 -1021 -2419 -987
rect -2201 -1021 -2185 -987
rect -2435 -1037 -2185 -1021
rect -2127 -987 -1877 -940
rect -2127 -1021 -2111 -987
rect -1893 -1021 -1877 -987
rect -2127 -1037 -1877 -1021
rect -1819 -987 -1569 -940
rect -1819 -1021 -1803 -987
rect -1585 -1021 -1569 -987
rect -1819 -1037 -1569 -1021
rect -1511 -987 -1261 -940
rect -1511 -1021 -1495 -987
rect -1277 -1021 -1261 -987
rect -1511 -1037 -1261 -1021
rect -1203 -987 -953 -940
rect -1203 -1021 -1187 -987
rect -969 -1021 -953 -987
rect -1203 -1037 -953 -1021
rect -895 -987 -645 -940
rect -895 -1021 -879 -987
rect -661 -1021 -645 -987
rect -895 -1037 -645 -1021
rect -587 -987 -337 -940
rect -587 -1021 -571 -987
rect -353 -1021 -337 -987
rect -587 -1037 -337 -1021
rect -279 -987 -29 -940
rect -279 -1021 -263 -987
rect -45 -1021 -29 -987
rect -279 -1037 -29 -1021
rect 29 -987 279 -940
rect 29 -1021 45 -987
rect 263 -1021 279 -987
rect 29 -1037 279 -1021
rect 337 -987 587 -940
rect 337 -1021 353 -987
rect 571 -1021 587 -987
rect 337 -1037 587 -1021
rect 645 -987 895 -940
rect 645 -1021 661 -987
rect 879 -1021 895 -987
rect 645 -1037 895 -1021
rect 953 -987 1203 -940
rect 953 -1021 969 -987
rect 1187 -1021 1203 -987
rect 953 -1037 1203 -1021
rect 1261 -987 1511 -940
rect 1261 -1021 1277 -987
rect 1495 -1021 1511 -987
rect 1261 -1037 1511 -1021
rect 1569 -987 1819 -940
rect 1569 -1021 1585 -987
rect 1803 -1021 1819 -987
rect 1569 -1037 1819 -1021
rect 1877 -987 2127 -940
rect 1877 -1021 1893 -987
rect 2111 -1021 2127 -987
rect 1877 -1037 2127 -1021
rect 2185 -987 2435 -940
rect 2185 -1021 2201 -987
rect 2419 -1021 2435 -987
rect 2185 -1037 2435 -1021
<< polycont >>
rect -2419 987 -2201 1021
rect -2111 987 -1893 1021
rect -1803 987 -1585 1021
rect -1495 987 -1277 1021
rect -1187 987 -969 1021
rect -879 987 -661 1021
rect -571 987 -353 1021
rect -263 987 -45 1021
rect 45 987 263 1021
rect 353 987 571 1021
rect 661 987 879 1021
rect 969 987 1187 1021
rect 1277 987 1495 1021
rect 1585 987 1803 1021
rect 1893 987 2111 1021
rect 2201 987 2419 1021
rect -2419 -1021 -2201 -987
rect -2111 -1021 -1893 -987
rect -1803 -1021 -1585 -987
rect -1495 -1021 -1277 -987
rect -1187 -1021 -969 -987
rect -879 -1021 -661 -987
rect -571 -1021 -353 -987
rect -263 -1021 -45 -987
rect 45 -1021 263 -987
rect 353 -1021 571 -987
rect 661 -1021 879 -987
rect 969 -1021 1187 -987
rect 1277 -1021 1495 -987
rect 1585 -1021 1803 -987
rect 1893 -1021 2111 -987
rect 2201 -1021 2419 -987
<< locali >>
rect -2615 1125 -2519 1159
rect 2519 1125 2615 1159
rect -2615 1063 -2581 1125
rect 2581 1063 2615 1125
rect -2435 987 -2419 1021
rect -2201 987 -2185 1021
rect -2127 987 -2111 1021
rect -1893 987 -1877 1021
rect -1819 987 -1803 1021
rect -1585 987 -1569 1021
rect -1511 987 -1495 1021
rect -1277 987 -1261 1021
rect -1203 987 -1187 1021
rect -969 987 -953 1021
rect -895 987 -879 1021
rect -661 987 -645 1021
rect -587 987 -571 1021
rect -353 987 -337 1021
rect -279 987 -263 1021
rect -45 987 -29 1021
rect 29 987 45 1021
rect 263 987 279 1021
rect 337 987 353 1021
rect 571 987 587 1021
rect 645 987 661 1021
rect 879 987 895 1021
rect 953 987 969 1021
rect 1187 987 1203 1021
rect 1261 987 1277 1021
rect 1495 987 1511 1021
rect 1569 987 1585 1021
rect 1803 987 1819 1021
rect 1877 987 1893 1021
rect 2111 987 2127 1021
rect 2185 987 2201 1021
rect 2419 987 2435 1021
rect -2481 928 -2447 944
rect -2481 -944 -2447 -928
rect -2173 928 -2139 944
rect -2173 -944 -2139 -928
rect -1865 928 -1831 944
rect -1865 -944 -1831 -928
rect -1557 928 -1523 944
rect -1557 -944 -1523 -928
rect -1249 928 -1215 944
rect -1249 -944 -1215 -928
rect -941 928 -907 944
rect -941 -944 -907 -928
rect -633 928 -599 944
rect -633 -944 -599 -928
rect -325 928 -291 944
rect -325 -944 -291 -928
rect -17 928 17 944
rect -17 -944 17 -928
rect 291 928 325 944
rect 291 -944 325 -928
rect 599 928 633 944
rect 599 -944 633 -928
rect 907 928 941 944
rect 907 -944 941 -928
rect 1215 928 1249 944
rect 1215 -944 1249 -928
rect 1523 928 1557 944
rect 1523 -944 1557 -928
rect 1831 928 1865 944
rect 1831 -944 1865 -928
rect 2139 928 2173 944
rect 2139 -944 2173 -928
rect 2447 928 2481 944
rect 2447 -944 2481 -928
rect -2435 -1021 -2419 -987
rect -2201 -1021 -2185 -987
rect -2127 -1021 -2111 -987
rect -1893 -1021 -1877 -987
rect -1819 -1021 -1803 -987
rect -1585 -1021 -1569 -987
rect -1511 -1021 -1495 -987
rect -1277 -1021 -1261 -987
rect -1203 -1021 -1187 -987
rect -969 -1021 -953 -987
rect -895 -1021 -879 -987
rect -661 -1021 -645 -987
rect -587 -1021 -571 -987
rect -353 -1021 -337 -987
rect -279 -1021 -263 -987
rect -45 -1021 -29 -987
rect 29 -1021 45 -987
rect 263 -1021 279 -987
rect 337 -1021 353 -987
rect 571 -1021 587 -987
rect 645 -1021 661 -987
rect 879 -1021 895 -987
rect 953 -1021 969 -987
rect 1187 -1021 1203 -987
rect 1261 -1021 1277 -987
rect 1495 -1021 1511 -987
rect 1569 -1021 1585 -987
rect 1803 -1021 1819 -987
rect 1877 -1021 1893 -987
rect 2111 -1021 2127 -987
rect 2185 -1021 2201 -987
rect 2419 -1021 2435 -987
rect -2615 -1125 -2581 -1063
rect 2581 -1125 2615 -1063
rect -2615 -1159 -2519 -1125
rect 2519 -1159 2615 -1125
<< viali >>
rect -2419 987 -2201 1021
rect -2111 987 -1893 1021
rect -1803 987 -1585 1021
rect -1495 987 -1277 1021
rect -1187 987 -969 1021
rect -879 987 -661 1021
rect -571 987 -353 1021
rect -263 987 -45 1021
rect 45 987 263 1021
rect 353 987 571 1021
rect 661 987 879 1021
rect 969 987 1187 1021
rect 1277 987 1495 1021
rect 1585 987 1803 1021
rect 1893 987 2111 1021
rect 2201 987 2419 1021
rect -2481 -928 -2447 928
rect -2173 -928 -2139 928
rect -1865 -928 -1831 928
rect -1557 -928 -1523 928
rect -1249 -928 -1215 928
rect -941 -928 -907 928
rect -633 -928 -599 928
rect -325 -928 -291 928
rect -17 -928 17 928
rect 291 -928 325 928
rect 599 -928 633 928
rect 907 -928 941 928
rect 1215 -928 1249 928
rect 1523 -928 1557 928
rect 1831 -928 1865 928
rect 2139 -928 2173 928
rect 2447 -928 2481 928
rect -2419 -1021 -2201 -987
rect -2111 -1021 -1893 -987
rect -1803 -1021 -1585 -987
rect -1495 -1021 -1277 -987
rect -1187 -1021 -969 -987
rect -879 -1021 -661 -987
rect -571 -1021 -353 -987
rect -263 -1021 -45 -987
rect 45 -1021 263 -987
rect 353 -1021 571 -987
rect 661 -1021 879 -987
rect 969 -1021 1187 -987
rect 1277 -1021 1495 -987
rect 1585 -1021 1803 -987
rect 1893 -1021 2111 -987
rect 2201 -1021 2419 -987
<< metal1 >>
rect -2431 1021 -2189 1027
rect -2431 987 -2419 1021
rect -2201 987 -2189 1021
rect -2431 981 -2189 987
rect -2123 1021 -1881 1027
rect -2123 987 -2111 1021
rect -1893 987 -1881 1021
rect -2123 981 -1881 987
rect -1815 1021 -1573 1027
rect -1815 987 -1803 1021
rect -1585 987 -1573 1021
rect -1815 981 -1573 987
rect -1507 1021 -1265 1027
rect -1507 987 -1495 1021
rect -1277 987 -1265 1021
rect -1507 981 -1265 987
rect -1199 1021 -957 1027
rect -1199 987 -1187 1021
rect -969 987 -957 1021
rect -1199 981 -957 987
rect -891 1021 -649 1027
rect -891 987 -879 1021
rect -661 987 -649 1021
rect -891 981 -649 987
rect -583 1021 -341 1027
rect -583 987 -571 1021
rect -353 987 -341 1021
rect -583 981 -341 987
rect -275 1021 -33 1027
rect -275 987 -263 1021
rect -45 987 -33 1021
rect -275 981 -33 987
rect 33 1021 275 1027
rect 33 987 45 1021
rect 263 987 275 1021
rect 33 981 275 987
rect 341 1021 583 1027
rect 341 987 353 1021
rect 571 987 583 1021
rect 341 981 583 987
rect 649 1021 891 1027
rect 649 987 661 1021
rect 879 987 891 1021
rect 649 981 891 987
rect 957 1021 1199 1027
rect 957 987 969 1021
rect 1187 987 1199 1021
rect 957 981 1199 987
rect 1265 1021 1507 1027
rect 1265 987 1277 1021
rect 1495 987 1507 1021
rect 1265 981 1507 987
rect 1573 1021 1815 1027
rect 1573 987 1585 1021
rect 1803 987 1815 1021
rect 1573 981 1815 987
rect 1881 1021 2123 1027
rect 1881 987 1893 1021
rect 2111 987 2123 1021
rect 1881 981 2123 987
rect 2189 1021 2431 1027
rect 2189 987 2201 1021
rect 2419 987 2431 1021
rect 2189 981 2431 987
rect -2487 928 -2441 940
rect -2487 -928 -2481 928
rect -2447 -928 -2441 928
rect -2487 -940 -2441 -928
rect -2179 928 -2133 940
rect -2179 -928 -2173 928
rect -2139 -928 -2133 928
rect -2179 -940 -2133 -928
rect -1871 928 -1825 940
rect -1871 -928 -1865 928
rect -1831 -928 -1825 928
rect -1871 -940 -1825 -928
rect -1563 928 -1517 940
rect -1563 -928 -1557 928
rect -1523 -928 -1517 928
rect -1563 -940 -1517 -928
rect -1255 928 -1209 940
rect -1255 -928 -1249 928
rect -1215 -928 -1209 928
rect -1255 -940 -1209 -928
rect -947 928 -901 940
rect -947 -928 -941 928
rect -907 -928 -901 928
rect -947 -940 -901 -928
rect -639 928 -593 940
rect -639 -928 -633 928
rect -599 -928 -593 928
rect -639 -940 -593 -928
rect -331 928 -285 940
rect -331 -928 -325 928
rect -291 -928 -285 928
rect -331 -940 -285 -928
rect -23 928 23 940
rect -23 -928 -17 928
rect 17 -928 23 928
rect -23 -940 23 -928
rect 285 928 331 940
rect 285 -928 291 928
rect 325 -928 331 928
rect 285 -940 331 -928
rect 593 928 639 940
rect 593 -928 599 928
rect 633 -928 639 928
rect 593 -940 639 -928
rect 901 928 947 940
rect 901 -928 907 928
rect 941 -928 947 928
rect 901 -940 947 -928
rect 1209 928 1255 940
rect 1209 -928 1215 928
rect 1249 -928 1255 928
rect 1209 -940 1255 -928
rect 1517 928 1563 940
rect 1517 -928 1523 928
rect 1557 -928 1563 928
rect 1517 -940 1563 -928
rect 1825 928 1871 940
rect 1825 -928 1831 928
rect 1865 -928 1871 928
rect 1825 -940 1871 -928
rect 2133 928 2179 940
rect 2133 -928 2139 928
rect 2173 -928 2179 928
rect 2133 -940 2179 -928
rect 2441 928 2487 940
rect 2441 -928 2447 928
rect 2481 -928 2487 928
rect 2441 -940 2487 -928
rect -2431 -987 -2189 -981
rect -2431 -1021 -2419 -987
rect -2201 -1021 -2189 -987
rect -2431 -1027 -2189 -1021
rect -2123 -987 -1881 -981
rect -2123 -1021 -2111 -987
rect -1893 -1021 -1881 -987
rect -2123 -1027 -1881 -1021
rect -1815 -987 -1573 -981
rect -1815 -1021 -1803 -987
rect -1585 -1021 -1573 -987
rect -1815 -1027 -1573 -1021
rect -1507 -987 -1265 -981
rect -1507 -1021 -1495 -987
rect -1277 -1021 -1265 -987
rect -1507 -1027 -1265 -1021
rect -1199 -987 -957 -981
rect -1199 -1021 -1187 -987
rect -969 -1021 -957 -987
rect -1199 -1027 -957 -1021
rect -891 -987 -649 -981
rect -891 -1021 -879 -987
rect -661 -1021 -649 -987
rect -891 -1027 -649 -1021
rect -583 -987 -341 -981
rect -583 -1021 -571 -987
rect -353 -1021 -341 -987
rect -583 -1027 -341 -1021
rect -275 -987 -33 -981
rect -275 -1021 -263 -987
rect -45 -1021 -33 -987
rect -275 -1027 -33 -1021
rect 33 -987 275 -981
rect 33 -1021 45 -987
rect 263 -1021 275 -987
rect 33 -1027 275 -1021
rect 341 -987 583 -981
rect 341 -1021 353 -987
rect 571 -1021 583 -987
rect 341 -1027 583 -1021
rect 649 -987 891 -981
rect 649 -1021 661 -987
rect 879 -1021 891 -987
rect 649 -1027 891 -1021
rect 957 -987 1199 -981
rect 957 -1021 969 -987
rect 1187 -1021 1199 -987
rect 957 -1027 1199 -1021
rect 1265 -987 1507 -981
rect 1265 -1021 1277 -987
rect 1495 -1021 1507 -987
rect 1265 -1027 1507 -1021
rect 1573 -987 1815 -981
rect 1573 -1021 1585 -987
rect 1803 -1021 1815 -987
rect 1573 -1027 1815 -1021
rect 1881 -987 2123 -981
rect 1881 -1021 1893 -987
rect 2111 -1021 2123 -987
rect 1881 -1027 2123 -1021
rect 2189 -987 2431 -981
rect 2189 -1021 2201 -987
rect 2419 -1021 2431 -987
rect 2189 -1027 2431 -1021
<< properties >>
string FIXED_BBOX -2598 -1142 2598 1142
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9.4 l 1.25 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
