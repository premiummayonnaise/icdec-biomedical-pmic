magic
tech sky130A
magscale 1 2
timestamp 1770371891
<< nwell >>
rect 23396 -19582 30396 -18602
rect 20256 -22582 33536 -19582
rect 20256 -24322 22756 -22582
rect 20256 -28182 20536 -24322
rect 31036 -24322 33536 -22582
rect 33256 -28182 33536 -24322
rect 20256 -28462 23636 -28182
rect 23356 -29182 23636 -28462
rect 30116 -28462 33536 -28182
rect 30116 -29182 30396 -28462
rect 23356 -29462 30396 -29182
<< pwell >>
rect 22796 -24362 30996 -22622
rect 20556 -24382 33256 -24362
rect 20556 -26682 33236 -24382
rect 20556 -26702 31136 -26682
rect 32316 -26702 33236 -26682
rect 20556 -28162 33236 -26702
rect 23636 -29182 30116 -28182
<< mvnmos >>
rect 21474 -26254 21724 -24754
rect 21782 -26254 22032 -24754
rect 22090 -26254 22340 -24754
rect 22398 -26254 22648 -24754
rect 23414 -24094 23514 -23144
rect 23572 -24094 23672 -23144
rect 23854 -24094 23954 -23144
rect 24012 -24094 24112 -23144
rect 24294 -24094 24394 -23144
rect 24452 -24094 24552 -23144
rect 25214 -24094 25314 -23144
rect 25372 -24094 25472 -23144
rect 25654 -24094 25754 -23144
rect 25812 -24094 25912 -23144
rect 26094 -24094 26194 -23144
rect 26252 -24094 26352 -23144
rect 27414 -24094 27514 -23144
rect 27572 -24094 27672 -23144
rect 27854 -24094 27954 -23144
rect 28012 -24094 28112 -23144
rect 28294 -24094 28394 -23144
rect 28452 -24094 28552 -23144
rect 29214 -24094 29314 -23144
rect 29372 -24094 29472 -23144
rect 29654 -24094 29754 -23144
rect 29812 -24094 29912 -23144
rect 30094 -24094 30194 -23144
rect 30252 -24094 30352 -23144
rect 23414 -25796 23514 -24846
rect 23572 -25796 23672 -24846
rect 23854 -25796 23954 -24846
rect 24012 -25796 24112 -24846
rect 24294 -25796 24394 -24846
rect 24452 -25796 24552 -24846
rect 25214 -25796 25314 -24846
rect 25372 -25796 25472 -24846
rect 25654 -25796 25754 -24846
rect 25812 -25796 25912 -24846
rect 26094 -25796 26194 -24846
rect 26252 -25796 26352 -24846
rect 27414 -25796 27514 -24846
rect 27572 -25796 27672 -24846
rect 27854 -25796 27954 -24846
rect 28012 -25796 28112 -24846
rect 28294 -25796 28394 -24846
rect 28452 -25796 28552 -24846
rect 29214 -25796 29314 -24846
rect 29372 -25796 29472 -24846
rect 29654 -25796 29754 -24846
rect 29812 -25796 29912 -24846
rect 30094 -25796 30194 -24846
rect 30252 -25796 30352 -24846
rect 23994 -27896 24094 -26396
rect 24152 -27896 24252 -26396
rect 24434 -27896 24684 -26396
rect 24742 -27896 24992 -26396
rect 25050 -27896 25300 -26396
rect 25358 -27896 25608 -26396
rect 25666 -27896 25916 -26396
rect 25974 -27896 26224 -26396
rect 26282 -27896 26532 -26396
rect 26590 -27896 26840 -26396
rect 26898 -27896 27148 -26396
rect 27206 -27896 27456 -26396
rect 27514 -27896 27764 -26396
rect 27822 -27896 28072 -26396
rect 28130 -27896 28380 -26396
rect 28438 -27896 28688 -26396
rect 28746 -27896 28996 -26396
rect 29054 -27896 29304 -26396
rect 29494 -27896 29594 -26396
rect 29652 -27896 29752 -26396
rect 31134 -26274 31384 -24774
rect 31442 -26274 31692 -24774
rect 31750 -26274 32000 -24774
rect 32058 -26274 32308 -24774
<< mvpmos >>
rect 20960 -22222 21210 -20222
rect 21268 -22222 21518 -20222
rect 21576 -22222 21826 -20222
rect 21884 -22222 22134 -20222
rect 22192 -22222 22442 -20222
rect 22500 -22222 22750 -20222
rect 22808 -22222 23058 -20222
rect 23116 -22222 23366 -20222
rect 23960 -21742 24060 -19862
rect 24118 -21742 24218 -19862
rect 24395 -21747 24645 -19867
rect 24703 -21747 24953 -19867
rect 25011 -21747 25261 -19867
rect 25319 -21747 25569 -19867
rect 25627 -21747 25877 -19867
rect 25935 -21747 26185 -19867
rect 26243 -21747 26493 -19867
rect 26551 -21747 26801 -19867
rect 26859 -21747 27109 -19867
rect 27167 -21747 27417 -19867
rect 27475 -21747 27725 -19867
rect 27783 -21747 28033 -19867
rect 28091 -21747 28341 -19867
rect 28399 -21747 28649 -19867
rect 28707 -21747 28957 -19867
rect 29015 -21747 29265 -19867
rect 29500 -21742 29600 -19862
rect 29658 -21742 29758 -19862
rect 30400 -22222 30650 -20222
rect 30708 -22222 30958 -20222
rect 31016 -22222 31266 -20222
rect 31324 -22222 31574 -20222
rect 31632 -22222 31882 -20222
rect 31940 -22222 32190 -20222
rect 32248 -22222 32498 -20222
rect 32556 -22222 32806 -20222
rect 21920 -23922 22100 -22922
rect 22158 -23922 22338 -22922
rect 31500 -23902 31680 -22902
rect 31738 -23902 31918 -22902
<< mvndiff >>
rect 21416 -24766 21474 -24754
rect 21416 -26242 21428 -24766
rect 21462 -26242 21474 -24766
rect 21416 -26254 21474 -26242
rect 21724 -24766 21782 -24754
rect 21724 -26242 21736 -24766
rect 21770 -26242 21782 -24766
rect 21724 -26254 21782 -26242
rect 22032 -24766 22090 -24754
rect 22032 -26242 22044 -24766
rect 22078 -26242 22090 -24766
rect 22032 -26254 22090 -26242
rect 22340 -24766 22398 -24754
rect 22340 -26242 22352 -24766
rect 22386 -26242 22398 -24766
rect 22340 -26254 22398 -26242
rect 22648 -24766 22706 -24754
rect 22648 -26242 22660 -24766
rect 22694 -26242 22706 -24766
rect 22648 -26254 22706 -26242
rect 23356 -23156 23414 -23144
rect 23356 -24082 23368 -23156
rect 23402 -24082 23414 -23156
rect 23356 -24094 23414 -24082
rect 23514 -23156 23572 -23144
rect 23514 -24082 23526 -23156
rect 23560 -24082 23572 -23156
rect 23514 -24094 23572 -24082
rect 23672 -23156 23730 -23144
rect 23672 -24082 23684 -23156
rect 23718 -24082 23730 -23156
rect 23672 -24094 23730 -24082
rect 23796 -23156 23854 -23144
rect 23796 -24082 23808 -23156
rect 23842 -24082 23854 -23156
rect 23796 -24094 23854 -24082
rect 23954 -23156 24012 -23144
rect 23954 -24082 23966 -23156
rect 24000 -24082 24012 -23156
rect 23954 -24094 24012 -24082
rect 24112 -23156 24170 -23144
rect 24112 -24082 24124 -23156
rect 24158 -24082 24170 -23156
rect 24112 -24094 24170 -24082
rect 24236 -23156 24294 -23144
rect 24236 -24082 24248 -23156
rect 24282 -24082 24294 -23156
rect 24236 -24094 24294 -24082
rect 24394 -23156 24452 -23144
rect 24394 -24082 24406 -23156
rect 24440 -24082 24452 -23156
rect 24394 -24094 24452 -24082
rect 24552 -23156 24610 -23144
rect 24552 -24082 24564 -23156
rect 24598 -24082 24610 -23156
rect 24552 -24094 24610 -24082
rect 25156 -23156 25214 -23144
rect 25156 -24082 25168 -23156
rect 25202 -24082 25214 -23156
rect 25156 -24094 25214 -24082
rect 25314 -23156 25372 -23144
rect 25314 -24082 25326 -23156
rect 25360 -24082 25372 -23156
rect 25314 -24094 25372 -24082
rect 25472 -23156 25530 -23144
rect 25472 -24082 25484 -23156
rect 25518 -24082 25530 -23156
rect 25472 -24094 25530 -24082
rect 25596 -23156 25654 -23144
rect 25596 -24082 25608 -23156
rect 25642 -24082 25654 -23156
rect 25596 -24094 25654 -24082
rect 25754 -23156 25812 -23144
rect 25754 -24082 25766 -23156
rect 25800 -24082 25812 -23156
rect 25754 -24094 25812 -24082
rect 25912 -23156 25970 -23144
rect 25912 -24082 25924 -23156
rect 25958 -24082 25970 -23156
rect 25912 -24094 25970 -24082
rect 26036 -23156 26094 -23144
rect 26036 -24082 26048 -23156
rect 26082 -24082 26094 -23156
rect 26036 -24094 26094 -24082
rect 26194 -23156 26252 -23144
rect 26194 -24082 26206 -23156
rect 26240 -24082 26252 -23156
rect 26194 -24094 26252 -24082
rect 26352 -23156 26410 -23144
rect 26352 -24082 26364 -23156
rect 26398 -24082 26410 -23156
rect 26352 -24094 26410 -24082
rect 27356 -23156 27414 -23144
rect 27356 -24082 27368 -23156
rect 27402 -24082 27414 -23156
rect 27356 -24094 27414 -24082
rect 27514 -23156 27572 -23144
rect 27514 -24082 27526 -23156
rect 27560 -24082 27572 -23156
rect 27514 -24094 27572 -24082
rect 27672 -23156 27730 -23144
rect 27672 -24082 27684 -23156
rect 27718 -24082 27730 -23156
rect 27672 -24094 27730 -24082
rect 27796 -23156 27854 -23144
rect 27796 -24082 27808 -23156
rect 27842 -24082 27854 -23156
rect 27796 -24094 27854 -24082
rect 27954 -23156 28012 -23144
rect 27954 -24082 27966 -23156
rect 28000 -24082 28012 -23156
rect 27954 -24094 28012 -24082
rect 28112 -23156 28170 -23144
rect 28112 -24082 28124 -23156
rect 28158 -24082 28170 -23156
rect 28112 -24094 28170 -24082
rect 28236 -23156 28294 -23144
rect 28236 -24082 28248 -23156
rect 28282 -24082 28294 -23156
rect 28236 -24094 28294 -24082
rect 28394 -23156 28452 -23144
rect 28394 -24082 28406 -23156
rect 28440 -24082 28452 -23156
rect 28394 -24094 28452 -24082
rect 28552 -23156 28610 -23144
rect 28552 -24082 28564 -23156
rect 28598 -24082 28610 -23156
rect 28552 -24094 28610 -24082
rect 29156 -23156 29214 -23144
rect 29156 -24082 29168 -23156
rect 29202 -24082 29214 -23156
rect 29156 -24094 29214 -24082
rect 29314 -23156 29372 -23144
rect 29314 -24082 29326 -23156
rect 29360 -24082 29372 -23156
rect 29314 -24094 29372 -24082
rect 29472 -23156 29530 -23144
rect 29472 -24082 29484 -23156
rect 29518 -24082 29530 -23156
rect 29472 -24094 29530 -24082
rect 29596 -23156 29654 -23144
rect 29596 -24082 29608 -23156
rect 29642 -24082 29654 -23156
rect 29596 -24094 29654 -24082
rect 29754 -23156 29812 -23144
rect 29754 -24082 29766 -23156
rect 29800 -24082 29812 -23156
rect 29754 -24094 29812 -24082
rect 29912 -23156 29970 -23144
rect 29912 -24082 29924 -23156
rect 29958 -24082 29970 -23156
rect 29912 -24094 29970 -24082
rect 30036 -23156 30094 -23144
rect 30036 -24082 30048 -23156
rect 30082 -24082 30094 -23156
rect 30036 -24094 30094 -24082
rect 30194 -23156 30252 -23144
rect 30194 -24082 30206 -23156
rect 30240 -24082 30252 -23156
rect 30194 -24094 30252 -24082
rect 30352 -23156 30410 -23144
rect 30352 -24082 30364 -23156
rect 30398 -24082 30410 -23156
rect 30352 -24094 30410 -24082
rect 23356 -24858 23414 -24846
rect 23356 -25784 23368 -24858
rect 23402 -25784 23414 -24858
rect 23356 -25796 23414 -25784
rect 23514 -24858 23572 -24846
rect 23514 -25784 23526 -24858
rect 23560 -25784 23572 -24858
rect 23514 -25796 23572 -25784
rect 23672 -24858 23730 -24846
rect 23672 -25784 23684 -24858
rect 23718 -25784 23730 -24858
rect 23672 -25796 23730 -25784
rect 23796 -24858 23854 -24846
rect 23796 -25784 23808 -24858
rect 23842 -25784 23854 -24858
rect 23796 -25796 23854 -25784
rect 23954 -24858 24012 -24846
rect 23954 -25784 23966 -24858
rect 24000 -25784 24012 -24858
rect 23954 -25796 24012 -25784
rect 24112 -24858 24170 -24846
rect 24112 -25784 24124 -24858
rect 24158 -25784 24170 -24858
rect 24112 -25796 24170 -25784
rect 24236 -24858 24294 -24846
rect 24236 -25784 24248 -24858
rect 24282 -25784 24294 -24858
rect 24236 -25796 24294 -25784
rect 24394 -24858 24452 -24846
rect 24394 -25784 24406 -24858
rect 24440 -25784 24452 -24858
rect 24394 -25796 24452 -25784
rect 24552 -24858 24610 -24846
rect 24552 -25784 24564 -24858
rect 24598 -25784 24610 -24858
rect 24552 -25796 24610 -25784
rect 25156 -24858 25214 -24846
rect 25156 -25784 25168 -24858
rect 25202 -25784 25214 -24858
rect 25156 -25796 25214 -25784
rect 25314 -24858 25372 -24846
rect 25314 -25784 25326 -24858
rect 25360 -25784 25372 -24858
rect 25314 -25796 25372 -25784
rect 25472 -24858 25530 -24846
rect 25472 -25784 25484 -24858
rect 25518 -25784 25530 -24858
rect 25472 -25796 25530 -25784
rect 25596 -24858 25654 -24846
rect 25596 -25784 25608 -24858
rect 25642 -25784 25654 -24858
rect 25596 -25796 25654 -25784
rect 25754 -24858 25812 -24846
rect 25754 -25784 25766 -24858
rect 25800 -25784 25812 -24858
rect 25754 -25796 25812 -25784
rect 25912 -24858 25970 -24846
rect 25912 -25784 25924 -24858
rect 25958 -25784 25970 -24858
rect 25912 -25796 25970 -25784
rect 26036 -24858 26094 -24846
rect 26036 -25784 26048 -24858
rect 26082 -25784 26094 -24858
rect 26036 -25796 26094 -25784
rect 26194 -24858 26252 -24846
rect 26194 -25784 26206 -24858
rect 26240 -25784 26252 -24858
rect 26194 -25796 26252 -25784
rect 26352 -24858 26410 -24846
rect 26352 -25784 26364 -24858
rect 26398 -25784 26410 -24858
rect 26352 -25796 26410 -25784
rect 27356 -24858 27414 -24846
rect 27356 -25784 27368 -24858
rect 27402 -25784 27414 -24858
rect 27356 -25796 27414 -25784
rect 27514 -24858 27572 -24846
rect 27514 -25784 27526 -24858
rect 27560 -25784 27572 -24858
rect 27514 -25796 27572 -25784
rect 27672 -24858 27730 -24846
rect 27672 -25784 27684 -24858
rect 27718 -25784 27730 -24858
rect 27672 -25796 27730 -25784
rect 27796 -24858 27854 -24846
rect 27796 -25784 27808 -24858
rect 27842 -25784 27854 -24858
rect 27796 -25796 27854 -25784
rect 27954 -24858 28012 -24846
rect 27954 -25784 27966 -24858
rect 28000 -25784 28012 -24858
rect 27954 -25796 28012 -25784
rect 28112 -24858 28170 -24846
rect 28112 -25784 28124 -24858
rect 28158 -25784 28170 -24858
rect 28112 -25796 28170 -25784
rect 28236 -24858 28294 -24846
rect 28236 -25784 28248 -24858
rect 28282 -25784 28294 -24858
rect 28236 -25796 28294 -25784
rect 28394 -24858 28452 -24846
rect 28394 -25784 28406 -24858
rect 28440 -25784 28452 -24858
rect 28394 -25796 28452 -25784
rect 28552 -24858 28610 -24846
rect 28552 -25784 28564 -24858
rect 28598 -25784 28610 -24858
rect 28552 -25796 28610 -25784
rect 29156 -24858 29214 -24846
rect 29156 -25784 29168 -24858
rect 29202 -25784 29214 -24858
rect 29156 -25796 29214 -25784
rect 29314 -24858 29372 -24846
rect 29314 -25784 29326 -24858
rect 29360 -25784 29372 -24858
rect 29314 -25796 29372 -25784
rect 29472 -24858 29530 -24846
rect 29472 -25784 29484 -24858
rect 29518 -25784 29530 -24858
rect 29472 -25796 29530 -25784
rect 29596 -24858 29654 -24846
rect 29596 -25784 29608 -24858
rect 29642 -25784 29654 -24858
rect 29596 -25796 29654 -25784
rect 29754 -24858 29812 -24846
rect 29754 -25784 29766 -24858
rect 29800 -25784 29812 -24858
rect 29754 -25796 29812 -25784
rect 29912 -24858 29970 -24846
rect 29912 -25784 29924 -24858
rect 29958 -25784 29970 -24858
rect 29912 -25796 29970 -25784
rect 30036 -24858 30094 -24846
rect 30036 -25784 30048 -24858
rect 30082 -25784 30094 -24858
rect 30036 -25796 30094 -25784
rect 30194 -24858 30252 -24846
rect 30194 -25784 30206 -24858
rect 30240 -25784 30252 -24858
rect 30194 -25796 30252 -25784
rect 30352 -24858 30410 -24846
rect 30352 -25784 30364 -24858
rect 30398 -25784 30410 -24858
rect 30352 -25796 30410 -25784
rect 23936 -26408 23994 -26396
rect 23936 -27884 23948 -26408
rect 23982 -27884 23994 -26408
rect 23936 -27896 23994 -27884
rect 24094 -26408 24152 -26396
rect 24094 -27884 24106 -26408
rect 24140 -27884 24152 -26408
rect 24094 -27896 24152 -27884
rect 24252 -26408 24310 -26396
rect 24252 -27884 24264 -26408
rect 24298 -27884 24310 -26408
rect 24252 -27896 24310 -27884
rect 24376 -26408 24434 -26396
rect 24376 -27884 24388 -26408
rect 24422 -27884 24434 -26408
rect 24376 -27896 24434 -27884
rect 24684 -26408 24742 -26396
rect 24684 -27884 24696 -26408
rect 24730 -27884 24742 -26408
rect 24684 -27896 24742 -27884
rect 24992 -26408 25050 -26396
rect 24992 -27884 25004 -26408
rect 25038 -27884 25050 -26408
rect 24992 -27896 25050 -27884
rect 25300 -26408 25358 -26396
rect 25300 -27884 25312 -26408
rect 25346 -27884 25358 -26408
rect 25300 -27896 25358 -27884
rect 25608 -26408 25666 -26396
rect 25608 -27884 25620 -26408
rect 25654 -27884 25666 -26408
rect 25608 -27896 25666 -27884
rect 25916 -26408 25974 -26396
rect 25916 -27884 25928 -26408
rect 25962 -27884 25974 -26408
rect 25916 -27896 25974 -27884
rect 26224 -26408 26282 -26396
rect 26224 -27884 26236 -26408
rect 26270 -27884 26282 -26408
rect 26224 -27896 26282 -27884
rect 26532 -26408 26590 -26396
rect 26532 -27884 26544 -26408
rect 26578 -27884 26590 -26408
rect 26532 -27896 26590 -27884
rect 26840 -26408 26898 -26396
rect 26840 -27884 26852 -26408
rect 26886 -27884 26898 -26408
rect 26840 -27896 26898 -27884
rect 27148 -26408 27206 -26396
rect 27148 -27884 27160 -26408
rect 27194 -27884 27206 -26408
rect 27148 -27896 27206 -27884
rect 27456 -26408 27514 -26396
rect 27456 -27884 27468 -26408
rect 27502 -27884 27514 -26408
rect 27456 -27896 27514 -27884
rect 27764 -26408 27822 -26396
rect 27764 -27884 27776 -26408
rect 27810 -27884 27822 -26408
rect 27764 -27896 27822 -27884
rect 28072 -26408 28130 -26396
rect 28072 -27884 28084 -26408
rect 28118 -27884 28130 -26408
rect 28072 -27896 28130 -27884
rect 28380 -26408 28438 -26396
rect 28380 -27884 28392 -26408
rect 28426 -27884 28438 -26408
rect 28380 -27896 28438 -27884
rect 28688 -26408 28746 -26396
rect 28688 -27884 28700 -26408
rect 28734 -27884 28746 -26408
rect 28688 -27896 28746 -27884
rect 28996 -26408 29054 -26396
rect 28996 -27884 29008 -26408
rect 29042 -27884 29054 -26408
rect 28996 -27896 29054 -27884
rect 29304 -26408 29362 -26396
rect 29304 -27884 29316 -26408
rect 29350 -27884 29362 -26408
rect 29304 -27896 29362 -27884
rect 29436 -26408 29494 -26396
rect 29436 -27884 29448 -26408
rect 29482 -27884 29494 -26408
rect 29436 -27896 29494 -27884
rect 29594 -26408 29652 -26396
rect 29594 -27884 29606 -26408
rect 29640 -27884 29652 -26408
rect 29594 -27896 29652 -27884
rect 29752 -26408 29810 -26396
rect 29752 -27884 29764 -26408
rect 29798 -27884 29810 -26408
rect 29752 -27896 29810 -27884
rect 31076 -24786 31134 -24774
rect 31076 -26262 31088 -24786
rect 31122 -26262 31134 -24786
rect 31076 -26274 31134 -26262
rect 31384 -24786 31442 -24774
rect 31384 -26262 31396 -24786
rect 31430 -26262 31442 -24786
rect 31384 -26274 31442 -26262
rect 31692 -24786 31750 -24774
rect 31692 -26262 31704 -24786
rect 31738 -26262 31750 -24786
rect 31692 -26274 31750 -26262
rect 32000 -24786 32058 -24774
rect 32000 -26262 32012 -24786
rect 32046 -26262 32058 -24786
rect 32000 -26274 32058 -26262
rect 32308 -24786 32366 -24774
rect 32308 -26262 32320 -24786
rect 32354 -26262 32366 -24786
rect 32308 -26274 32366 -26262
<< mvpdiff >>
rect 20902 -20234 20960 -20222
rect 20902 -22210 20914 -20234
rect 20948 -22210 20960 -20234
rect 20902 -22222 20960 -22210
rect 21210 -20234 21268 -20222
rect 21210 -22210 21222 -20234
rect 21256 -22210 21268 -20234
rect 21210 -22222 21268 -22210
rect 21518 -20234 21576 -20222
rect 21518 -22210 21530 -20234
rect 21564 -22210 21576 -20234
rect 21518 -22222 21576 -22210
rect 21826 -20234 21884 -20222
rect 21826 -22210 21838 -20234
rect 21872 -22210 21884 -20234
rect 21826 -22222 21884 -22210
rect 22134 -20234 22192 -20222
rect 22134 -22210 22146 -20234
rect 22180 -22210 22192 -20234
rect 22134 -22222 22192 -22210
rect 22442 -20234 22500 -20222
rect 22442 -22210 22454 -20234
rect 22488 -22210 22500 -20234
rect 22442 -22222 22500 -22210
rect 22750 -20234 22808 -20222
rect 22750 -22210 22762 -20234
rect 22796 -22210 22808 -20234
rect 22750 -22222 22808 -22210
rect 23058 -20234 23116 -20222
rect 23058 -22210 23070 -20234
rect 23104 -22210 23116 -20234
rect 23058 -22222 23116 -22210
rect 23366 -20234 23424 -20222
rect 23366 -22210 23378 -20234
rect 23412 -22210 23424 -20234
rect 23366 -22222 23424 -22210
rect 23902 -19874 23960 -19862
rect 23902 -21730 23914 -19874
rect 23948 -21730 23960 -19874
rect 23902 -21742 23960 -21730
rect 24060 -19874 24118 -19862
rect 24060 -21730 24072 -19874
rect 24106 -21730 24118 -19874
rect 24060 -21742 24118 -21730
rect 24218 -19874 24276 -19862
rect 24218 -21730 24230 -19874
rect 24264 -21730 24276 -19874
rect 24218 -21742 24276 -21730
rect 24337 -20065 24395 -19867
rect 24337 -21549 24349 -20065
rect 24383 -21549 24395 -20065
rect 24337 -21747 24395 -21549
rect 24645 -20065 24703 -19867
rect 24645 -21549 24657 -20065
rect 24691 -21549 24703 -20065
rect 24645 -21747 24703 -21549
rect 24953 -20065 25011 -19867
rect 24953 -21549 24965 -20065
rect 24999 -21549 25011 -20065
rect 24953 -21747 25011 -21549
rect 25261 -20065 25319 -19867
rect 25261 -21549 25273 -20065
rect 25307 -21549 25319 -20065
rect 25261 -21747 25319 -21549
rect 25569 -20065 25627 -19867
rect 25569 -21549 25581 -20065
rect 25615 -21549 25627 -20065
rect 25569 -21747 25627 -21549
rect 25877 -20065 25935 -19867
rect 25877 -21549 25889 -20065
rect 25923 -21549 25935 -20065
rect 25877 -21747 25935 -21549
rect 26185 -20065 26243 -19867
rect 26185 -21549 26197 -20065
rect 26231 -21549 26243 -20065
rect 26185 -21747 26243 -21549
rect 26493 -20065 26551 -19867
rect 26493 -21549 26505 -20065
rect 26539 -21549 26551 -20065
rect 26493 -21747 26551 -21549
rect 26801 -20065 26859 -19867
rect 26801 -21549 26813 -20065
rect 26847 -21549 26859 -20065
rect 26801 -21747 26859 -21549
rect 27109 -20065 27167 -19867
rect 27109 -21549 27121 -20065
rect 27155 -21549 27167 -20065
rect 27109 -21747 27167 -21549
rect 27417 -20065 27475 -19867
rect 27417 -21549 27429 -20065
rect 27463 -21549 27475 -20065
rect 27417 -21747 27475 -21549
rect 27725 -20065 27783 -19867
rect 27725 -21549 27737 -20065
rect 27771 -21549 27783 -20065
rect 27725 -21747 27783 -21549
rect 28033 -20065 28091 -19867
rect 28033 -21549 28045 -20065
rect 28079 -21549 28091 -20065
rect 28033 -21747 28091 -21549
rect 28341 -20065 28399 -19867
rect 28341 -21549 28353 -20065
rect 28387 -21549 28399 -20065
rect 28341 -21747 28399 -21549
rect 28649 -20065 28707 -19867
rect 28649 -21549 28661 -20065
rect 28695 -21549 28707 -20065
rect 28649 -21747 28707 -21549
rect 28957 -20065 29015 -19867
rect 28957 -21549 28969 -20065
rect 29003 -21549 29015 -20065
rect 28957 -21747 29015 -21549
rect 29265 -20065 29323 -19867
rect 29265 -21549 29277 -20065
rect 29311 -21549 29323 -20065
rect 29265 -21747 29323 -21549
rect 29442 -19874 29500 -19862
rect 29442 -21730 29454 -19874
rect 29488 -21730 29500 -19874
rect 29442 -21742 29500 -21730
rect 29600 -19874 29658 -19862
rect 29600 -21730 29612 -19874
rect 29646 -21730 29658 -19874
rect 29600 -21742 29658 -21730
rect 29758 -19874 29816 -19862
rect 29758 -21730 29770 -19874
rect 29804 -21730 29816 -19874
rect 29758 -21742 29816 -21730
rect 30342 -20234 30400 -20222
rect 30342 -22210 30354 -20234
rect 30388 -22210 30400 -20234
rect 30342 -22222 30400 -22210
rect 30650 -20234 30708 -20222
rect 30650 -22210 30662 -20234
rect 30696 -22210 30708 -20234
rect 30650 -22222 30708 -22210
rect 30958 -20234 31016 -20222
rect 30958 -22210 30970 -20234
rect 31004 -22210 31016 -20234
rect 30958 -22222 31016 -22210
rect 31266 -20234 31324 -20222
rect 31266 -22210 31278 -20234
rect 31312 -22210 31324 -20234
rect 31266 -22222 31324 -22210
rect 31574 -20234 31632 -20222
rect 31574 -22210 31586 -20234
rect 31620 -22210 31632 -20234
rect 31574 -22222 31632 -22210
rect 31882 -20234 31940 -20222
rect 31882 -22210 31894 -20234
rect 31928 -22210 31940 -20234
rect 31882 -22222 31940 -22210
rect 32190 -20234 32248 -20222
rect 32190 -22210 32202 -20234
rect 32236 -22210 32248 -20234
rect 32190 -22222 32248 -22210
rect 32498 -20234 32556 -20222
rect 32498 -22210 32510 -20234
rect 32544 -22210 32556 -20234
rect 32498 -22222 32556 -22210
rect 32806 -20234 32864 -20222
rect 32806 -22210 32818 -20234
rect 32852 -22210 32864 -20234
rect 32806 -22222 32864 -22210
rect 21862 -22934 21920 -22922
rect 21862 -23910 21874 -22934
rect 21908 -23910 21920 -22934
rect 21862 -23922 21920 -23910
rect 22100 -22934 22158 -22922
rect 22100 -23910 22112 -22934
rect 22146 -23910 22158 -22934
rect 22100 -23922 22158 -23910
rect 22338 -22934 22396 -22922
rect 22338 -23910 22350 -22934
rect 22384 -23910 22396 -22934
rect 22338 -23922 22396 -23910
rect 31442 -22914 31500 -22902
rect 31442 -23890 31454 -22914
rect 31488 -23890 31500 -22914
rect 31442 -23902 31500 -23890
rect 31680 -22914 31738 -22902
rect 31680 -23890 31692 -22914
rect 31726 -23890 31738 -22914
rect 31680 -23902 31738 -23890
rect 31918 -22914 31976 -22902
rect 31918 -23890 31930 -22914
rect 31964 -23890 31976 -22914
rect 31918 -23902 31976 -23890
<< mvndiffc >>
rect 21428 -26242 21462 -24766
rect 21736 -26242 21770 -24766
rect 22044 -26242 22078 -24766
rect 22352 -26242 22386 -24766
rect 22660 -26242 22694 -24766
rect 23368 -24082 23402 -23156
rect 23526 -24082 23560 -23156
rect 23684 -24082 23718 -23156
rect 23808 -24082 23842 -23156
rect 23966 -24082 24000 -23156
rect 24124 -24082 24158 -23156
rect 24248 -24082 24282 -23156
rect 24406 -24082 24440 -23156
rect 24564 -24082 24598 -23156
rect 25168 -24082 25202 -23156
rect 25326 -24082 25360 -23156
rect 25484 -24082 25518 -23156
rect 25608 -24082 25642 -23156
rect 25766 -24082 25800 -23156
rect 25924 -24082 25958 -23156
rect 26048 -24082 26082 -23156
rect 26206 -24082 26240 -23156
rect 26364 -24082 26398 -23156
rect 27368 -24082 27402 -23156
rect 27526 -24082 27560 -23156
rect 27684 -24082 27718 -23156
rect 27808 -24082 27842 -23156
rect 27966 -24082 28000 -23156
rect 28124 -24082 28158 -23156
rect 28248 -24082 28282 -23156
rect 28406 -24082 28440 -23156
rect 28564 -24082 28598 -23156
rect 29168 -24082 29202 -23156
rect 29326 -24082 29360 -23156
rect 29484 -24082 29518 -23156
rect 29608 -24082 29642 -23156
rect 29766 -24082 29800 -23156
rect 29924 -24082 29958 -23156
rect 30048 -24082 30082 -23156
rect 30206 -24082 30240 -23156
rect 30364 -24082 30398 -23156
rect 23368 -25784 23402 -24858
rect 23526 -25784 23560 -24858
rect 23684 -25784 23718 -24858
rect 23808 -25784 23842 -24858
rect 23966 -25784 24000 -24858
rect 24124 -25784 24158 -24858
rect 24248 -25784 24282 -24858
rect 24406 -25784 24440 -24858
rect 24564 -25784 24598 -24858
rect 25168 -25784 25202 -24858
rect 25326 -25784 25360 -24858
rect 25484 -25784 25518 -24858
rect 25608 -25784 25642 -24858
rect 25766 -25784 25800 -24858
rect 25924 -25784 25958 -24858
rect 26048 -25784 26082 -24858
rect 26206 -25784 26240 -24858
rect 26364 -25784 26398 -24858
rect 27368 -25784 27402 -24858
rect 27526 -25784 27560 -24858
rect 27684 -25784 27718 -24858
rect 27808 -25784 27842 -24858
rect 27966 -25784 28000 -24858
rect 28124 -25784 28158 -24858
rect 28248 -25784 28282 -24858
rect 28406 -25784 28440 -24858
rect 28564 -25784 28598 -24858
rect 29168 -25784 29202 -24858
rect 29326 -25784 29360 -24858
rect 29484 -25784 29518 -24858
rect 29608 -25784 29642 -24858
rect 29766 -25784 29800 -24858
rect 29924 -25784 29958 -24858
rect 30048 -25784 30082 -24858
rect 30206 -25784 30240 -24858
rect 30364 -25784 30398 -24858
rect 23948 -27884 23982 -26408
rect 24106 -27884 24140 -26408
rect 24264 -27884 24298 -26408
rect 24388 -27884 24422 -26408
rect 24696 -27884 24730 -26408
rect 25004 -27884 25038 -26408
rect 25312 -27884 25346 -26408
rect 25620 -27884 25654 -26408
rect 25928 -27884 25962 -26408
rect 26236 -27884 26270 -26408
rect 26544 -27884 26578 -26408
rect 26852 -27884 26886 -26408
rect 27160 -27884 27194 -26408
rect 27468 -27884 27502 -26408
rect 27776 -27884 27810 -26408
rect 28084 -27884 28118 -26408
rect 28392 -27884 28426 -26408
rect 28700 -27884 28734 -26408
rect 29008 -27884 29042 -26408
rect 29316 -27884 29350 -26408
rect 29448 -27884 29482 -26408
rect 29606 -27884 29640 -26408
rect 29764 -27884 29798 -26408
rect 31088 -26262 31122 -24786
rect 31396 -26262 31430 -24786
rect 31704 -26262 31738 -24786
rect 32012 -26262 32046 -24786
rect 32320 -26262 32354 -24786
<< mvpdiffc >>
rect 20914 -22210 20948 -20234
rect 21222 -22210 21256 -20234
rect 21530 -22210 21564 -20234
rect 21838 -22210 21872 -20234
rect 22146 -22210 22180 -20234
rect 22454 -22210 22488 -20234
rect 22762 -22210 22796 -20234
rect 23070 -22210 23104 -20234
rect 23378 -22210 23412 -20234
rect 23914 -21730 23948 -19874
rect 24072 -21730 24106 -19874
rect 24230 -21730 24264 -19874
rect 24349 -21549 24383 -20065
rect 24657 -21549 24691 -20065
rect 24965 -21549 24999 -20065
rect 25273 -21549 25307 -20065
rect 25581 -21549 25615 -20065
rect 25889 -21549 25923 -20065
rect 26197 -21549 26231 -20065
rect 26505 -21549 26539 -20065
rect 26813 -21549 26847 -20065
rect 27121 -21549 27155 -20065
rect 27429 -21549 27463 -20065
rect 27737 -21549 27771 -20065
rect 28045 -21549 28079 -20065
rect 28353 -21549 28387 -20065
rect 28661 -21549 28695 -20065
rect 28969 -21549 29003 -20065
rect 29277 -21549 29311 -20065
rect 29454 -21730 29488 -19874
rect 29612 -21730 29646 -19874
rect 29770 -21730 29804 -19874
rect 30354 -22210 30388 -20234
rect 30662 -22210 30696 -20234
rect 30970 -22210 31004 -20234
rect 31278 -22210 31312 -20234
rect 31586 -22210 31620 -20234
rect 31894 -22210 31928 -20234
rect 32202 -22210 32236 -20234
rect 32510 -22210 32544 -20234
rect 32818 -22210 32852 -20234
rect 21874 -23910 21908 -22934
rect 22112 -23910 22146 -22934
rect 22350 -23910 22384 -22934
rect 31454 -23890 31488 -22914
rect 31692 -23890 31726 -22914
rect 31930 -23890 31964 -22914
<< psubdiff >>
rect 22996 -22742 30796 -22722
rect 22996 -22802 23116 -22742
rect 30676 -22802 30796 -22742
rect 22996 -22822 30796 -22802
rect 22996 -22842 23096 -22822
rect 21216 -24562 22916 -24542
rect 21216 -24622 21336 -24562
rect 22796 -24622 22916 -24562
rect 21216 -24642 22916 -24622
rect 21216 -24662 21316 -24642
rect 21216 -26422 21236 -24662
rect 21296 -26422 21316 -24662
rect 22816 -24662 22916 -24642
rect 21216 -26442 21316 -26422
rect 22816 -26422 22836 -24662
rect 22896 -26422 22916 -24662
rect 22996 -26102 23016 -22842
rect 23076 -26102 23096 -22842
rect 30696 -22842 30796 -22822
rect 23196 -22942 24796 -22922
rect 23196 -23002 23236 -22942
rect 24756 -23002 24796 -22942
rect 23196 -23022 24796 -23002
rect 23196 -24222 23296 -23022
rect 24696 -24222 24796 -23022
rect 23196 -24322 24796 -24222
rect 24996 -22942 26596 -22922
rect 24996 -23002 25036 -22942
rect 26556 -23002 26596 -22942
rect 24996 -23022 26596 -23002
rect 24996 -24222 25096 -23022
rect 26496 -24222 26596 -23022
rect 24996 -24322 26596 -24222
rect 27196 -22942 28796 -22922
rect 27196 -23002 27236 -22942
rect 28756 -23002 28796 -22942
rect 27196 -23022 28796 -23002
rect 27196 -24222 27296 -23022
rect 28696 -24222 28796 -23022
rect 27196 -24322 28796 -24222
rect 28996 -22942 30596 -22922
rect 28996 -23002 29036 -22942
rect 30556 -23002 30596 -22942
rect 28996 -23022 30596 -23002
rect 28996 -24222 29096 -23022
rect 30496 -24222 30596 -23022
rect 28996 -24322 30596 -24222
rect 23196 -24722 24796 -24622
rect 23196 -25922 23296 -24722
rect 24696 -25922 24796 -24722
rect 23196 -25942 24796 -25922
rect 23196 -26002 23236 -25942
rect 24756 -26002 24796 -25942
rect 23196 -26022 24796 -26002
rect 24996 -24722 26596 -24622
rect 24996 -25922 25096 -24722
rect 26496 -25922 26596 -24722
rect 24996 -25942 26596 -25922
rect 24996 -26002 25036 -25942
rect 26556 -26002 26596 -25942
rect 24996 -26022 26596 -26002
rect 27196 -24722 28796 -24622
rect 27196 -25922 27296 -24722
rect 28696 -25922 28796 -24722
rect 27196 -25942 28796 -25922
rect 27196 -26002 27236 -25942
rect 28756 -26002 28796 -25942
rect 27196 -26022 28796 -26002
rect 28996 -24722 30596 -24622
rect 28996 -25922 29096 -24722
rect 30496 -25922 30596 -24722
rect 28996 -25942 30596 -25922
rect 28996 -26002 29036 -25942
rect 30556 -26002 30596 -25942
rect 28996 -26022 30596 -26002
rect 22996 -26122 23096 -26102
rect 30696 -26102 30716 -22842
rect 30776 -26102 30796 -22842
rect 30696 -26122 30796 -26102
rect 22996 -26142 30796 -26122
rect 22996 -26202 23116 -26142
rect 30676 -26202 30796 -26142
rect 22996 -26222 30796 -26202
rect 30876 -24582 32576 -24562
rect 30876 -24642 30996 -24582
rect 32456 -24642 32576 -24582
rect 30876 -24662 32576 -24642
rect 30876 -24682 30976 -24662
rect 22816 -26442 22916 -26422
rect 21216 -26462 22916 -26442
rect 21216 -26522 21336 -26462
rect 22796 -26522 22916 -26462
rect 21216 -26542 22916 -26522
rect 23696 -26242 23796 -26222
rect 23696 -28002 23716 -26242
rect 23776 -28002 23796 -26242
rect 29896 -26242 29996 -26222
rect 23696 -28022 23796 -28002
rect 29896 -28002 29916 -26242
rect 29976 -28002 29996 -26242
rect 30876 -26422 30896 -24682
rect 30956 -26422 30976 -24682
rect 32476 -24682 32576 -24662
rect 30876 -26442 30976 -26422
rect 32476 -26422 32496 -24682
rect 32556 -26422 32576 -24682
rect 32476 -26442 32576 -26422
rect 30876 -26462 32576 -26442
rect 30876 -26522 30996 -26462
rect 32456 -26522 32576 -26462
rect 30876 -26542 32576 -26522
rect 29896 -28022 29996 -28002
rect 23696 -28042 29996 -28022
rect 23696 -28102 23816 -28042
rect 29876 -28102 29996 -28042
rect 23696 -28122 29996 -28102
<< nsubdiff >>
rect 23436 -18662 30356 -18642
rect 23436 -19622 23476 -18662
rect 20296 -19642 23476 -19622
rect 20296 -19802 20496 -19642
rect 23416 -19802 23476 -19642
rect 23596 -18822 23636 -18662
rect 30156 -18822 30196 -18662
rect 23596 -18842 30196 -18822
rect 23596 -19802 23636 -18842
rect 20296 -19822 23636 -19802
rect 23736 -19662 30036 -19642
rect 23736 -19722 23856 -19662
rect 29916 -19722 30036 -19662
rect 23736 -19742 30036 -19722
rect 23736 -19762 23836 -19742
rect 20296 -19842 20496 -19822
rect 20296 -28202 20316 -19842
rect 20476 -28202 20496 -19842
rect 20736 -20042 23636 -20022
rect 20736 -20102 20856 -20042
rect 23516 -20102 23636 -20042
rect 20736 -20122 23636 -20102
rect 20736 -20142 20836 -20122
rect 20736 -22402 20756 -20142
rect 20816 -22402 20836 -20142
rect 23536 -20142 23636 -20122
rect 20736 -22422 20836 -22402
rect 23536 -22402 23556 -20142
rect 23616 -22402 23636 -20142
rect 23736 -21922 23756 -19762
rect 23816 -21922 23836 -19762
rect 29936 -19762 30036 -19742
rect 23736 -21942 23836 -21922
rect 29936 -21922 29956 -19762
rect 30016 -21922 30036 -19762
rect 30156 -19802 30196 -18842
rect 30316 -19622 30356 -18662
rect 30316 -19642 33496 -19622
rect 30316 -19802 30356 -19642
rect 33276 -19802 33496 -19642
rect 30156 -19822 33496 -19802
rect 33296 -19842 33496 -19822
rect 29936 -21942 30036 -21922
rect 23736 -21962 30036 -21942
rect 23736 -22022 23856 -21962
rect 29916 -22022 30036 -21962
rect 23736 -22042 30036 -22022
rect 30136 -20042 33036 -20022
rect 30136 -20102 30256 -20042
rect 32916 -20102 33036 -20042
rect 30136 -20122 33036 -20102
rect 30136 -20142 30236 -20122
rect 23536 -22422 23636 -22402
rect 20736 -22442 23636 -22422
rect 20736 -22502 20856 -22442
rect 23516 -22502 23636 -22442
rect 20736 -22522 23636 -22502
rect 30136 -22402 30156 -20142
rect 30216 -22402 30236 -20142
rect 32936 -20142 33036 -20122
rect 30136 -22422 30236 -22402
rect 32936 -22402 32956 -20142
rect 33016 -22402 33036 -20142
rect 32936 -22422 33036 -22402
rect 30136 -22442 33036 -22422
rect 30136 -22502 30256 -22442
rect 32916 -22502 33036 -22442
rect 30136 -22522 33036 -22502
rect 21596 -22742 22596 -22722
rect 21596 -22802 21716 -22742
rect 22476 -22802 22596 -22742
rect 21596 -22822 22596 -22802
rect 21596 -22842 21696 -22822
rect 21596 -24102 21616 -22842
rect 21676 -24102 21696 -22842
rect 22496 -22842 22596 -22822
rect 21596 -24122 21696 -24102
rect 22496 -24102 22516 -22842
rect 22576 -24102 22596 -22842
rect 22496 -24122 22596 -24102
rect 21596 -24142 22596 -24122
rect 21596 -24202 21716 -24142
rect 22476 -24202 22596 -24142
rect 21596 -24222 22596 -24202
rect 31196 -22742 32196 -22722
rect 31196 -22802 31316 -22742
rect 32076 -22802 32196 -22742
rect 31196 -22822 32196 -22802
rect 31196 -22842 31296 -22822
rect 31196 -24102 31216 -22842
rect 31276 -24102 31296 -22842
rect 32096 -22842 32196 -22822
rect 31196 -24122 31296 -24102
rect 32096 -24102 32116 -22842
rect 32176 -24102 32196 -22842
rect 32096 -24122 32196 -24102
rect 31196 -24142 32196 -24122
rect 31196 -24202 31316 -24142
rect 32076 -24202 32196 -24142
rect 31196 -24222 32196 -24202
rect 20296 -28222 20496 -28202
rect 33296 -28202 33316 -19842
rect 33476 -28202 33496 -19842
rect 33296 -28222 33496 -28202
rect 20296 -28242 23596 -28222
rect 20296 -28402 20516 -28242
rect 23376 -28402 23436 -28242
rect 20296 -28422 23436 -28402
rect 23396 -29402 23436 -28422
rect 23556 -29222 23596 -28242
rect 30156 -28242 33496 -28222
rect 30156 -29222 30196 -28242
rect 23556 -29242 30196 -29222
rect 23556 -29402 23596 -29242
rect 30156 -29402 30196 -29242
rect 30316 -28402 30356 -28242
rect 33276 -28402 33496 -28242
rect 30316 -28422 33496 -28402
rect 30316 -29402 30356 -28422
rect 23396 -29422 30356 -29402
<< psubdiffcont >>
rect 23116 -22802 30676 -22742
rect 21336 -24622 22796 -24562
rect 21236 -26422 21296 -24662
rect 22836 -26422 22896 -24662
rect 23016 -26102 23076 -22842
rect 23236 -23002 24756 -22942
rect 25036 -23002 26556 -22942
rect 27236 -23002 28756 -22942
rect 29036 -23002 30556 -22942
rect 23236 -26002 24756 -25942
rect 25036 -26002 26556 -25942
rect 27236 -26002 28756 -25942
rect 29036 -26002 30556 -25942
rect 30716 -26102 30776 -22842
rect 23116 -26202 30676 -26142
rect 30996 -24642 32456 -24582
rect 21336 -26522 22796 -26462
rect 23716 -28002 23776 -26242
rect 29916 -28002 29976 -26242
rect 30896 -26422 30956 -24682
rect 32496 -26422 32556 -24682
rect 30996 -26522 32456 -26462
rect 23816 -28102 29876 -28042
<< nsubdiffcont >>
rect 20496 -19802 23416 -19642
rect 23476 -19802 23596 -18662
rect 23636 -18822 30156 -18662
rect 23856 -19722 29916 -19662
rect 20316 -28202 20476 -19842
rect 20856 -20102 23516 -20042
rect 20756 -22402 20816 -20142
rect 23556 -22402 23616 -20142
rect 23756 -21922 23816 -19762
rect 29956 -21922 30016 -19762
rect 30196 -19802 30316 -18662
rect 30356 -19802 33276 -19642
rect 23856 -22022 29916 -21962
rect 30256 -20102 32916 -20042
rect 20856 -22502 23516 -22442
rect 30156 -22402 30216 -20142
rect 32956 -22402 33016 -20142
rect 30256 -22502 32916 -22442
rect 21716 -22802 22476 -22742
rect 21616 -24102 21676 -22842
rect 22516 -24102 22576 -22842
rect 21716 -24202 22476 -24142
rect 31316 -22802 32076 -22742
rect 31216 -24102 31276 -22842
rect 32116 -24102 32176 -22842
rect 31316 -24202 32076 -24142
rect 33316 -28202 33476 -19842
rect 20516 -28402 23376 -28242
rect 23436 -29402 23556 -28242
rect 23596 -29402 30156 -29242
rect 30196 -29402 30316 -28242
rect 30356 -28402 33276 -28242
<< poly >>
rect 20856 -22342 20886 -20172
rect 20960 -20222 21210 -20196
rect 21268 -20222 21518 -20196
rect 21576 -20222 21826 -20196
rect 21884 -20222 22134 -20196
rect 22192 -20222 22442 -20196
rect 22500 -20222 22750 -20196
rect 22808 -20222 23058 -20196
rect 23116 -20222 23366 -20196
rect 20960 -22269 21210 -22222
rect 20960 -22303 20976 -22269
rect 21194 -22303 21210 -22269
rect 20960 -22319 21210 -22303
rect 21268 -22269 21518 -22222
rect 21268 -22303 21284 -22269
rect 21502 -22303 21518 -22269
rect 21268 -22319 21518 -22303
rect 21576 -22269 21826 -22222
rect 21576 -22303 21592 -22269
rect 21810 -22303 21826 -22269
rect 21576 -22319 21826 -22303
rect 21884 -22269 22134 -22222
rect 21884 -22303 21900 -22269
rect 22118 -22303 22134 -22269
rect 21884 -22319 22134 -22303
rect 22192 -22269 22442 -22222
rect 22192 -22303 22208 -22269
rect 22426 -22303 22442 -22269
rect 22192 -22319 22442 -22303
rect 22500 -22269 22750 -22222
rect 22500 -22303 22516 -22269
rect 22734 -22303 22750 -22269
rect 22500 -22319 22750 -22303
rect 22808 -22269 23058 -22222
rect 22808 -22303 22824 -22269
rect 23042 -22303 23058 -22269
rect 22808 -22319 23058 -22303
rect 23116 -22269 23366 -22222
rect 23116 -22303 23132 -22269
rect 23350 -22303 23366 -22269
rect 23116 -22319 23366 -22303
rect 23446 -22342 23476 -20172
rect 23960 -19862 24060 -19836
rect 24118 -19862 24218 -19836
rect 24395 -19867 24645 -19841
rect 24703 -19867 24953 -19841
rect 25011 -19867 25261 -19841
rect 25319 -19867 25569 -19841
rect 25627 -19867 25877 -19841
rect 25935 -19867 26185 -19841
rect 26243 -19867 26493 -19841
rect 26551 -19867 26801 -19841
rect 26859 -19867 27109 -19841
rect 27167 -19867 27417 -19841
rect 27475 -19867 27725 -19841
rect 27783 -19867 28033 -19841
rect 28091 -19867 28341 -19841
rect 28399 -19867 28649 -19841
rect 28707 -19867 28957 -19841
rect 29015 -19867 29265 -19841
rect 29500 -19862 29600 -19836
rect 29658 -19862 29758 -19836
rect 23960 -21789 24060 -21742
rect 23960 -21823 23976 -21789
rect 24044 -21823 24060 -21789
rect 23960 -21839 24060 -21823
rect 24118 -21789 24218 -21742
rect 24118 -21823 24134 -21789
rect 24202 -21823 24218 -21789
rect 24118 -21839 24218 -21823
rect 24395 -21794 24645 -21747
rect 24395 -21828 24411 -21794
rect 24629 -21828 24645 -21794
rect 24395 -21844 24645 -21828
rect 24703 -21794 24953 -21747
rect 24703 -21828 24719 -21794
rect 24937 -21828 24953 -21794
rect 24703 -21844 24953 -21828
rect 25011 -21794 25261 -21747
rect 25011 -21828 25027 -21794
rect 25245 -21828 25261 -21794
rect 25011 -21844 25261 -21828
rect 25319 -21794 25569 -21747
rect 25319 -21828 25335 -21794
rect 25553 -21828 25569 -21794
rect 25319 -21844 25569 -21828
rect 25627 -21794 25877 -21747
rect 25627 -21828 25643 -21794
rect 25861 -21828 25877 -21794
rect 25627 -21844 25877 -21828
rect 25935 -21794 26185 -21747
rect 25935 -21828 25951 -21794
rect 26169 -21828 26185 -21794
rect 25935 -21844 26185 -21828
rect 26243 -21794 26493 -21747
rect 26243 -21828 26259 -21794
rect 26477 -21828 26493 -21794
rect 26243 -21844 26493 -21828
rect 26551 -21794 26801 -21747
rect 26551 -21828 26567 -21794
rect 26785 -21828 26801 -21794
rect 26551 -21844 26801 -21828
rect 26859 -21794 27109 -21747
rect 26859 -21828 26875 -21794
rect 27093 -21828 27109 -21794
rect 26859 -21844 27109 -21828
rect 27167 -21794 27417 -21747
rect 27167 -21828 27183 -21794
rect 27401 -21828 27417 -21794
rect 27167 -21844 27417 -21828
rect 27475 -21794 27725 -21747
rect 27475 -21828 27491 -21794
rect 27709 -21828 27725 -21794
rect 27475 -21844 27725 -21828
rect 27783 -21794 28033 -21747
rect 27783 -21828 27799 -21794
rect 28017 -21828 28033 -21794
rect 27783 -21844 28033 -21828
rect 28091 -21794 28341 -21747
rect 28091 -21828 28107 -21794
rect 28325 -21828 28341 -21794
rect 28091 -21844 28341 -21828
rect 28399 -21794 28649 -21747
rect 28399 -21828 28415 -21794
rect 28633 -21828 28649 -21794
rect 28399 -21844 28649 -21828
rect 28707 -21794 28957 -21747
rect 28707 -21828 28723 -21794
rect 28941 -21828 28957 -21794
rect 28707 -21844 28957 -21828
rect 29015 -21794 29265 -21747
rect 29015 -21828 29031 -21794
rect 29249 -21828 29265 -21794
rect 29015 -21844 29265 -21828
rect 29500 -21789 29600 -21742
rect 29500 -21823 29516 -21789
rect 29584 -21823 29600 -21789
rect 29500 -21839 29600 -21823
rect 29658 -21789 29758 -21742
rect 29658 -21823 29674 -21789
rect 29742 -21823 29758 -21789
rect 29658 -21839 29758 -21823
rect 30296 -22342 30326 -20182
rect 30400 -20222 30650 -20196
rect 30708 -20222 30958 -20196
rect 31016 -20222 31266 -20196
rect 31324 -20222 31574 -20196
rect 31632 -20222 31882 -20196
rect 31940 -20222 32190 -20196
rect 32248 -20222 32498 -20196
rect 32556 -20222 32806 -20196
rect 30400 -22269 30650 -22222
rect 30400 -22303 30416 -22269
rect 30634 -22303 30650 -22269
rect 30400 -22319 30650 -22303
rect 30708 -22269 30958 -22222
rect 30708 -22303 30724 -22269
rect 30942 -22303 30958 -22269
rect 30708 -22319 30958 -22303
rect 31016 -22269 31266 -22222
rect 31016 -22303 31032 -22269
rect 31250 -22303 31266 -22269
rect 31016 -22319 31266 -22303
rect 31324 -22269 31574 -22222
rect 31324 -22303 31340 -22269
rect 31558 -22303 31574 -22269
rect 31324 -22319 31574 -22303
rect 31632 -22269 31882 -22222
rect 31632 -22303 31648 -22269
rect 31866 -22303 31882 -22269
rect 31632 -22319 31882 -22303
rect 31940 -22269 32190 -22222
rect 31940 -22303 31956 -22269
rect 32174 -22303 32190 -22269
rect 31940 -22319 32190 -22303
rect 32248 -22269 32498 -22222
rect 32248 -22303 32264 -22269
rect 32482 -22303 32498 -22269
rect 32248 -22319 32498 -22303
rect 32556 -22269 32806 -22222
rect 32556 -22303 32572 -22269
rect 32790 -22303 32806 -22269
rect 32556 -22319 32806 -22303
rect 32886 -22342 32916 -20182
rect 21816 -24042 21846 -22892
rect 21920 -22922 22100 -22896
rect 22158 -22922 22338 -22896
rect 21920 -23969 22100 -23922
rect 21920 -24003 21936 -23969
rect 22084 -24003 22100 -23969
rect 21920 -24019 22100 -24003
rect 22158 -23969 22338 -23922
rect 22158 -24003 22174 -23969
rect 22322 -24003 22338 -23969
rect 22158 -24019 22338 -24003
rect 22416 -24042 22446 -22892
rect 21336 -26342 21396 -24722
rect 21474 -24754 21724 -24728
rect 21782 -24754 22032 -24728
rect 22090 -24754 22340 -24728
rect 22398 -24754 22648 -24728
rect 21474 -26292 21724 -26254
rect 21474 -26326 21490 -26292
rect 21708 -26326 21724 -26292
rect 21474 -26342 21724 -26326
rect 21782 -26292 22032 -26254
rect 21782 -26326 21798 -26292
rect 22016 -26326 22032 -26292
rect 21782 -26342 22032 -26326
rect 22090 -26292 22340 -26254
rect 22090 -26326 22106 -26292
rect 22324 -26326 22340 -26292
rect 22090 -26342 22340 -26326
rect 22398 -26292 22648 -26254
rect 22398 -26326 22414 -26292
rect 22632 -26326 22648 -26292
rect 22398 -26342 22648 -26326
rect 22726 -26342 22786 -24722
rect 23414 -23144 23514 -23118
rect 23572 -23144 23672 -23118
rect 23854 -23144 23954 -23118
rect 24012 -23144 24112 -23118
rect 24294 -23144 24394 -23118
rect 24452 -23144 24552 -23118
rect 23414 -24132 23514 -24094
rect 23414 -24166 23430 -24132
rect 23498 -24166 23514 -24132
rect 23414 -24182 23514 -24166
rect 23572 -24132 23672 -24094
rect 23572 -24166 23588 -24132
rect 23656 -24166 23672 -24132
rect 23572 -24182 23672 -24166
rect 23854 -24132 23954 -24094
rect 23854 -24166 23870 -24132
rect 23938 -24166 23954 -24132
rect 23854 -24182 23954 -24166
rect 24012 -24132 24112 -24094
rect 24012 -24166 24028 -24132
rect 24096 -24166 24112 -24132
rect 24012 -24182 24112 -24166
rect 24294 -24132 24394 -24094
rect 24294 -24166 24310 -24132
rect 24378 -24166 24394 -24132
rect 24294 -24182 24394 -24166
rect 24452 -24132 24552 -24094
rect 24452 -24166 24468 -24132
rect 24536 -24166 24552 -24132
rect 24452 -24182 24552 -24166
rect 25214 -23144 25314 -23118
rect 25372 -23144 25472 -23118
rect 25654 -23144 25754 -23118
rect 25812 -23144 25912 -23118
rect 26094 -23144 26194 -23118
rect 26252 -23144 26352 -23118
rect 25214 -24132 25314 -24094
rect 25214 -24166 25230 -24132
rect 25298 -24166 25314 -24132
rect 25214 -24182 25314 -24166
rect 25372 -24132 25472 -24094
rect 25372 -24166 25388 -24132
rect 25456 -24166 25472 -24132
rect 25372 -24182 25472 -24166
rect 25654 -24132 25754 -24094
rect 25654 -24166 25670 -24132
rect 25738 -24166 25754 -24132
rect 25654 -24182 25754 -24166
rect 25812 -24132 25912 -24094
rect 25812 -24166 25828 -24132
rect 25896 -24166 25912 -24132
rect 25812 -24182 25912 -24166
rect 26094 -24132 26194 -24094
rect 26094 -24166 26110 -24132
rect 26178 -24166 26194 -24132
rect 26094 -24182 26194 -24166
rect 26252 -24132 26352 -24094
rect 26252 -24166 26268 -24132
rect 26336 -24166 26352 -24132
rect 26252 -24182 26352 -24166
rect 27414 -23144 27514 -23118
rect 27572 -23144 27672 -23118
rect 27854 -23144 27954 -23118
rect 28012 -23144 28112 -23118
rect 28294 -23144 28394 -23118
rect 28452 -23144 28552 -23118
rect 27414 -24132 27514 -24094
rect 27414 -24166 27430 -24132
rect 27498 -24166 27514 -24132
rect 27414 -24182 27514 -24166
rect 27572 -24132 27672 -24094
rect 27572 -24166 27588 -24132
rect 27656 -24166 27672 -24132
rect 27572 -24182 27672 -24166
rect 27854 -24132 27954 -24094
rect 27854 -24166 27870 -24132
rect 27938 -24166 27954 -24132
rect 27854 -24182 27954 -24166
rect 28012 -24132 28112 -24094
rect 28012 -24166 28028 -24132
rect 28096 -24166 28112 -24132
rect 28012 -24182 28112 -24166
rect 28294 -24132 28394 -24094
rect 28294 -24166 28310 -24132
rect 28378 -24166 28394 -24132
rect 28294 -24182 28394 -24166
rect 28452 -24132 28552 -24094
rect 28452 -24166 28468 -24132
rect 28536 -24166 28552 -24132
rect 28452 -24182 28552 -24166
rect 29214 -23144 29314 -23118
rect 29372 -23144 29472 -23118
rect 29654 -23144 29754 -23118
rect 29812 -23144 29912 -23118
rect 30094 -23144 30194 -23118
rect 30252 -23144 30352 -23118
rect 29214 -24132 29314 -24094
rect 29214 -24166 29230 -24132
rect 29298 -24166 29314 -24132
rect 29214 -24182 29314 -24166
rect 29372 -24132 29472 -24094
rect 29372 -24166 29388 -24132
rect 29456 -24166 29472 -24132
rect 29372 -24182 29472 -24166
rect 29654 -24132 29754 -24094
rect 29654 -24166 29670 -24132
rect 29738 -24166 29754 -24132
rect 29654 -24182 29754 -24166
rect 29812 -24132 29912 -24094
rect 29812 -24166 29828 -24132
rect 29896 -24166 29912 -24132
rect 29812 -24182 29912 -24166
rect 30094 -24132 30194 -24094
rect 30094 -24166 30110 -24132
rect 30178 -24166 30194 -24132
rect 30094 -24182 30194 -24166
rect 30252 -24132 30352 -24094
rect 30252 -24166 30268 -24132
rect 30336 -24166 30352 -24132
rect 30252 -24182 30352 -24166
rect 23414 -24774 23514 -24758
rect 23414 -24808 23430 -24774
rect 23498 -24808 23514 -24774
rect 23414 -24846 23514 -24808
rect 23572 -24774 23672 -24758
rect 23572 -24808 23588 -24774
rect 23656 -24808 23672 -24774
rect 23572 -24846 23672 -24808
rect 23854 -24774 23954 -24758
rect 23854 -24808 23870 -24774
rect 23938 -24808 23954 -24774
rect 23854 -24846 23954 -24808
rect 24012 -24774 24112 -24758
rect 24012 -24808 24028 -24774
rect 24096 -24808 24112 -24774
rect 24012 -24846 24112 -24808
rect 24294 -24774 24394 -24758
rect 24294 -24808 24310 -24774
rect 24378 -24808 24394 -24774
rect 24294 -24846 24394 -24808
rect 24452 -24774 24552 -24758
rect 24452 -24808 24468 -24774
rect 24536 -24808 24552 -24774
rect 24452 -24846 24552 -24808
rect 23414 -25822 23514 -25796
rect 23572 -25822 23672 -25796
rect 23854 -25822 23954 -25796
rect 24012 -25822 24112 -25796
rect 24294 -25822 24394 -25796
rect 24452 -25822 24552 -25796
rect 25214 -24774 25314 -24758
rect 25214 -24808 25230 -24774
rect 25298 -24808 25314 -24774
rect 25214 -24846 25314 -24808
rect 25372 -24774 25472 -24758
rect 25372 -24808 25388 -24774
rect 25456 -24808 25472 -24774
rect 25372 -24846 25472 -24808
rect 25654 -24774 25754 -24758
rect 25654 -24808 25670 -24774
rect 25738 -24808 25754 -24774
rect 25654 -24846 25754 -24808
rect 25812 -24774 25912 -24758
rect 25812 -24808 25828 -24774
rect 25896 -24808 25912 -24774
rect 25812 -24846 25912 -24808
rect 26094 -24774 26194 -24758
rect 26094 -24808 26110 -24774
rect 26178 -24808 26194 -24774
rect 26094 -24846 26194 -24808
rect 26252 -24774 26352 -24758
rect 26252 -24808 26268 -24774
rect 26336 -24808 26352 -24774
rect 26252 -24846 26352 -24808
rect 25214 -25822 25314 -25796
rect 25372 -25822 25472 -25796
rect 25654 -25822 25754 -25796
rect 25812 -25822 25912 -25796
rect 26094 -25822 26194 -25796
rect 26252 -25822 26352 -25796
rect 27414 -24774 27514 -24758
rect 27414 -24808 27430 -24774
rect 27498 -24808 27514 -24774
rect 27414 -24846 27514 -24808
rect 27572 -24774 27672 -24758
rect 27572 -24808 27588 -24774
rect 27656 -24808 27672 -24774
rect 27572 -24846 27672 -24808
rect 27854 -24774 27954 -24758
rect 27854 -24808 27870 -24774
rect 27938 -24808 27954 -24774
rect 27854 -24846 27954 -24808
rect 28012 -24774 28112 -24758
rect 28012 -24808 28028 -24774
rect 28096 -24808 28112 -24774
rect 28012 -24846 28112 -24808
rect 28294 -24774 28394 -24758
rect 28294 -24808 28310 -24774
rect 28378 -24808 28394 -24774
rect 28294 -24846 28394 -24808
rect 28452 -24774 28552 -24758
rect 28452 -24808 28468 -24774
rect 28536 -24808 28552 -24774
rect 28452 -24846 28552 -24808
rect 27414 -25822 27514 -25796
rect 27572 -25822 27672 -25796
rect 27854 -25822 27954 -25796
rect 28012 -25822 28112 -25796
rect 28294 -25822 28394 -25796
rect 28452 -25822 28552 -25796
rect 29214 -24774 29314 -24758
rect 29214 -24808 29230 -24774
rect 29298 -24808 29314 -24774
rect 29214 -24846 29314 -24808
rect 29372 -24774 29472 -24758
rect 29372 -24808 29388 -24774
rect 29456 -24808 29472 -24774
rect 29372 -24846 29472 -24808
rect 29654 -24774 29754 -24758
rect 29654 -24808 29670 -24774
rect 29738 -24808 29754 -24774
rect 29654 -24846 29754 -24808
rect 29812 -24774 29912 -24758
rect 29812 -24808 29828 -24774
rect 29896 -24808 29912 -24774
rect 29812 -24846 29912 -24808
rect 30094 -24774 30194 -24758
rect 30094 -24808 30110 -24774
rect 30178 -24808 30194 -24774
rect 30094 -24846 30194 -24808
rect 30252 -24774 30352 -24758
rect 30252 -24808 30268 -24774
rect 30336 -24808 30352 -24774
rect 30252 -24846 30352 -24808
rect 29214 -25822 29314 -25796
rect 29372 -25822 29472 -25796
rect 29654 -25822 29754 -25796
rect 29812 -25822 29912 -25796
rect 30094 -25822 30194 -25796
rect 30252 -25822 30352 -25796
rect 31396 -24012 31426 -22862
rect 31500 -22902 31680 -22876
rect 31738 -22902 31918 -22876
rect 31500 -23949 31680 -23902
rect 31500 -23983 31516 -23949
rect 31664 -23983 31680 -23949
rect 31500 -23999 31680 -23983
rect 31738 -23949 31918 -23902
rect 31738 -23983 31754 -23949
rect 31902 -23983 31918 -23949
rect 31738 -23999 31918 -23983
rect 31996 -24012 32026 -22862
rect 23994 -26324 24094 -26308
rect 23994 -26358 24010 -26324
rect 24078 -26358 24094 -26324
rect 23994 -26396 24094 -26358
rect 24152 -26324 24252 -26308
rect 24152 -26358 24168 -26324
rect 24236 -26358 24252 -26324
rect 24152 -26396 24252 -26358
rect 24434 -26324 24684 -26308
rect 24434 -26358 24450 -26324
rect 24668 -26358 24684 -26324
rect 24434 -26396 24684 -26358
rect 24742 -26324 24992 -26308
rect 24742 -26358 24758 -26324
rect 24976 -26358 24992 -26324
rect 24742 -26396 24992 -26358
rect 25050 -26324 25300 -26308
rect 25050 -26358 25066 -26324
rect 25284 -26358 25300 -26324
rect 25050 -26396 25300 -26358
rect 25358 -26324 25608 -26308
rect 25358 -26358 25374 -26324
rect 25592 -26358 25608 -26324
rect 25358 -26396 25608 -26358
rect 25666 -26324 25916 -26308
rect 25666 -26358 25682 -26324
rect 25900 -26358 25916 -26324
rect 25666 -26396 25916 -26358
rect 25974 -26324 26224 -26308
rect 25974 -26358 25990 -26324
rect 26208 -26358 26224 -26324
rect 25974 -26396 26224 -26358
rect 26282 -26324 26532 -26308
rect 26282 -26358 26298 -26324
rect 26516 -26358 26532 -26324
rect 26282 -26396 26532 -26358
rect 26590 -26324 26840 -26308
rect 26590 -26358 26606 -26324
rect 26824 -26358 26840 -26324
rect 26590 -26396 26840 -26358
rect 26898 -26324 27148 -26308
rect 26898 -26358 26914 -26324
rect 27132 -26358 27148 -26324
rect 26898 -26396 27148 -26358
rect 27206 -26324 27456 -26308
rect 27206 -26358 27222 -26324
rect 27440 -26358 27456 -26324
rect 27206 -26396 27456 -26358
rect 27514 -26324 27764 -26308
rect 27514 -26358 27530 -26324
rect 27748 -26358 27764 -26324
rect 27514 -26396 27764 -26358
rect 27822 -26324 28072 -26308
rect 27822 -26358 27838 -26324
rect 28056 -26358 28072 -26324
rect 27822 -26396 28072 -26358
rect 28130 -26324 28380 -26308
rect 28130 -26358 28146 -26324
rect 28364 -26358 28380 -26324
rect 28130 -26396 28380 -26358
rect 28438 -26324 28688 -26308
rect 28438 -26358 28454 -26324
rect 28672 -26358 28688 -26324
rect 28438 -26396 28688 -26358
rect 28746 -26324 28996 -26308
rect 28746 -26358 28762 -26324
rect 28980 -26358 28996 -26324
rect 28746 -26396 28996 -26358
rect 29054 -26324 29304 -26308
rect 29054 -26358 29070 -26324
rect 29288 -26358 29304 -26324
rect 29054 -26396 29304 -26358
rect 29494 -26324 29594 -26308
rect 29494 -26358 29510 -26324
rect 29578 -26358 29594 -26324
rect 29494 -26396 29594 -26358
rect 29652 -26324 29752 -26308
rect 29652 -26358 29668 -26324
rect 29736 -26358 29752 -26324
rect 29652 -26396 29752 -26358
rect 23994 -27922 24094 -27896
rect 24152 -27922 24252 -27896
rect 24434 -27922 24684 -27896
rect 24742 -27922 24992 -27896
rect 25050 -27922 25300 -27896
rect 25358 -27922 25608 -27896
rect 25666 -27922 25916 -27896
rect 25974 -27922 26224 -27896
rect 26282 -27922 26532 -27896
rect 26590 -27922 26840 -27896
rect 26898 -27922 27148 -27896
rect 27206 -27922 27456 -27896
rect 27514 -27922 27764 -27896
rect 27822 -27922 28072 -27896
rect 28130 -27922 28380 -27896
rect 28438 -27922 28688 -27896
rect 28746 -27922 28996 -27896
rect 29054 -27922 29304 -27896
rect 29494 -27922 29594 -27896
rect 29652 -27922 29752 -27896
rect 30996 -26362 31056 -24742
rect 31134 -24774 31384 -24748
rect 31442 -24774 31692 -24748
rect 31750 -24774 32000 -24748
rect 32058 -24774 32308 -24748
rect 31134 -26312 31384 -26274
rect 31134 -26346 31150 -26312
rect 31368 -26346 31384 -26312
rect 31134 -26362 31384 -26346
rect 31442 -26312 31692 -26274
rect 31442 -26346 31458 -26312
rect 31676 -26346 31692 -26312
rect 31442 -26362 31692 -26346
rect 31750 -26312 32000 -26274
rect 31750 -26346 31766 -26312
rect 31984 -26346 32000 -26312
rect 31750 -26362 32000 -26346
rect 32058 -26312 32308 -26274
rect 32058 -26346 32074 -26312
rect 32292 -26346 32308 -26312
rect 32058 -26362 32308 -26346
rect 32386 -26362 32446 -24742
<< polycont >>
rect 20976 -22303 21194 -22269
rect 21284 -22303 21502 -22269
rect 21592 -22303 21810 -22269
rect 21900 -22303 22118 -22269
rect 22208 -22303 22426 -22269
rect 22516 -22303 22734 -22269
rect 22824 -22303 23042 -22269
rect 23132 -22303 23350 -22269
rect 23976 -21823 24044 -21789
rect 24134 -21823 24202 -21789
rect 24411 -21828 24629 -21794
rect 24719 -21828 24937 -21794
rect 25027 -21828 25245 -21794
rect 25335 -21828 25553 -21794
rect 25643 -21828 25861 -21794
rect 25951 -21828 26169 -21794
rect 26259 -21828 26477 -21794
rect 26567 -21828 26785 -21794
rect 26875 -21828 27093 -21794
rect 27183 -21828 27401 -21794
rect 27491 -21828 27709 -21794
rect 27799 -21828 28017 -21794
rect 28107 -21828 28325 -21794
rect 28415 -21828 28633 -21794
rect 28723 -21828 28941 -21794
rect 29031 -21828 29249 -21794
rect 29516 -21823 29584 -21789
rect 29674 -21823 29742 -21789
rect 30416 -22303 30634 -22269
rect 30724 -22303 30942 -22269
rect 31032 -22303 31250 -22269
rect 31340 -22303 31558 -22269
rect 31648 -22303 31866 -22269
rect 31956 -22303 32174 -22269
rect 32264 -22303 32482 -22269
rect 32572 -22303 32790 -22269
rect 21936 -24003 22084 -23969
rect 22174 -24003 22322 -23969
rect 21490 -26326 21708 -26292
rect 21798 -26326 22016 -26292
rect 22106 -26326 22324 -26292
rect 22414 -26326 22632 -26292
rect 23430 -24166 23498 -24132
rect 23588 -24166 23656 -24132
rect 23870 -24166 23938 -24132
rect 24028 -24166 24096 -24132
rect 24310 -24166 24378 -24132
rect 24468 -24166 24536 -24132
rect 25230 -24166 25298 -24132
rect 25388 -24166 25456 -24132
rect 25670 -24166 25738 -24132
rect 25828 -24166 25896 -24132
rect 26110 -24166 26178 -24132
rect 26268 -24166 26336 -24132
rect 27430 -24166 27498 -24132
rect 27588 -24166 27656 -24132
rect 27870 -24166 27938 -24132
rect 28028 -24166 28096 -24132
rect 28310 -24166 28378 -24132
rect 28468 -24166 28536 -24132
rect 29230 -24166 29298 -24132
rect 29388 -24166 29456 -24132
rect 29670 -24166 29738 -24132
rect 29828 -24166 29896 -24132
rect 30110 -24166 30178 -24132
rect 30268 -24166 30336 -24132
rect 23430 -24808 23498 -24774
rect 23588 -24808 23656 -24774
rect 23870 -24808 23938 -24774
rect 24028 -24808 24096 -24774
rect 24310 -24808 24378 -24774
rect 24468 -24808 24536 -24774
rect 25230 -24808 25298 -24774
rect 25388 -24808 25456 -24774
rect 25670 -24808 25738 -24774
rect 25828 -24808 25896 -24774
rect 26110 -24808 26178 -24774
rect 26268 -24808 26336 -24774
rect 27430 -24808 27498 -24774
rect 27588 -24808 27656 -24774
rect 27870 -24808 27938 -24774
rect 28028 -24808 28096 -24774
rect 28310 -24808 28378 -24774
rect 28468 -24808 28536 -24774
rect 29230 -24808 29298 -24774
rect 29388 -24808 29456 -24774
rect 29670 -24808 29738 -24774
rect 29828 -24808 29896 -24774
rect 30110 -24808 30178 -24774
rect 30268 -24808 30336 -24774
rect 31516 -23983 31664 -23949
rect 31754 -23983 31902 -23949
rect 24010 -26358 24078 -26324
rect 24168 -26358 24236 -26324
rect 24450 -26358 24668 -26324
rect 24758 -26358 24976 -26324
rect 25066 -26358 25284 -26324
rect 25374 -26358 25592 -26324
rect 25682 -26358 25900 -26324
rect 25990 -26358 26208 -26324
rect 26298 -26358 26516 -26324
rect 26606 -26358 26824 -26324
rect 26914 -26358 27132 -26324
rect 27222 -26358 27440 -26324
rect 27530 -26358 27748 -26324
rect 27838 -26358 28056 -26324
rect 28146 -26358 28364 -26324
rect 28454 -26358 28672 -26324
rect 28762 -26358 28980 -26324
rect 29070 -26358 29288 -26324
rect 29510 -26358 29578 -26324
rect 29668 -26358 29736 -26324
rect 31150 -26346 31368 -26312
rect 31458 -26346 31676 -26312
rect 31766 -26346 31984 -26312
rect 32074 -26346 32292 -26312
<< locali >>
rect 23436 -18662 30356 -18642
rect 23436 -19622 23476 -18662
rect 20296 -19642 23476 -19622
rect 20296 -19802 20496 -19642
rect 23416 -19802 23476 -19642
rect 23596 -18822 23636 -18662
rect 30156 -18822 30196 -18662
rect 23596 -18922 30196 -18822
rect 23596 -19002 23656 -18922
rect 23736 -19002 23776 -18922
rect 23856 -19002 23896 -18922
rect 23976 -19002 24016 -18922
rect 24096 -19002 24136 -18922
rect 24216 -19002 24256 -18922
rect 24336 -19002 24376 -18922
rect 24456 -19002 24496 -18922
rect 24576 -19002 24616 -18922
rect 24696 -19002 24736 -18922
rect 24816 -19002 24856 -18922
rect 24936 -19002 24976 -18922
rect 25056 -19002 25096 -18922
rect 25176 -19002 25216 -18922
rect 25296 -19002 25336 -18922
rect 25416 -19002 25456 -18922
rect 25536 -19002 25576 -18922
rect 25656 -19002 25696 -18922
rect 25776 -19002 25816 -18922
rect 25896 -19002 25936 -18922
rect 26016 -19002 26056 -18922
rect 26136 -19002 26176 -18922
rect 26256 -19002 26296 -18922
rect 26376 -19002 26416 -18922
rect 26496 -19002 26536 -18922
rect 26616 -19002 26656 -18922
rect 26736 -19002 26776 -18922
rect 26856 -19002 26896 -18922
rect 26976 -19002 27016 -18922
rect 27096 -19002 27136 -18922
rect 27216 -19002 27256 -18922
rect 27336 -19002 27376 -18922
rect 27456 -19002 27496 -18922
rect 27576 -19002 27616 -18922
rect 27696 -19002 27736 -18922
rect 27816 -19002 27856 -18922
rect 27936 -19002 27976 -18922
rect 28056 -19002 28096 -18922
rect 28176 -19002 28216 -18922
rect 28296 -19002 28336 -18922
rect 28416 -19002 28456 -18922
rect 28536 -19002 28576 -18922
rect 28656 -19002 28696 -18922
rect 28776 -19002 28816 -18922
rect 28896 -19002 28936 -18922
rect 29016 -19002 29056 -18922
rect 29136 -19002 29176 -18922
rect 29256 -19002 29296 -18922
rect 29376 -19002 29416 -18922
rect 29496 -19002 29536 -18922
rect 29616 -19002 29656 -18922
rect 29736 -19002 29776 -18922
rect 29856 -19002 29896 -18922
rect 29976 -19002 30016 -18922
rect 30096 -19002 30196 -18922
rect 23596 -19042 30196 -19002
rect 23596 -19122 23656 -19042
rect 23736 -19122 23776 -19042
rect 23856 -19122 23896 -19042
rect 23976 -19122 24016 -19042
rect 24096 -19122 24136 -19042
rect 24216 -19122 24256 -19042
rect 24336 -19122 24376 -19042
rect 24456 -19122 24496 -19042
rect 24576 -19122 24616 -19042
rect 24696 -19122 24736 -19042
rect 24816 -19122 24856 -19042
rect 24936 -19122 24976 -19042
rect 25056 -19122 25096 -19042
rect 25176 -19122 25216 -19042
rect 25296 -19122 25336 -19042
rect 25416 -19122 25456 -19042
rect 25536 -19122 25576 -19042
rect 25656 -19122 25696 -19042
rect 25776 -19122 25816 -19042
rect 25896 -19122 25936 -19042
rect 26016 -19122 26056 -19042
rect 26136 -19122 26176 -19042
rect 26256 -19122 26296 -19042
rect 26376 -19122 26416 -19042
rect 26496 -19122 26536 -19042
rect 26616 -19122 26656 -19042
rect 26736 -19122 26776 -19042
rect 26856 -19122 26896 -19042
rect 26976 -19122 27016 -19042
rect 27096 -19122 27136 -19042
rect 27216 -19122 27256 -19042
rect 27336 -19122 27376 -19042
rect 27456 -19122 27496 -19042
rect 27576 -19122 27616 -19042
rect 27696 -19122 27736 -19042
rect 27816 -19122 27856 -19042
rect 27936 -19122 27976 -19042
rect 28056 -19122 28096 -19042
rect 28176 -19122 28216 -19042
rect 28296 -19122 28336 -19042
rect 28416 -19122 28456 -19042
rect 28536 -19122 28576 -19042
rect 28656 -19122 28696 -19042
rect 28776 -19122 28816 -19042
rect 28896 -19122 28936 -19042
rect 29016 -19122 29056 -19042
rect 29136 -19122 29176 -19042
rect 29256 -19122 29296 -19042
rect 29376 -19122 29416 -19042
rect 29496 -19122 29536 -19042
rect 29616 -19122 29656 -19042
rect 29736 -19122 29776 -19042
rect 29856 -19122 29896 -19042
rect 29976 -19122 30016 -19042
rect 30096 -19122 30196 -19042
rect 23596 -19162 30196 -19122
rect 23596 -19242 23656 -19162
rect 23736 -19242 23776 -19162
rect 23856 -19242 23896 -19162
rect 23976 -19242 24016 -19162
rect 24096 -19242 24136 -19162
rect 24216 -19242 24256 -19162
rect 24336 -19242 24376 -19162
rect 24456 -19242 24496 -19162
rect 24576 -19242 24616 -19162
rect 24696 -19242 24736 -19162
rect 24816 -19242 24856 -19162
rect 24936 -19242 24976 -19162
rect 25056 -19242 25096 -19162
rect 25176 -19242 25216 -19162
rect 25296 -19242 25336 -19162
rect 25416 -19242 25456 -19162
rect 25536 -19242 25576 -19162
rect 25656 -19242 25696 -19162
rect 25776 -19242 25816 -19162
rect 25896 -19242 25936 -19162
rect 26016 -19242 26056 -19162
rect 26136 -19242 26176 -19162
rect 26256 -19242 26296 -19162
rect 26376 -19242 26416 -19162
rect 26496 -19242 26536 -19162
rect 26616 -19242 26656 -19162
rect 26736 -19242 26776 -19162
rect 26856 -19242 26896 -19162
rect 26976 -19242 27016 -19162
rect 27096 -19242 27136 -19162
rect 27216 -19242 27256 -19162
rect 27336 -19242 27376 -19162
rect 27456 -19242 27496 -19162
rect 27576 -19242 27616 -19162
rect 27696 -19242 27736 -19162
rect 27816 -19242 27856 -19162
rect 27936 -19242 27976 -19162
rect 28056 -19242 28096 -19162
rect 28176 -19242 28216 -19162
rect 28296 -19242 28336 -19162
rect 28416 -19242 28456 -19162
rect 28536 -19242 28576 -19162
rect 28656 -19242 28696 -19162
rect 28776 -19242 28816 -19162
rect 28896 -19242 28936 -19162
rect 29016 -19242 29056 -19162
rect 29136 -19242 29176 -19162
rect 29256 -19242 29296 -19162
rect 29376 -19242 29416 -19162
rect 29496 -19242 29536 -19162
rect 29616 -19242 29656 -19162
rect 29736 -19242 29776 -19162
rect 29856 -19242 29896 -19162
rect 29976 -19242 30016 -19162
rect 30096 -19242 30196 -19162
rect 23596 -19282 30196 -19242
rect 23596 -19362 23656 -19282
rect 23736 -19362 23776 -19282
rect 23856 -19362 23896 -19282
rect 23976 -19362 24016 -19282
rect 24096 -19362 24136 -19282
rect 24216 -19362 24256 -19282
rect 24336 -19362 24376 -19282
rect 24456 -19362 24496 -19282
rect 24576 -19362 24616 -19282
rect 24696 -19362 24736 -19282
rect 24816 -19362 24856 -19282
rect 24936 -19362 24976 -19282
rect 25056 -19362 25096 -19282
rect 25176 -19362 25216 -19282
rect 25296 -19362 25336 -19282
rect 25416 -19362 25456 -19282
rect 25536 -19362 25576 -19282
rect 25656 -19362 25696 -19282
rect 25776 -19362 25816 -19282
rect 25896 -19362 25936 -19282
rect 26016 -19362 26056 -19282
rect 26136 -19362 26176 -19282
rect 26256 -19362 26296 -19282
rect 26376 -19362 26416 -19282
rect 26496 -19362 26536 -19282
rect 26616 -19362 26656 -19282
rect 26736 -19362 26776 -19282
rect 26856 -19362 26896 -19282
rect 26976 -19362 27016 -19282
rect 27096 -19362 27136 -19282
rect 27216 -19362 27256 -19282
rect 27336 -19362 27376 -19282
rect 27456 -19362 27496 -19282
rect 27576 -19362 27616 -19282
rect 27696 -19362 27736 -19282
rect 27816 -19362 27856 -19282
rect 27936 -19362 27976 -19282
rect 28056 -19362 28096 -19282
rect 28176 -19362 28216 -19282
rect 28296 -19362 28336 -19282
rect 28416 -19362 28456 -19282
rect 28536 -19362 28576 -19282
rect 28656 -19362 28696 -19282
rect 28776 -19362 28816 -19282
rect 28896 -19362 28936 -19282
rect 29016 -19362 29056 -19282
rect 29136 -19362 29176 -19282
rect 29256 -19362 29296 -19282
rect 29376 -19362 29416 -19282
rect 29496 -19362 29536 -19282
rect 29616 -19362 29656 -19282
rect 29736 -19362 29776 -19282
rect 29856 -19362 29896 -19282
rect 29976 -19362 30016 -19282
rect 30096 -19362 30196 -19282
rect 23596 -19402 30196 -19362
rect 23596 -19482 23656 -19402
rect 23736 -19482 23776 -19402
rect 23856 -19482 23896 -19402
rect 23976 -19482 24016 -19402
rect 24096 -19482 24136 -19402
rect 24216 -19482 24256 -19402
rect 24336 -19482 24376 -19402
rect 24456 -19482 24496 -19402
rect 24576 -19482 24616 -19402
rect 24696 -19482 24736 -19402
rect 24816 -19482 24856 -19402
rect 24936 -19482 24976 -19402
rect 25056 -19482 25096 -19402
rect 25176 -19482 25216 -19402
rect 25296 -19482 25336 -19402
rect 25416 -19482 25456 -19402
rect 25536 -19482 25576 -19402
rect 25656 -19482 25696 -19402
rect 25776 -19482 25816 -19402
rect 25896 -19482 25936 -19402
rect 26016 -19482 26056 -19402
rect 26136 -19482 26176 -19402
rect 26256 -19482 26296 -19402
rect 26376 -19482 26416 -19402
rect 26496 -19482 26536 -19402
rect 26616 -19482 26656 -19402
rect 26736 -19482 26776 -19402
rect 26856 -19482 26896 -19402
rect 26976 -19482 27016 -19402
rect 27096 -19482 27136 -19402
rect 27216 -19482 27256 -19402
rect 27336 -19482 27376 -19402
rect 27456 -19482 27496 -19402
rect 27576 -19482 27616 -19402
rect 27696 -19482 27736 -19402
rect 27816 -19482 27856 -19402
rect 27936 -19482 27976 -19402
rect 28056 -19482 28096 -19402
rect 28176 -19482 28216 -19402
rect 28296 -19482 28336 -19402
rect 28416 -19482 28456 -19402
rect 28536 -19482 28576 -19402
rect 28656 -19482 28696 -19402
rect 28776 -19482 28816 -19402
rect 28896 -19482 28936 -19402
rect 29016 -19482 29056 -19402
rect 29136 -19482 29176 -19402
rect 29256 -19482 29296 -19402
rect 29376 -19482 29416 -19402
rect 29496 -19482 29536 -19402
rect 29616 -19482 29656 -19402
rect 29736 -19482 29776 -19402
rect 29856 -19482 29896 -19402
rect 29976 -19482 30016 -19402
rect 30096 -19482 30196 -19402
rect 23596 -19522 30196 -19482
rect 23596 -19602 23656 -19522
rect 23736 -19602 23776 -19522
rect 23856 -19602 23896 -19522
rect 23976 -19602 24016 -19522
rect 24096 -19602 24136 -19522
rect 24216 -19602 24256 -19522
rect 24336 -19602 24376 -19522
rect 24456 -19602 24496 -19522
rect 24576 -19602 24616 -19522
rect 24696 -19602 24736 -19522
rect 24816 -19602 24856 -19522
rect 24936 -19602 24976 -19522
rect 25056 -19602 25096 -19522
rect 25176 -19602 25216 -19522
rect 25296 -19602 25336 -19522
rect 25416 -19602 25456 -19522
rect 25536 -19602 25576 -19522
rect 25656 -19602 25696 -19522
rect 25776 -19602 25816 -19522
rect 25896 -19602 25936 -19522
rect 26016 -19602 26056 -19522
rect 26136 -19602 26176 -19522
rect 26256 -19602 26296 -19522
rect 26376 -19602 26416 -19522
rect 26496 -19602 26536 -19522
rect 26616 -19602 26656 -19522
rect 26736 -19602 26776 -19522
rect 26856 -19602 26896 -19522
rect 26976 -19602 27016 -19522
rect 27096 -19602 27136 -19522
rect 27216 -19602 27256 -19522
rect 27336 -19602 27376 -19522
rect 27456 -19602 27496 -19522
rect 27576 -19602 27616 -19522
rect 27696 -19602 27736 -19522
rect 27816 -19602 27856 -19522
rect 27936 -19602 27976 -19522
rect 28056 -19602 28096 -19522
rect 28176 -19602 28216 -19522
rect 28296 -19602 28336 -19522
rect 28416 -19602 28456 -19522
rect 28536 -19602 28576 -19522
rect 28656 -19602 28696 -19522
rect 28776 -19602 28816 -19522
rect 28896 -19602 28936 -19522
rect 29016 -19602 29056 -19522
rect 29136 -19602 29176 -19522
rect 29256 -19602 29296 -19522
rect 29376 -19602 29416 -19522
rect 29496 -19602 29536 -19522
rect 29616 -19602 29656 -19522
rect 29736 -19602 29776 -19522
rect 29856 -19602 29896 -19522
rect 29976 -19602 30016 -19522
rect 30096 -19602 30196 -19522
rect 23596 -19662 30196 -19602
rect 23596 -19722 23856 -19662
rect 29916 -19722 30196 -19662
rect 23596 -19742 30196 -19722
rect 23596 -19762 23836 -19742
rect 23596 -19802 23756 -19762
rect 20296 -19842 23756 -19802
rect 20296 -28202 20316 -19842
rect 20476 -20042 23756 -19842
rect 20476 -20102 20856 -20042
rect 23516 -20102 23756 -20042
rect 20476 -20122 23756 -20102
rect 20476 -20142 20836 -20122
rect 20476 -22402 20756 -20142
rect 20816 -22402 20836 -20142
rect 20914 -20234 20948 -20218
rect 20914 -22226 20948 -22210
rect 21156 -20234 21316 -20122
rect 21156 -22210 21222 -20234
rect 21256 -22210 21316 -20234
rect 21156 -22222 21316 -22210
rect 21530 -20234 21564 -20218
rect 21222 -22226 21256 -22222
rect 21530 -22226 21564 -22210
rect 21776 -20234 21936 -20122
rect 21776 -22210 21838 -20234
rect 21872 -22210 21936 -20234
rect 21776 -22222 21936 -22210
rect 22146 -20234 22180 -20218
rect 21838 -22226 21872 -22222
rect 22146 -22226 22180 -22210
rect 22376 -20234 22536 -20122
rect 22376 -22210 22454 -20234
rect 22488 -22210 22536 -20234
rect 22376 -22222 22536 -22210
rect 22762 -20234 22796 -20218
rect 22454 -22226 22488 -22222
rect 22762 -22226 22796 -22210
rect 22996 -20234 23156 -20122
rect 23536 -20142 23756 -20122
rect 22996 -22210 23070 -20234
rect 23104 -22210 23156 -20234
rect 22996 -22222 23156 -22210
rect 23378 -20234 23412 -20218
rect 23070 -22226 23104 -22222
rect 23378 -22226 23412 -22210
rect 20960 -22303 20976 -22269
rect 21194 -22303 21210 -22269
rect 21268 -22303 21284 -22269
rect 21502 -22303 21518 -22269
rect 21576 -22303 21592 -22269
rect 21810 -22303 21826 -22269
rect 21884 -22303 21900 -22269
rect 22118 -22303 22134 -22269
rect 22192 -22303 22208 -22269
rect 22426 -22303 22442 -22269
rect 22500 -22303 22516 -22269
rect 22734 -22303 22750 -22269
rect 22808 -22303 22824 -22269
rect 23042 -22303 23058 -22269
rect 23116 -22303 23132 -22269
rect 23350 -22303 23366 -22269
rect 20476 -22422 20836 -22402
rect 23536 -22402 23556 -20142
rect 23616 -21922 23756 -20142
rect 23816 -21922 23836 -19762
rect 23916 -19858 23976 -19742
rect 24076 -19858 24136 -19742
rect 24236 -19858 24296 -19742
rect 23914 -19874 23976 -19858
rect 23948 -21730 23976 -19874
rect 23914 -21746 23976 -21730
rect 24072 -19874 24136 -19858
rect 24106 -21730 24136 -19874
rect 24072 -21746 24136 -21730
rect 24230 -19874 24296 -19858
rect 24264 -21730 24296 -19874
rect 24356 -20049 24496 -19862
rect 24349 -20065 24496 -20049
rect 24383 -21549 24496 -20065
rect 24349 -21565 24496 -21549
rect 24230 -21746 24296 -21730
rect 23916 -21782 23976 -21746
rect 24076 -21782 24136 -21746
rect 24236 -21782 24296 -21746
rect 23916 -21789 24296 -21782
rect 23916 -21823 23976 -21789
rect 24044 -21823 24134 -21789
rect 24202 -21823 24296 -21789
rect 23916 -21842 24296 -21823
rect 24356 -21782 24496 -21565
rect 24596 -20065 24736 -19742
rect 24596 -21549 24657 -20065
rect 24691 -21549 24736 -20065
rect 24596 -21642 24736 -21549
rect 24965 -20065 24999 -20049
rect 24965 -21565 24999 -21549
rect 25216 -20065 25356 -19742
rect 25216 -21549 25273 -20065
rect 25307 -21549 25356 -20065
rect 25216 -21642 25356 -21549
rect 25516 -20065 25656 -19862
rect 25516 -21549 25581 -20065
rect 25615 -21549 25656 -20065
rect 25516 -21782 25656 -21549
rect 25836 -20065 25976 -19742
rect 25836 -21549 25889 -20065
rect 25923 -21549 25976 -20065
rect 25836 -21642 25976 -21549
rect 26197 -20065 26231 -20049
rect 26197 -21565 26231 -21549
rect 26456 -20065 26596 -19742
rect 26456 -21549 26505 -20065
rect 26539 -21549 26596 -20065
rect 26456 -21642 26596 -21549
rect 26756 -20065 26896 -19862
rect 26756 -21549 26813 -20065
rect 26847 -21549 26896 -20065
rect 26756 -21782 26896 -21549
rect 27076 -20065 27216 -19742
rect 27076 -21549 27121 -20065
rect 27155 -21549 27216 -20065
rect 27076 -21642 27216 -21549
rect 27429 -20065 27463 -20049
rect 27429 -21565 27463 -21549
rect 27676 -20065 27816 -19742
rect 27676 -21549 27737 -20065
rect 27771 -21549 27816 -20065
rect 27676 -21622 27816 -21549
rect 27976 -20065 28116 -19862
rect 27976 -21549 28045 -20065
rect 28079 -21549 28116 -20065
rect 27976 -21782 28116 -21549
rect 28296 -20065 28436 -19742
rect 28296 -21549 28353 -20065
rect 28387 -21549 28436 -20065
rect 28296 -21622 28436 -21549
rect 28661 -20065 28695 -20049
rect 28661 -21565 28695 -21549
rect 28916 -20065 29056 -19742
rect 29416 -19858 29476 -19742
rect 29576 -19858 29636 -19742
rect 29736 -19858 29796 -19742
rect 29936 -19762 30196 -19742
rect 28916 -21549 28969 -20065
rect 29003 -21549 29056 -20065
rect 28916 -21622 29056 -21549
rect 29216 -20065 29356 -19862
rect 29216 -21549 29277 -20065
rect 29311 -21549 29356 -20065
rect 29216 -21782 29356 -21549
rect 24356 -21794 29356 -21782
rect 24356 -21828 24411 -21794
rect 24629 -21828 24719 -21794
rect 24937 -21828 25027 -21794
rect 25245 -21828 25335 -21794
rect 25553 -21828 25643 -21794
rect 25861 -21828 25951 -21794
rect 26169 -21828 26259 -21794
rect 26477 -21828 26567 -21794
rect 26785 -21828 26875 -21794
rect 27093 -21828 27183 -21794
rect 27401 -21828 27491 -21794
rect 27709 -21828 27799 -21794
rect 28017 -21828 28107 -21794
rect 28325 -21828 28415 -21794
rect 28633 -21828 28723 -21794
rect 28941 -21828 29031 -21794
rect 29249 -21828 29356 -21794
rect 24356 -21842 29356 -21828
rect 29416 -19874 29488 -19858
rect 29416 -21730 29454 -19874
rect 29416 -21746 29488 -21730
rect 29576 -19874 29646 -19858
rect 29576 -21730 29612 -19874
rect 29576 -21746 29646 -21730
rect 29736 -19874 29804 -19858
rect 29736 -21730 29770 -19874
rect 29736 -21746 29804 -21730
rect 29416 -21782 29476 -21746
rect 29576 -21782 29636 -21746
rect 29736 -21782 29796 -21746
rect 29416 -21789 29796 -21782
rect 29416 -21823 29516 -21789
rect 29584 -21823 29674 -21789
rect 29742 -21823 29796 -21789
rect 29416 -21842 29796 -21823
rect 23616 -21942 23836 -21922
rect 29936 -21922 29956 -19762
rect 30016 -19802 30196 -19762
rect 30316 -19622 30356 -18662
rect 30316 -19642 33496 -19622
rect 30316 -19802 30356 -19642
rect 33276 -19802 33496 -19642
rect 30016 -19842 33496 -19802
rect 30016 -20042 33316 -19842
rect 30016 -20102 30256 -20042
rect 32916 -20102 33316 -20042
rect 30016 -20122 33316 -20102
rect 30016 -20142 30236 -20122
rect 30016 -21922 30156 -20142
rect 29936 -21942 30156 -21922
rect 23616 -21962 30156 -21942
rect 23616 -22022 23856 -21962
rect 29916 -22022 30156 -21962
rect 23616 -22402 30156 -22022
rect 30216 -22402 30236 -20142
rect 30354 -20234 30388 -20218
rect 30354 -22226 30388 -22210
rect 30616 -20234 30776 -20122
rect 30616 -22210 30662 -20234
rect 30696 -22210 30776 -20234
rect 30616 -22222 30776 -22210
rect 30970 -20234 31004 -20218
rect 30662 -22226 30696 -22222
rect 30970 -22226 31004 -22210
rect 31216 -20234 31376 -20122
rect 31216 -22210 31278 -20234
rect 31312 -22210 31376 -20234
rect 31216 -22222 31376 -22210
rect 31586 -20234 31620 -20218
rect 31278 -22226 31312 -22222
rect 31586 -22226 31620 -22210
rect 31836 -20234 31996 -20122
rect 31836 -22210 31894 -20234
rect 31928 -22210 31996 -20234
rect 31836 -22222 31996 -22210
rect 32202 -20234 32236 -20218
rect 31894 -22226 31928 -22222
rect 32202 -22226 32236 -22210
rect 32436 -20234 32596 -20122
rect 32936 -20142 33316 -20122
rect 32436 -22210 32510 -20234
rect 32544 -22210 32596 -20234
rect 32436 -22222 32596 -22210
rect 32818 -20234 32852 -20218
rect 32510 -22226 32544 -22222
rect 32818 -22226 32852 -22210
rect 30400 -22303 30416 -22269
rect 30634 -22303 30650 -22269
rect 30708 -22303 30724 -22269
rect 30942 -22303 30958 -22269
rect 31016 -22303 31032 -22269
rect 31250 -22303 31266 -22269
rect 31324 -22303 31340 -22269
rect 31558 -22303 31574 -22269
rect 31632 -22303 31648 -22269
rect 31866 -22303 31882 -22269
rect 31940 -22303 31956 -22269
rect 32174 -22303 32190 -22269
rect 32248 -22303 32264 -22269
rect 32482 -22303 32498 -22269
rect 32556 -22303 32572 -22269
rect 32790 -22303 32806 -22269
rect 23536 -22422 30236 -22402
rect 32936 -22402 32956 -20142
rect 33016 -22402 33316 -20142
rect 32936 -22422 33316 -22402
rect 20476 -22442 33316 -22422
rect 20476 -22502 20856 -22442
rect 23516 -22502 30256 -22442
rect 32916 -22502 33316 -22442
rect 20476 -22582 33316 -22502
rect 20476 -22742 22756 -22582
rect 20476 -22802 21716 -22742
rect 22476 -22802 22756 -22742
rect 20476 -22822 22756 -22802
rect 20476 -22842 21696 -22822
rect 20476 -24102 21616 -22842
rect 21676 -24102 21696 -22842
rect 22496 -22842 22756 -22822
rect 21874 -22934 21908 -22918
rect 21874 -23926 21908 -23910
rect 22112 -22934 22146 -22918
rect 22112 -23926 22146 -23910
rect 22350 -22934 22384 -22918
rect 22350 -23926 22384 -23910
rect 21920 -24003 21936 -23969
rect 22084 -24003 22100 -23969
rect 22158 -24003 22174 -23969
rect 22322 -24003 22338 -23969
rect 20476 -24122 21696 -24102
rect 22496 -24102 22516 -22842
rect 22576 -24102 22756 -22842
rect 22496 -24122 22756 -24102
rect 20476 -24142 22756 -24122
rect 20476 -24202 21716 -24142
rect 22476 -24202 22756 -24142
rect 20476 -24322 22756 -24202
rect 22796 -22742 30996 -22622
rect 22796 -22802 23116 -22742
rect 30676 -22802 30996 -22742
rect 22796 -22822 30996 -22802
rect 22796 -22842 26596 -22822
rect 20476 -28202 20496 -24322
rect 22796 -24362 23016 -22842
rect 20536 -24402 23016 -24362
rect 20536 -24482 21936 -24402
rect 22016 -24482 22076 -24402
rect 22176 -24482 22236 -24402
rect 22316 -24482 23016 -24402
rect 20536 -24562 23016 -24482
rect 20536 -24622 21336 -24562
rect 22796 -24622 23016 -24562
rect 20536 -24642 23016 -24622
rect 20536 -24662 21316 -24642
rect 20536 -26422 21236 -24662
rect 21296 -26422 21316 -24662
rect 21428 -24766 21462 -24750
rect 21676 -24766 21836 -24642
rect 21676 -26242 21736 -24766
rect 21770 -26242 21836 -24766
rect 22044 -24766 22078 -24750
rect 22296 -24766 22456 -24642
rect 22816 -24662 23016 -24642
rect 22296 -26242 22352 -24766
rect 22386 -26242 22456 -24766
rect 22660 -24766 22694 -24750
rect 21428 -26258 21462 -26242
rect 21736 -26258 21770 -26242
rect 22044 -26258 22078 -26242
rect 22352 -26258 22386 -26242
rect 22660 -26258 22694 -26242
rect 21474 -26326 21490 -26292
rect 21708 -26326 21724 -26292
rect 21782 -26326 21798 -26292
rect 22016 -26326 22032 -26292
rect 22090 -26326 22106 -26292
rect 22324 -26326 22340 -26292
rect 22398 -26326 22414 -26292
rect 22632 -26326 22648 -26292
rect 20536 -26442 21316 -26422
rect 22816 -26422 22836 -24662
rect 22896 -26102 23016 -24662
rect 23076 -22942 26596 -22842
rect 27196 -22842 30996 -22822
rect 23076 -23002 23236 -22942
rect 24756 -23002 25036 -22942
rect 26556 -23002 26596 -22942
rect 23076 -23022 26596 -23002
rect 26636 -22922 27156 -22862
rect 26636 -23002 26716 -22922
rect 26796 -23002 26856 -22922
rect 26936 -23002 26996 -22922
rect 27076 -23002 27156 -22922
rect 23076 -25922 23156 -23022
rect 23356 -23156 23416 -23022
rect 23356 -24082 23368 -23156
rect 23402 -24082 23416 -23156
rect 23356 -24102 23416 -24082
rect 23516 -23156 23576 -23022
rect 23516 -24082 23526 -23156
rect 23560 -24082 23576 -23156
rect 23516 -24102 23576 -24082
rect 23676 -23156 23736 -23022
rect 23676 -24082 23684 -23156
rect 23718 -24082 23736 -23156
rect 23676 -24102 23736 -24082
rect 23808 -23156 23842 -23140
rect 23808 -24098 23842 -24082
rect 23966 -23156 24000 -23140
rect 23966 -24098 24000 -24082
rect 24124 -23156 24158 -23140
rect 24124 -24098 24158 -24082
rect 24236 -23156 24296 -23022
rect 24236 -24082 24248 -23156
rect 24282 -24082 24296 -23156
rect 23356 -24132 23736 -24102
rect 24236 -24102 24296 -24082
rect 24396 -23156 24456 -23022
rect 24396 -24082 24406 -23156
rect 24440 -24082 24456 -23156
rect 24396 -24102 24456 -24082
rect 24556 -23156 24616 -23022
rect 24556 -24082 24564 -23156
rect 24598 -24082 24616 -23156
rect 24556 -24102 24616 -24082
rect 24236 -24132 24616 -24102
rect 23356 -24166 23430 -24132
rect 23498 -24166 23588 -24132
rect 23656 -24166 23736 -24132
rect 23854 -24166 23870 -24132
rect 23938 -24166 23954 -24132
rect 24012 -24166 24028 -24132
rect 24096 -24166 24112 -24132
rect 24236 -24166 24310 -24132
rect 24378 -24166 24468 -24132
rect 24536 -24166 24616 -24132
rect 23356 -24182 23736 -24166
rect 24236 -24182 24616 -24166
rect 24796 -23082 24996 -23062
rect 24796 -23162 24856 -23082
rect 24936 -23162 24996 -23082
rect 24796 -23202 24996 -23162
rect 24796 -23282 24856 -23202
rect 24936 -23282 24996 -23202
rect 24796 -23322 24996 -23282
rect 24796 -23402 24856 -23322
rect 24936 -23402 24996 -23322
rect 24796 -23442 24996 -23402
rect 24796 -23522 24856 -23442
rect 24936 -23522 24996 -23442
rect 24796 -23562 24996 -23522
rect 24796 -23642 24856 -23562
rect 24936 -23642 24996 -23562
rect 24796 -23682 24996 -23642
rect 24796 -23762 24856 -23682
rect 24936 -23762 24996 -23682
rect 24796 -23802 24996 -23762
rect 24796 -23882 24856 -23802
rect 24936 -23882 24996 -23802
rect 24796 -23922 24996 -23882
rect 24796 -24002 24856 -23922
rect 24936 -24002 24996 -23922
rect 24796 -24042 24996 -24002
rect 24796 -24122 24856 -24042
rect 24936 -24122 24996 -24042
rect 24796 -24162 24996 -24122
rect 24796 -24242 24856 -24162
rect 24936 -24242 24996 -24162
rect 25156 -23156 25216 -23022
rect 25156 -24082 25168 -23156
rect 25202 -24082 25216 -23156
rect 25156 -24102 25216 -24082
rect 25316 -23156 25376 -23022
rect 25316 -24082 25326 -23156
rect 25360 -24082 25376 -23156
rect 25316 -24102 25376 -24082
rect 25476 -23156 25536 -23022
rect 25476 -24082 25484 -23156
rect 25518 -24082 25536 -23156
rect 25476 -24102 25536 -24082
rect 25608 -23156 25642 -23140
rect 25608 -24098 25642 -24082
rect 25766 -23156 25800 -23140
rect 25766 -24098 25800 -24082
rect 25924 -23156 25958 -23140
rect 25924 -24098 25958 -24082
rect 26036 -23156 26096 -23022
rect 26036 -24082 26048 -23156
rect 26082 -24082 26096 -23156
rect 25156 -24132 25536 -24102
rect 26036 -24102 26096 -24082
rect 26196 -23156 26256 -23022
rect 26196 -24082 26206 -23156
rect 26240 -24082 26256 -23156
rect 26196 -24102 26256 -24082
rect 26356 -23156 26416 -23022
rect 26356 -24082 26364 -23156
rect 26398 -24082 26416 -23156
rect 26356 -24102 26416 -24082
rect 26036 -24132 26416 -24102
rect 25156 -24166 25230 -24132
rect 25298 -24166 25388 -24132
rect 25456 -24166 25536 -24132
rect 25654 -24166 25670 -24132
rect 25738 -24166 25754 -24132
rect 25812 -24166 25828 -24132
rect 25896 -24166 25912 -24132
rect 26036 -24166 26110 -24132
rect 26178 -24166 26268 -24132
rect 26336 -24166 26416 -24132
rect 25156 -24182 25536 -24166
rect 26036 -24182 26416 -24166
rect 26636 -23042 27156 -23002
rect 27196 -22942 30716 -22842
rect 27196 -23002 27236 -22942
rect 28756 -23002 29036 -22942
rect 30556 -23002 30716 -22942
rect 27196 -23022 30716 -23002
rect 26636 -23122 26716 -23042
rect 26796 -23122 26856 -23042
rect 26936 -23122 26996 -23042
rect 27076 -23122 27156 -23042
rect 26636 -23162 27156 -23122
rect 26636 -23242 26716 -23162
rect 26796 -23242 26856 -23162
rect 26936 -23242 26996 -23162
rect 27076 -23242 27156 -23162
rect 26636 -23282 27156 -23242
rect 26636 -23362 26716 -23282
rect 26796 -23362 26856 -23282
rect 26936 -23362 26996 -23282
rect 27076 -23362 27156 -23282
rect 26636 -23402 27156 -23362
rect 26636 -23482 26716 -23402
rect 26796 -23482 26856 -23402
rect 26936 -23482 26996 -23402
rect 27076 -23482 27156 -23402
rect 26636 -23522 27156 -23482
rect 26636 -23602 26716 -23522
rect 26796 -23602 26856 -23522
rect 26936 -23602 26996 -23522
rect 27076 -23602 27156 -23522
rect 26636 -23642 27156 -23602
rect 26636 -23722 26716 -23642
rect 26796 -23722 26856 -23642
rect 26936 -23722 26996 -23642
rect 27076 -23722 27156 -23642
rect 26636 -23762 27156 -23722
rect 26636 -23842 26716 -23762
rect 26796 -23842 26856 -23762
rect 26936 -23842 26996 -23762
rect 27076 -23842 27156 -23762
rect 26636 -23882 27156 -23842
rect 26636 -23962 26716 -23882
rect 26796 -23962 26856 -23882
rect 26936 -23962 26996 -23882
rect 27076 -23962 27156 -23882
rect 26636 -24002 27156 -23962
rect 26636 -24082 26716 -24002
rect 26796 -24082 26856 -24002
rect 26936 -24082 26996 -24002
rect 27076 -24082 27156 -24002
rect 26636 -24122 27156 -24082
rect 24796 -24282 24996 -24242
rect 24796 -24322 24856 -24282
rect 23196 -24362 24856 -24322
rect 24936 -24322 24996 -24282
rect 26636 -24202 26716 -24122
rect 26796 -24202 26856 -24122
rect 26936 -24202 26996 -24122
rect 27076 -24202 27156 -24122
rect 27356 -23156 27416 -23022
rect 27356 -24082 27368 -23156
rect 27402 -24082 27416 -23156
rect 27356 -24102 27416 -24082
rect 27516 -23156 27576 -23022
rect 27516 -24082 27526 -23156
rect 27560 -24082 27576 -23156
rect 27516 -24102 27576 -24082
rect 27676 -23156 27736 -23022
rect 27676 -24082 27684 -23156
rect 27718 -24082 27736 -23156
rect 27676 -24102 27736 -24082
rect 27808 -23156 27842 -23140
rect 27808 -24098 27842 -24082
rect 27966 -23156 28000 -23140
rect 27966 -24098 28000 -24082
rect 28124 -23156 28158 -23140
rect 28124 -24098 28158 -24082
rect 28236 -23156 28296 -23022
rect 28236 -24082 28248 -23156
rect 28282 -24082 28296 -23156
rect 27356 -24132 27736 -24102
rect 28236 -24102 28296 -24082
rect 28396 -23156 28456 -23022
rect 28396 -24082 28406 -23156
rect 28440 -24082 28456 -23156
rect 28396 -24102 28456 -24082
rect 28556 -23156 28616 -23022
rect 28556 -24082 28564 -23156
rect 28598 -24082 28616 -23156
rect 28556 -24102 28616 -24082
rect 28236 -24132 28616 -24102
rect 27356 -24166 27430 -24132
rect 27498 -24166 27588 -24132
rect 27656 -24166 27736 -24132
rect 27854 -24166 27870 -24132
rect 27938 -24166 27954 -24132
rect 28012 -24166 28028 -24132
rect 28096 -24166 28112 -24132
rect 28236 -24166 28310 -24132
rect 28378 -24166 28468 -24132
rect 28536 -24166 28616 -24132
rect 27356 -24182 27736 -24166
rect 28236 -24182 28616 -24166
rect 28796 -23082 28996 -23062
rect 28796 -23162 28856 -23082
rect 28936 -23162 28996 -23082
rect 28796 -23202 28996 -23162
rect 28796 -23282 28856 -23202
rect 28936 -23282 28996 -23202
rect 28796 -23322 28996 -23282
rect 28796 -23402 28856 -23322
rect 28936 -23402 28996 -23322
rect 28796 -23442 28996 -23402
rect 28796 -23522 28856 -23442
rect 28936 -23522 28996 -23442
rect 28796 -23562 28996 -23522
rect 28796 -23642 28856 -23562
rect 28936 -23642 28996 -23562
rect 28796 -23682 28996 -23642
rect 28796 -23762 28856 -23682
rect 28936 -23762 28996 -23682
rect 28796 -23802 28996 -23762
rect 28796 -23882 28856 -23802
rect 28936 -23882 28996 -23802
rect 28796 -23922 28996 -23882
rect 28796 -24002 28856 -23922
rect 28936 -24002 28996 -23922
rect 28796 -24042 28996 -24002
rect 28796 -24122 28856 -24042
rect 28936 -24122 28996 -24042
rect 28796 -24162 28996 -24122
rect 26636 -24242 27156 -24202
rect 26636 -24322 26716 -24242
rect 26796 -24322 26856 -24242
rect 26936 -24322 26996 -24242
rect 27076 -24322 27156 -24242
rect 28796 -24242 28856 -24162
rect 28936 -24242 28996 -24162
rect 29156 -23156 29216 -23022
rect 29156 -24082 29168 -23156
rect 29202 -24082 29216 -23156
rect 29156 -24102 29216 -24082
rect 29316 -23156 29376 -23022
rect 29316 -24082 29326 -23156
rect 29360 -24082 29376 -23156
rect 29316 -24102 29376 -24082
rect 29476 -23156 29536 -23022
rect 29476 -24082 29484 -23156
rect 29518 -24082 29536 -23156
rect 29476 -24102 29536 -24082
rect 29608 -23156 29642 -23140
rect 29608 -24098 29642 -24082
rect 29766 -23156 29800 -23140
rect 29766 -24098 29800 -24082
rect 29924 -23156 29958 -23140
rect 29924 -24098 29958 -24082
rect 30036 -23156 30096 -23022
rect 30036 -24082 30048 -23156
rect 30082 -24082 30096 -23156
rect 29156 -24132 29536 -24102
rect 30036 -24102 30096 -24082
rect 30196 -23156 30256 -23022
rect 30196 -24082 30206 -23156
rect 30240 -24082 30256 -23156
rect 30196 -24102 30256 -24082
rect 30356 -23156 30416 -23022
rect 30356 -24082 30364 -23156
rect 30398 -24082 30416 -23156
rect 30356 -24102 30416 -24082
rect 30036 -24132 30416 -24102
rect 29156 -24166 29230 -24132
rect 29298 -24166 29388 -24132
rect 29456 -24166 29536 -24132
rect 29654 -24166 29670 -24132
rect 29738 -24166 29754 -24132
rect 29812 -24166 29828 -24132
rect 29896 -24166 29912 -24132
rect 30036 -24166 30110 -24132
rect 30178 -24166 30268 -24132
rect 30336 -24166 30416 -24132
rect 29156 -24182 29536 -24166
rect 30036 -24182 30416 -24166
rect 28796 -24282 28996 -24242
rect 28796 -24322 28856 -24282
rect 24936 -24362 28856 -24322
rect 28936 -24322 28996 -24282
rect 28936 -24362 30596 -24322
rect 23196 -24442 23236 -24362
rect 23316 -24442 23356 -24362
rect 23436 -24442 23476 -24362
rect 23556 -24442 23596 -24362
rect 23676 -24442 23716 -24362
rect 23796 -24442 23836 -24362
rect 23916 -24442 23956 -24362
rect 24036 -24442 24076 -24362
rect 24156 -24442 24196 -24362
rect 24276 -24442 24316 -24362
rect 24396 -24442 24436 -24362
rect 24516 -24442 24556 -24362
rect 24636 -24442 24676 -24362
rect 24756 -24402 25036 -24362
rect 24756 -24442 24856 -24402
rect 23196 -24482 24856 -24442
rect 24936 -24442 25036 -24402
rect 25116 -24442 25156 -24362
rect 25236 -24442 25276 -24362
rect 25356 -24442 25396 -24362
rect 25476 -24442 25516 -24362
rect 25596 -24442 25636 -24362
rect 25716 -24442 25756 -24362
rect 25836 -24442 25876 -24362
rect 25956 -24442 25996 -24362
rect 26076 -24442 26116 -24362
rect 26196 -24442 26236 -24362
rect 26316 -24442 26356 -24362
rect 26436 -24442 26476 -24362
rect 26556 -24442 26596 -24362
rect 26676 -24442 26716 -24362
rect 26796 -24442 26856 -24362
rect 26936 -24442 26996 -24362
rect 27076 -24442 27116 -24362
rect 27196 -24442 27236 -24362
rect 27316 -24442 27356 -24362
rect 27436 -24442 27476 -24362
rect 27556 -24442 27596 -24362
rect 27676 -24442 27716 -24362
rect 27796 -24442 27836 -24362
rect 27916 -24442 27956 -24362
rect 28036 -24442 28076 -24362
rect 28156 -24442 28196 -24362
rect 28276 -24442 28316 -24362
rect 28396 -24442 28436 -24362
rect 28516 -24442 28556 -24362
rect 28636 -24442 28676 -24362
rect 28756 -24402 29036 -24362
rect 28756 -24442 28856 -24402
rect 24936 -24482 28856 -24442
rect 28936 -24442 29036 -24402
rect 29116 -24442 29156 -24362
rect 29236 -24442 29276 -24362
rect 29356 -24442 29396 -24362
rect 29476 -24442 29516 -24362
rect 29596 -24442 29636 -24362
rect 29716 -24442 29756 -24362
rect 29836 -24442 29876 -24362
rect 29956 -24442 29996 -24362
rect 30076 -24442 30116 -24362
rect 30196 -24442 30236 -24362
rect 30316 -24442 30356 -24362
rect 30436 -24442 30476 -24362
rect 30556 -24442 30596 -24362
rect 28936 -24482 30596 -24442
rect 23196 -24502 26716 -24482
rect 23196 -24582 23236 -24502
rect 23316 -24582 23356 -24502
rect 23436 -24582 23476 -24502
rect 23556 -24582 23596 -24502
rect 23676 -24582 23716 -24502
rect 23796 -24582 23836 -24502
rect 23916 -24582 23956 -24502
rect 24036 -24582 24076 -24502
rect 24156 -24582 24196 -24502
rect 24276 -24582 24316 -24502
rect 24396 -24582 24436 -24502
rect 24516 -24582 24556 -24502
rect 24636 -24582 24676 -24502
rect 24756 -24522 25036 -24502
rect 24756 -24582 24856 -24522
rect 23196 -24602 24856 -24582
rect 24936 -24582 25036 -24522
rect 25116 -24582 25156 -24502
rect 25236 -24582 25276 -24502
rect 25356 -24582 25396 -24502
rect 25476 -24582 25516 -24502
rect 25596 -24582 25636 -24502
rect 25716 -24582 25756 -24502
rect 25836 -24582 25876 -24502
rect 25956 -24582 25996 -24502
rect 26076 -24582 26116 -24502
rect 26196 -24582 26236 -24502
rect 26316 -24582 26356 -24502
rect 26436 -24582 26476 -24502
rect 26556 -24582 26596 -24502
rect 26676 -24562 26716 -24502
rect 26796 -24562 26856 -24482
rect 26936 -24562 26996 -24482
rect 27076 -24502 30596 -24482
rect 27076 -24562 27116 -24502
rect 26676 -24582 27116 -24562
rect 27196 -24582 27236 -24502
rect 27316 -24582 27356 -24502
rect 27436 -24582 27476 -24502
rect 27556 -24582 27596 -24502
rect 27676 -24582 27716 -24502
rect 27796 -24582 27836 -24502
rect 27916 -24582 27956 -24502
rect 28036 -24582 28076 -24502
rect 28156 -24582 28196 -24502
rect 28276 -24582 28316 -24502
rect 28396 -24582 28436 -24502
rect 28516 -24582 28556 -24502
rect 28636 -24582 28676 -24502
rect 28756 -24522 29036 -24502
rect 28756 -24582 28856 -24522
rect 24936 -24602 28856 -24582
rect 28936 -24582 29036 -24522
rect 29116 -24582 29156 -24502
rect 29236 -24582 29276 -24502
rect 29356 -24582 29396 -24502
rect 29476 -24582 29516 -24502
rect 29596 -24582 29636 -24502
rect 29716 -24582 29756 -24502
rect 29836 -24582 29876 -24502
rect 29956 -24582 29996 -24502
rect 30076 -24582 30116 -24502
rect 30196 -24582 30236 -24502
rect 30316 -24582 30356 -24502
rect 30436 -24582 30476 -24502
rect 30556 -24582 30596 -24502
rect 28936 -24602 30596 -24582
rect 23196 -24622 26716 -24602
rect 24796 -24642 24996 -24622
rect 24796 -24722 24856 -24642
rect 24936 -24722 24996 -24642
rect 24796 -24762 24996 -24722
rect 26636 -24682 26716 -24622
rect 26796 -24682 26856 -24602
rect 26936 -24682 26996 -24602
rect 27076 -24622 30596 -24602
rect 27076 -24682 27156 -24622
rect 26636 -24722 27156 -24682
rect 23356 -24774 23736 -24762
rect 24236 -24774 24616 -24762
rect 23356 -24808 23430 -24774
rect 23498 -24808 23588 -24774
rect 23656 -24808 23736 -24774
rect 23854 -24808 23870 -24774
rect 23938 -24808 23954 -24774
rect 24012 -24808 24028 -24774
rect 24096 -24808 24112 -24774
rect 24236 -24808 24310 -24774
rect 24378 -24808 24468 -24774
rect 24536 -24808 24616 -24774
rect 23356 -24842 23736 -24808
rect 24236 -24842 24616 -24808
rect 23356 -24858 23416 -24842
rect 23356 -25784 23368 -24858
rect 23402 -25784 23416 -24858
rect 23356 -25922 23416 -25784
rect 23516 -24858 23576 -24842
rect 23516 -25784 23526 -24858
rect 23560 -25784 23576 -24858
rect 23516 -25922 23576 -25784
rect 23676 -24858 23736 -24842
rect 23676 -25784 23684 -24858
rect 23718 -25784 23736 -24858
rect 23676 -25922 23736 -25784
rect 23808 -24858 23842 -24842
rect 23808 -25800 23842 -25784
rect 23966 -24858 24000 -24842
rect 23966 -25800 24000 -25784
rect 24124 -24858 24158 -24842
rect 24124 -25800 24158 -25784
rect 24236 -24858 24296 -24842
rect 24236 -25784 24248 -24858
rect 24282 -25784 24296 -24858
rect 24236 -25922 24296 -25784
rect 24396 -24858 24456 -24842
rect 24396 -25784 24406 -24858
rect 24440 -25784 24456 -24858
rect 24396 -25922 24456 -25784
rect 24556 -24858 24616 -24842
rect 24556 -25784 24564 -24858
rect 24598 -25784 24616 -24858
rect 24556 -25922 24616 -25784
rect 24796 -24842 24856 -24762
rect 24936 -24842 24996 -24762
rect 24796 -24882 24996 -24842
rect 24796 -24962 24856 -24882
rect 24936 -24962 24996 -24882
rect 24796 -25002 24996 -24962
rect 24796 -25082 24856 -25002
rect 24936 -25082 24996 -25002
rect 24796 -25122 24996 -25082
rect 24796 -25202 24856 -25122
rect 24936 -25202 24996 -25122
rect 24796 -25242 24996 -25202
rect 24796 -25322 24856 -25242
rect 24936 -25322 24996 -25242
rect 24796 -25362 24996 -25322
rect 24796 -25442 24856 -25362
rect 24936 -25442 24996 -25362
rect 24796 -25482 24996 -25442
rect 24796 -25562 24856 -25482
rect 24936 -25562 24996 -25482
rect 24796 -25602 24996 -25562
rect 24796 -25682 24856 -25602
rect 24936 -25682 24996 -25602
rect 24796 -25722 24996 -25682
rect 24796 -25802 24856 -25722
rect 24936 -25802 24996 -25722
rect 24796 -25882 24996 -25802
rect 25156 -24774 25536 -24762
rect 26036 -24774 26416 -24762
rect 25156 -24808 25230 -24774
rect 25298 -24808 25388 -24774
rect 25456 -24808 25536 -24774
rect 25654 -24808 25670 -24774
rect 25738 -24808 25754 -24774
rect 25812 -24808 25828 -24774
rect 25896 -24808 25912 -24774
rect 26036 -24808 26110 -24774
rect 26178 -24808 26268 -24774
rect 26336 -24808 26416 -24774
rect 25156 -24842 25536 -24808
rect 26036 -24842 26416 -24808
rect 25156 -24858 25216 -24842
rect 25156 -25784 25168 -24858
rect 25202 -25784 25216 -24858
rect 25156 -25922 25216 -25784
rect 25316 -24858 25376 -24842
rect 25316 -25784 25326 -24858
rect 25360 -25784 25376 -24858
rect 25316 -25922 25376 -25784
rect 25476 -24858 25536 -24842
rect 25476 -25784 25484 -24858
rect 25518 -25784 25536 -24858
rect 25476 -25922 25536 -25784
rect 25608 -24858 25642 -24842
rect 25608 -25800 25642 -25784
rect 25766 -24858 25800 -24842
rect 25766 -25800 25800 -25784
rect 25924 -24858 25958 -24842
rect 25924 -25800 25958 -25784
rect 26036 -24858 26096 -24842
rect 26036 -25784 26048 -24858
rect 26082 -25784 26096 -24858
rect 26036 -25922 26096 -25784
rect 26196 -24858 26256 -24842
rect 26196 -25784 26206 -24858
rect 26240 -25784 26256 -24858
rect 26196 -25922 26256 -25784
rect 26356 -24858 26416 -24842
rect 26356 -25784 26364 -24858
rect 26398 -25784 26416 -24858
rect 26356 -25922 26416 -25784
rect 26636 -24802 26716 -24722
rect 26796 -24802 26856 -24722
rect 26936 -24802 26996 -24722
rect 27076 -24802 27156 -24722
rect 28796 -24642 28996 -24622
rect 28796 -24722 28856 -24642
rect 28936 -24722 28996 -24642
rect 28796 -24762 28996 -24722
rect 26636 -24842 27156 -24802
rect 26636 -24922 26716 -24842
rect 26796 -24922 26856 -24842
rect 26936 -24922 26996 -24842
rect 27076 -24922 27156 -24842
rect 26636 -24962 27156 -24922
rect 26636 -25042 26716 -24962
rect 26796 -25042 26856 -24962
rect 26936 -25042 26996 -24962
rect 27076 -25042 27156 -24962
rect 26636 -25082 27156 -25042
rect 26636 -25162 26716 -25082
rect 26796 -25162 26856 -25082
rect 26936 -25162 26996 -25082
rect 27076 -25162 27156 -25082
rect 26636 -25202 27156 -25162
rect 26636 -25282 26716 -25202
rect 26796 -25282 26856 -25202
rect 26936 -25282 26996 -25202
rect 27076 -25282 27156 -25202
rect 26636 -25322 27156 -25282
rect 26636 -25402 26716 -25322
rect 26796 -25402 26856 -25322
rect 26936 -25402 26996 -25322
rect 27076 -25402 27156 -25322
rect 26636 -25442 27156 -25402
rect 26636 -25522 26716 -25442
rect 26796 -25522 26856 -25442
rect 26936 -25522 26996 -25442
rect 27076 -25522 27156 -25442
rect 26636 -25562 27156 -25522
rect 26636 -25642 26716 -25562
rect 26796 -25642 26856 -25562
rect 26936 -25642 26996 -25562
rect 27076 -25642 27156 -25562
rect 26636 -25682 27156 -25642
rect 26636 -25762 26716 -25682
rect 26796 -25762 26856 -25682
rect 26936 -25762 26996 -25682
rect 27076 -25762 27156 -25682
rect 26636 -25802 27156 -25762
rect 26636 -25882 26716 -25802
rect 26796 -25882 26856 -25802
rect 26936 -25882 26996 -25802
rect 27076 -25882 27156 -25802
rect 26636 -25922 27156 -25882
rect 27356 -24774 27736 -24762
rect 28236 -24774 28616 -24762
rect 27356 -24808 27430 -24774
rect 27498 -24808 27588 -24774
rect 27656 -24808 27736 -24774
rect 27854 -24808 27870 -24774
rect 27938 -24808 27954 -24774
rect 28012 -24808 28028 -24774
rect 28096 -24808 28112 -24774
rect 28236 -24808 28310 -24774
rect 28378 -24808 28468 -24774
rect 28536 -24808 28616 -24774
rect 27356 -24842 27736 -24808
rect 28236 -24842 28616 -24808
rect 27356 -24858 27416 -24842
rect 27356 -25784 27368 -24858
rect 27402 -25784 27416 -24858
rect 27356 -25922 27416 -25784
rect 27516 -24858 27576 -24842
rect 27516 -25784 27526 -24858
rect 27560 -25784 27576 -24858
rect 27516 -25922 27576 -25784
rect 27676 -24858 27736 -24842
rect 27676 -25784 27684 -24858
rect 27718 -25784 27736 -24858
rect 27676 -25922 27736 -25784
rect 27808 -24858 27842 -24842
rect 27808 -25800 27842 -25784
rect 27966 -24858 28000 -24842
rect 27966 -25800 28000 -25784
rect 28124 -24858 28158 -24842
rect 28124 -25800 28158 -25784
rect 28236 -24858 28296 -24842
rect 28236 -25784 28248 -24858
rect 28282 -25784 28296 -24858
rect 28236 -25922 28296 -25784
rect 28396 -24858 28456 -24842
rect 28396 -25784 28406 -24858
rect 28440 -25784 28456 -24858
rect 28396 -25922 28456 -25784
rect 28556 -24858 28616 -24842
rect 28556 -25784 28564 -24858
rect 28598 -25784 28616 -24858
rect 28556 -25922 28616 -25784
rect 28796 -24842 28856 -24762
rect 28936 -24842 28996 -24762
rect 28796 -24882 28996 -24842
rect 28796 -24962 28856 -24882
rect 28936 -24962 28996 -24882
rect 28796 -25002 28996 -24962
rect 28796 -25082 28856 -25002
rect 28936 -25082 28996 -25002
rect 28796 -25122 28996 -25082
rect 28796 -25202 28856 -25122
rect 28936 -25202 28996 -25122
rect 28796 -25242 28996 -25202
rect 28796 -25322 28856 -25242
rect 28936 -25322 28996 -25242
rect 28796 -25362 28996 -25322
rect 28796 -25442 28856 -25362
rect 28936 -25442 28996 -25362
rect 28796 -25482 28996 -25442
rect 28796 -25562 28856 -25482
rect 28936 -25562 28996 -25482
rect 28796 -25602 28996 -25562
rect 28796 -25682 28856 -25602
rect 28936 -25682 28996 -25602
rect 28796 -25722 28996 -25682
rect 28796 -25802 28856 -25722
rect 28936 -25802 28996 -25722
rect 28796 -25882 28996 -25802
rect 29156 -24774 29536 -24762
rect 30036 -24774 30416 -24762
rect 29156 -24808 29230 -24774
rect 29298 -24808 29388 -24774
rect 29456 -24808 29536 -24774
rect 29654 -24808 29670 -24774
rect 29738 -24808 29754 -24774
rect 29812 -24808 29828 -24774
rect 29896 -24808 29912 -24774
rect 30036 -24808 30110 -24774
rect 30178 -24808 30268 -24774
rect 30336 -24808 30416 -24774
rect 29156 -24842 29536 -24808
rect 30036 -24842 30416 -24808
rect 29156 -24858 29216 -24842
rect 29156 -25784 29168 -24858
rect 29202 -25784 29216 -24858
rect 29156 -25922 29216 -25784
rect 29316 -24858 29376 -24842
rect 29316 -25784 29326 -24858
rect 29360 -25784 29376 -24858
rect 29316 -25922 29376 -25784
rect 29476 -24858 29536 -24842
rect 29476 -25784 29484 -24858
rect 29518 -25784 29536 -24858
rect 29476 -25922 29536 -25784
rect 29608 -24858 29642 -24842
rect 29608 -25800 29642 -25784
rect 29766 -24858 29800 -24842
rect 29766 -25800 29800 -25784
rect 29924 -24858 29958 -24842
rect 29924 -25800 29958 -25784
rect 30036 -24858 30096 -24842
rect 30036 -25784 30048 -24858
rect 30082 -25784 30096 -24858
rect 30036 -25922 30096 -25784
rect 30196 -24858 30256 -24842
rect 30196 -25784 30206 -24858
rect 30240 -25784 30256 -24858
rect 30196 -25922 30256 -25784
rect 30356 -24858 30416 -24842
rect 30356 -25784 30364 -24858
rect 30398 -25784 30416 -24858
rect 30356 -25922 30416 -25784
rect 30636 -25922 30716 -23022
rect 23076 -25942 26596 -25922
rect 23076 -26002 23236 -25942
rect 24756 -26002 25036 -25942
rect 26556 -26002 26596 -25942
rect 23076 -26102 26596 -26002
rect 26636 -26002 26716 -25922
rect 26796 -26002 26856 -25922
rect 26936 -26002 26996 -25922
rect 27076 -26002 27156 -25922
rect 26636 -26082 27156 -26002
rect 27196 -25942 30716 -25922
rect 27196 -26002 27236 -25942
rect 28756 -26002 29036 -25942
rect 30556 -26002 30716 -25942
rect 22896 -26122 26596 -26102
rect 27196 -26102 30716 -26002
rect 30776 -24362 30996 -22842
rect 31036 -22742 33316 -22582
rect 31036 -22802 31316 -22742
rect 32076 -22802 33316 -22742
rect 31036 -22822 33316 -22802
rect 31036 -22842 31296 -22822
rect 31036 -24102 31216 -22842
rect 31276 -24102 31296 -22842
rect 32096 -22842 33316 -22822
rect 31454 -22914 31488 -22898
rect 31454 -23906 31488 -23890
rect 31692 -22914 31726 -22898
rect 31692 -23906 31726 -23890
rect 31930 -22914 31964 -22898
rect 31930 -23906 31964 -23890
rect 31500 -23983 31516 -23949
rect 31664 -23983 31680 -23949
rect 31738 -23983 31754 -23949
rect 31902 -23983 31918 -23949
rect 31036 -24122 31296 -24102
rect 32096 -24102 32116 -22842
rect 32176 -24102 33316 -22842
rect 32096 -24122 33316 -24102
rect 31036 -24142 33316 -24122
rect 31036 -24202 31316 -24142
rect 32076 -24202 33316 -24142
rect 31036 -24322 33316 -24202
rect 30776 -24402 33256 -24362
rect 30776 -24482 31516 -24402
rect 31596 -24482 31636 -24402
rect 31776 -24482 31816 -24402
rect 31896 -24482 33256 -24402
rect 30776 -24582 33256 -24482
rect 30776 -24642 30996 -24582
rect 32456 -24642 33256 -24582
rect 30776 -24662 33256 -24642
rect 30776 -24682 30976 -24662
rect 30776 -26102 30896 -24682
rect 27196 -26122 30896 -26102
rect 22896 -26142 30896 -26122
rect 22896 -26202 23116 -26142
rect 30676 -26202 30896 -26142
rect 22896 -26222 30896 -26202
rect 22896 -26242 23796 -26222
rect 22896 -26422 23716 -26242
rect 22816 -26442 23716 -26422
rect 20536 -26462 23716 -26442
rect 20536 -26522 21336 -26462
rect 22796 -26522 23716 -26462
rect 20536 -28002 23716 -26522
rect 23776 -28002 23796 -26242
rect 29896 -26242 30896 -26222
rect 24376 -26302 29366 -26292
rect 20536 -28022 23796 -28002
rect 23936 -26324 24316 -26322
rect 23936 -26358 24010 -26324
rect 24078 -26358 24168 -26324
rect 24236 -26358 24316 -26324
rect 23936 -26402 24316 -26358
rect 23936 -26408 23996 -26402
rect 23936 -27884 23948 -26408
rect 23982 -27884 23996 -26408
rect 23936 -28022 23996 -27884
rect 24096 -26408 24156 -26402
rect 24096 -27884 24106 -26408
rect 24140 -27884 24156 -26408
rect 24096 -28022 24156 -27884
rect 24256 -26408 24316 -26402
rect 24256 -27884 24264 -26408
rect 24298 -27884 24316 -26408
rect 24256 -28022 24316 -27884
rect 24376 -26324 29376 -26302
rect 24376 -26358 24450 -26324
rect 24668 -26352 24758 -26324
rect 24668 -26358 24684 -26352
rect 24742 -26358 24758 -26352
rect 24976 -26352 25066 -26324
rect 24976 -26358 24992 -26352
rect 25050 -26358 25066 -26352
rect 25284 -26352 25374 -26324
rect 25284 -26358 25300 -26352
rect 25358 -26358 25374 -26352
rect 25592 -26358 25682 -26324
rect 25900 -26352 25990 -26324
rect 25900 -26358 25916 -26352
rect 25974 -26358 25990 -26352
rect 26208 -26352 26298 -26324
rect 26208 -26358 26224 -26352
rect 26282 -26358 26298 -26352
rect 26516 -26352 26606 -26324
rect 26516 -26358 26532 -26352
rect 26590 -26358 26606 -26352
rect 26824 -26358 26914 -26324
rect 27132 -26352 27222 -26324
rect 27132 -26358 27148 -26352
rect 27206 -26358 27222 -26352
rect 27440 -26352 27530 -26324
rect 27440 -26358 27456 -26352
rect 27514 -26358 27530 -26352
rect 27748 -26352 27838 -26324
rect 27748 -26358 27764 -26352
rect 27822 -26358 27838 -26352
rect 28056 -26358 28146 -26324
rect 28364 -26352 28454 -26324
rect 28364 -26358 28380 -26352
rect 28438 -26358 28454 -26352
rect 28672 -26352 28762 -26324
rect 28672 -26358 28688 -26352
rect 28746 -26358 28762 -26352
rect 28980 -26352 29070 -26324
rect 28980 -26358 28996 -26352
rect 29054 -26358 29070 -26352
rect 29288 -26358 29376 -26324
rect 24376 -26408 24536 -26358
rect 24696 -26402 24736 -26392
rect 24376 -27884 24388 -26408
rect 24422 -27884 24536 -26408
rect 24376 -27962 24536 -27884
rect 24636 -26408 24776 -26402
rect 24636 -27884 24696 -26408
rect 24730 -27884 24776 -26408
rect 24636 -28022 24776 -27884
rect 25004 -26408 25038 -26392
rect 25306 -26402 25346 -26392
rect 25004 -27900 25038 -27884
rect 25256 -26408 25396 -26402
rect 25256 -27884 25312 -26408
rect 25346 -27884 25396 -26408
rect 25256 -28022 25396 -27884
rect 25556 -26408 25716 -26358
rect 25926 -26402 25966 -26392
rect 25556 -27884 25620 -26408
rect 25654 -27884 25716 -26408
rect 25556 -27962 25716 -27884
rect 25876 -26408 26016 -26402
rect 25876 -27884 25928 -26408
rect 25962 -27884 26016 -26408
rect 25876 -28022 26016 -27884
rect 26236 -26408 26270 -26392
rect 26544 -26402 26578 -26392
rect 26236 -27900 26270 -27884
rect 26496 -26408 26636 -26402
rect 26496 -27884 26544 -26408
rect 26578 -27884 26636 -26408
rect 26496 -28022 26636 -27884
rect 26796 -26408 26956 -26358
rect 27160 -26402 27194 -26392
rect 26796 -27884 26852 -26408
rect 26886 -27884 26956 -26408
rect 26796 -27962 26956 -27884
rect 27096 -26408 27236 -26402
rect 27096 -27884 27160 -26408
rect 27194 -27884 27236 -26408
rect 27096 -28022 27236 -27884
rect 27468 -26408 27502 -26392
rect 27776 -26402 27810 -26392
rect 27468 -27900 27502 -27884
rect 27736 -26408 27876 -26402
rect 27736 -27884 27776 -26408
rect 27810 -27884 27876 -26408
rect 27736 -28022 27876 -27884
rect 28016 -26408 28176 -26358
rect 28392 -26402 28426 -26392
rect 28016 -27884 28084 -26408
rect 28118 -27884 28176 -26408
rect 28016 -27962 28176 -27884
rect 28336 -26408 28476 -26402
rect 28336 -27884 28392 -26408
rect 28426 -27884 28476 -26408
rect 28336 -28022 28476 -27884
rect 28700 -26408 28734 -26392
rect 29008 -26402 29042 -26392
rect 28700 -27900 28734 -27884
rect 28936 -26408 29076 -26402
rect 28936 -27884 29008 -26408
rect 29042 -27884 29076 -26408
rect 28936 -28022 29076 -27884
rect 29216 -26408 29376 -26358
rect 29216 -27884 29316 -26408
rect 29350 -27884 29376 -26408
rect 29216 -27962 29376 -27884
rect 29436 -26324 29816 -26322
rect 29436 -26358 29510 -26324
rect 29578 -26358 29668 -26324
rect 29736 -26358 29816 -26324
rect 29436 -26402 29816 -26358
rect 29436 -26408 29496 -26402
rect 29436 -27884 29448 -26408
rect 29482 -27884 29496 -26408
rect 29436 -28022 29496 -27884
rect 29596 -26408 29656 -26402
rect 29596 -27884 29606 -26408
rect 29640 -27884 29656 -26408
rect 29596 -28022 29656 -27884
rect 29756 -26408 29816 -26402
rect 29756 -27884 29764 -26408
rect 29798 -27884 29816 -26408
rect 29756 -28022 29816 -27884
rect 29896 -28002 29916 -26242
rect 29976 -26422 30896 -26242
rect 30956 -26422 30976 -24682
rect 31088 -24786 31122 -24770
rect 31336 -24786 31496 -24662
rect 31336 -26262 31396 -24786
rect 31430 -26262 31496 -24786
rect 31704 -24786 31738 -24770
rect 31936 -24786 32096 -24662
rect 32476 -24682 33256 -24662
rect 31936 -26262 32012 -24786
rect 32046 -26262 32096 -24786
rect 32320 -24786 32354 -24770
rect 31088 -26278 31122 -26262
rect 31396 -26278 31430 -26262
rect 31704 -26278 31738 -26262
rect 32012 -26278 32046 -26262
rect 32320 -26278 32354 -26262
rect 31134 -26346 31150 -26312
rect 31368 -26346 31384 -26312
rect 31442 -26346 31458 -26312
rect 31676 -26346 31692 -26312
rect 31750 -26346 31766 -26312
rect 31984 -26346 32000 -26312
rect 32058 -26346 32074 -26312
rect 32292 -26346 32308 -26312
rect 29976 -26442 30976 -26422
rect 32476 -26422 32496 -24682
rect 32556 -26422 33256 -24682
rect 32476 -26442 33256 -26422
rect 29976 -26462 33256 -26442
rect 29976 -26522 30996 -26462
rect 32456 -26522 33256 -26462
rect 29976 -28002 33256 -26522
rect 29896 -28022 33256 -28002
rect 20536 -28042 33256 -28022
rect 20536 -28102 23816 -28042
rect 29876 -28102 33256 -28042
rect 20536 -28182 33256 -28102
rect 20296 -28222 20496 -28202
rect 20296 -28242 23596 -28222
rect 20296 -28402 20516 -28242
rect 23376 -28402 23436 -28242
rect 20296 -28422 23436 -28402
rect 23396 -29402 23436 -28422
rect 23556 -29222 23596 -28242
rect 23636 -28242 30116 -28182
rect 33296 -28202 33316 -24322
rect 33476 -28202 33496 -19842
rect 33296 -28222 33496 -28202
rect 23636 -28322 23656 -28242
rect 23736 -28322 23776 -28242
rect 23856 -28322 23896 -28242
rect 23976 -28322 24016 -28242
rect 24096 -28322 24136 -28242
rect 24216 -28322 24256 -28242
rect 24336 -28322 24376 -28242
rect 24456 -28322 24496 -28242
rect 24576 -28322 24616 -28242
rect 24696 -28322 24736 -28242
rect 24816 -28322 24856 -28242
rect 24936 -28322 24976 -28242
rect 25056 -28322 25096 -28242
rect 25176 -28322 25216 -28242
rect 25296 -28322 25336 -28242
rect 25416 -28322 25456 -28242
rect 25536 -28322 25576 -28242
rect 25656 -28322 25696 -28242
rect 25776 -28322 25816 -28242
rect 25896 -28322 25936 -28242
rect 26016 -28322 26056 -28242
rect 26136 -28322 26176 -28242
rect 26256 -28322 26296 -28242
rect 26376 -28322 26416 -28242
rect 26496 -28322 26536 -28242
rect 26616 -28322 26656 -28242
rect 26736 -28322 26776 -28242
rect 26856 -28322 26896 -28242
rect 26976 -28322 27016 -28242
rect 27096 -28322 27136 -28242
rect 27216 -28322 27256 -28242
rect 27336 -28322 27376 -28242
rect 27456 -28322 27496 -28242
rect 27576 -28322 27616 -28242
rect 27696 -28322 27736 -28242
rect 27816 -28322 27856 -28242
rect 27936 -28322 27976 -28242
rect 28056 -28322 28096 -28242
rect 28176 -28322 28216 -28242
rect 28296 -28322 28336 -28242
rect 28416 -28322 28456 -28242
rect 28536 -28322 28576 -28242
rect 28656 -28322 28696 -28242
rect 28776 -28322 28816 -28242
rect 28896 -28322 28936 -28242
rect 29016 -28322 29056 -28242
rect 29136 -28322 29176 -28242
rect 29256 -28322 29296 -28242
rect 29376 -28322 29416 -28242
rect 29496 -28322 29536 -28242
rect 29616 -28322 29656 -28242
rect 29736 -28322 29776 -28242
rect 29856 -28322 29896 -28242
rect 29976 -28322 30016 -28242
rect 30096 -28322 30116 -28242
rect 23636 -28362 30116 -28322
rect 23636 -28442 23656 -28362
rect 23736 -28442 23776 -28362
rect 23856 -28442 23896 -28362
rect 23976 -28442 24016 -28362
rect 24096 -28442 24136 -28362
rect 24216 -28442 24256 -28362
rect 24336 -28442 24376 -28362
rect 24456 -28442 24496 -28362
rect 24576 -28442 24616 -28362
rect 24696 -28442 24736 -28362
rect 24816 -28442 24856 -28362
rect 24936 -28442 24976 -28362
rect 25056 -28442 25096 -28362
rect 25176 -28442 25216 -28362
rect 25296 -28442 25336 -28362
rect 25416 -28442 25456 -28362
rect 25536 -28442 25576 -28362
rect 25656 -28442 25696 -28362
rect 25776 -28442 25816 -28362
rect 25896 -28442 25936 -28362
rect 26016 -28442 26056 -28362
rect 26136 -28442 26176 -28362
rect 26256 -28442 26296 -28362
rect 26376 -28442 26416 -28362
rect 26496 -28442 26536 -28362
rect 26616 -28442 26656 -28362
rect 26736 -28442 26776 -28362
rect 26856 -28442 26896 -28362
rect 26976 -28442 27016 -28362
rect 27096 -28442 27136 -28362
rect 27216 -28442 27256 -28362
rect 27336 -28442 27376 -28362
rect 27456 -28442 27496 -28362
rect 27576 -28442 27616 -28362
rect 27696 -28442 27736 -28362
rect 27816 -28442 27856 -28362
rect 27936 -28442 27976 -28362
rect 28056 -28442 28096 -28362
rect 28176 -28442 28216 -28362
rect 28296 -28442 28336 -28362
rect 28416 -28442 28456 -28362
rect 28536 -28442 28576 -28362
rect 28656 -28442 28696 -28362
rect 28776 -28442 28816 -28362
rect 28896 -28442 28936 -28362
rect 29016 -28442 29056 -28362
rect 29136 -28442 29176 -28362
rect 29256 -28442 29296 -28362
rect 29376 -28442 29416 -28362
rect 29496 -28442 29536 -28362
rect 29616 -28442 29656 -28362
rect 29736 -28442 29776 -28362
rect 29856 -28442 29896 -28362
rect 29976 -28442 30016 -28362
rect 30096 -28442 30116 -28362
rect 23636 -28482 30116 -28442
rect 23636 -28562 23656 -28482
rect 23736 -28562 23776 -28482
rect 23856 -28562 23896 -28482
rect 23976 -28562 24016 -28482
rect 24096 -28562 24136 -28482
rect 24216 -28562 24256 -28482
rect 24336 -28562 24376 -28482
rect 24456 -28562 24496 -28482
rect 24576 -28562 24616 -28482
rect 24696 -28562 24736 -28482
rect 24816 -28562 24856 -28482
rect 24936 -28562 24976 -28482
rect 25056 -28562 25096 -28482
rect 25176 -28562 25216 -28482
rect 25296 -28562 25336 -28482
rect 25416 -28562 25456 -28482
rect 25536 -28562 25576 -28482
rect 25656 -28562 25696 -28482
rect 25776 -28562 25816 -28482
rect 25896 -28562 25936 -28482
rect 26016 -28562 26056 -28482
rect 26136 -28562 26176 -28482
rect 26256 -28562 26296 -28482
rect 26376 -28562 26416 -28482
rect 26496 -28562 26536 -28482
rect 26616 -28562 26656 -28482
rect 26736 -28562 26776 -28482
rect 26856 -28562 26896 -28482
rect 26976 -28562 27016 -28482
rect 27096 -28562 27136 -28482
rect 27216 -28562 27256 -28482
rect 27336 -28562 27376 -28482
rect 27456 -28562 27496 -28482
rect 27576 -28562 27616 -28482
rect 27696 -28562 27736 -28482
rect 27816 -28562 27856 -28482
rect 27936 -28562 27976 -28482
rect 28056 -28562 28096 -28482
rect 28176 -28562 28216 -28482
rect 28296 -28562 28336 -28482
rect 28416 -28562 28456 -28482
rect 28536 -28562 28576 -28482
rect 28656 -28562 28696 -28482
rect 28776 -28562 28816 -28482
rect 28896 -28562 28936 -28482
rect 29016 -28562 29056 -28482
rect 29136 -28562 29176 -28482
rect 29256 -28562 29296 -28482
rect 29376 -28562 29416 -28482
rect 29496 -28562 29536 -28482
rect 29616 -28562 29656 -28482
rect 29736 -28562 29776 -28482
rect 29856 -28562 29896 -28482
rect 29976 -28562 30016 -28482
rect 30096 -28562 30116 -28482
rect 23636 -28602 30116 -28562
rect 23636 -28682 23656 -28602
rect 23736 -28682 23776 -28602
rect 23856 -28682 23896 -28602
rect 23976 -28682 24016 -28602
rect 24096 -28682 24136 -28602
rect 24216 -28682 24256 -28602
rect 24336 -28682 24376 -28602
rect 24456 -28682 24496 -28602
rect 24576 -28682 24616 -28602
rect 24696 -28682 24736 -28602
rect 24816 -28682 24856 -28602
rect 24936 -28682 24976 -28602
rect 25056 -28682 25096 -28602
rect 25176 -28682 25216 -28602
rect 25296 -28682 25336 -28602
rect 25416 -28682 25456 -28602
rect 25536 -28682 25576 -28602
rect 25656 -28682 25696 -28602
rect 25776 -28682 25816 -28602
rect 25896 -28682 25936 -28602
rect 26016 -28682 26056 -28602
rect 26136 -28682 26176 -28602
rect 26256 -28682 26296 -28602
rect 26376 -28682 26416 -28602
rect 26496 -28682 26536 -28602
rect 26616 -28682 26656 -28602
rect 26736 -28682 26776 -28602
rect 26856 -28682 26896 -28602
rect 26976 -28682 27016 -28602
rect 27096 -28682 27136 -28602
rect 27216 -28682 27256 -28602
rect 27336 -28682 27376 -28602
rect 27456 -28682 27496 -28602
rect 27576 -28682 27616 -28602
rect 27696 -28682 27736 -28602
rect 27816 -28682 27856 -28602
rect 27936 -28682 27976 -28602
rect 28056 -28682 28096 -28602
rect 28176 -28682 28216 -28602
rect 28296 -28682 28336 -28602
rect 28416 -28682 28456 -28602
rect 28536 -28682 28576 -28602
rect 28656 -28682 28696 -28602
rect 28776 -28682 28816 -28602
rect 28896 -28682 28936 -28602
rect 29016 -28682 29056 -28602
rect 29136 -28682 29176 -28602
rect 29256 -28682 29296 -28602
rect 29376 -28682 29416 -28602
rect 29496 -28682 29536 -28602
rect 29616 -28682 29656 -28602
rect 29736 -28682 29776 -28602
rect 29856 -28682 29896 -28602
rect 29976 -28682 30016 -28602
rect 30096 -28682 30116 -28602
rect 23636 -28722 30116 -28682
rect 23636 -28802 23656 -28722
rect 23736 -28802 23776 -28722
rect 23856 -28802 23896 -28722
rect 23976 -28802 24016 -28722
rect 24096 -28802 24136 -28722
rect 24216 -28802 24256 -28722
rect 24336 -28802 24376 -28722
rect 24456 -28802 24496 -28722
rect 24576 -28802 24616 -28722
rect 24696 -28802 24736 -28722
rect 24816 -28802 24856 -28722
rect 24936 -28802 24976 -28722
rect 25056 -28802 25096 -28722
rect 25176 -28802 25216 -28722
rect 25296 -28802 25336 -28722
rect 25416 -28802 25456 -28722
rect 25536 -28802 25576 -28722
rect 25656 -28802 25696 -28722
rect 25776 -28802 25816 -28722
rect 25896 -28802 25936 -28722
rect 26016 -28802 26056 -28722
rect 26136 -28802 26176 -28722
rect 26256 -28802 26296 -28722
rect 26376 -28802 26416 -28722
rect 26496 -28802 26536 -28722
rect 26616 -28802 26656 -28722
rect 26736 -28802 26776 -28722
rect 26856 -28802 26896 -28722
rect 26976 -28802 27016 -28722
rect 27096 -28802 27136 -28722
rect 27216 -28802 27256 -28722
rect 27336 -28802 27376 -28722
rect 27456 -28802 27496 -28722
rect 27576 -28802 27616 -28722
rect 27696 -28802 27736 -28722
rect 27816 -28802 27856 -28722
rect 27936 -28802 27976 -28722
rect 28056 -28802 28096 -28722
rect 28176 -28802 28216 -28722
rect 28296 -28802 28336 -28722
rect 28416 -28802 28456 -28722
rect 28536 -28802 28576 -28722
rect 28656 -28802 28696 -28722
rect 28776 -28802 28816 -28722
rect 28896 -28802 28936 -28722
rect 29016 -28802 29056 -28722
rect 29136 -28802 29176 -28722
rect 29256 -28802 29296 -28722
rect 29376 -28802 29416 -28722
rect 29496 -28802 29536 -28722
rect 29616 -28802 29656 -28722
rect 29736 -28802 29776 -28722
rect 29856 -28802 29896 -28722
rect 29976 -28802 30016 -28722
rect 30096 -28802 30116 -28722
rect 23636 -28842 30116 -28802
rect 23636 -28922 23656 -28842
rect 23736 -28922 23776 -28842
rect 23856 -28922 23896 -28842
rect 23976 -28922 24016 -28842
rect 24096 -28922 24136 -28842
rect 24216 -28922 24256 -28842
rect 24336 -28922 24376 -28842
rect 24456 -28922 24496 -28842
rect 24576 -28922 24616 -28842
rect 24696 -28922 24736 -28842
rect 24816 -28922 24856 -28842
rect 24936 -28922 24976 -28842
rect 25056 -28922 25096 -28842
rect 25176 -28922 25216 -28842
rect 25296 -28922 25336 -28842
rect 25416 -28922 25456 -28842
rect 25536 -28922 25576 -28842
rect 25656 -28922 25696 -28842
rect 25776 -28922 25816 -28842
rect 25896 -28922 25936 -28842
rect 26016 -28922 26056 -28842
rect 26136 -28922 26176 -28842
rect 26256 -28922 26296 -28842
rect 26376 -28922 26416 -28842
rect 26496 -28922 26536 -28842
rect 26616 -28922 26656 -28842
rect 26736 -28922 26776 -28842
rect 26856 -28922 26896 -28842
rect 26976 -28922 27016 -28842
rect 27096 -28922 27136 -28842
rect 27216 -28922 27256 -28842
rect 27336 -28922 27376 -28842
rect 27456 -28922 27496 -28842
rect 27576 -28922 27616 -28842
rect 27696 -28922 27736 -28842
rect 27816 -28922 27856 -28842
rect 27936 -28922 27976 -28842
rect 28056 -28922 28096 -28842
rect 28176 -28922 28216 -28842
rect 28296 -28922 28336 -28842
rect 28416 -28922 28456 -28842
rect 28536 -28922 28576 -28842
rect 28656 -28922 28696 -28842
rect 28776 -28922 28816 -28842
rect 28896 -28922 28936 -28842
rect 29016 -28922 29056 -28842
rect 29136 -28922 29176 -28842
rect 29256 -28922 29296 -28842
rect 29376 -28922 29416 -28842
rect 29496 -28922 29536 -28842
rect 29616 -28922 29656 -28842
rect 29736 -28922 29776 -28842
rect 29856 -28922 29896 -28842
rect 29976 -28922 30016 -28842
rect 30096 -28922 30116 -28842
rect 23636 -28962 30116 -28922
rect 23636 -29042 23656 -28962
rect 23736 -29042 23776 -28962
rect 23856 -29042 23896 -28962
rect 23976 -29042 24016 -28962
rect 24096 -29042 24136 -28962
rect 24216 -29042 24256 -28962
rect 24336 -29042 24376 -28962
rect 24456 -29042 24496 -28962
rect 24576 -29042 24616 -28962
rect 24696 -29042 24736 -28962
rect 24816 -29042 24856 -28962
rect 24936 -29042 24976 -28962
rect 25056 -29042 25096 -28962
rect 25176 -29042 25216 -28962
rect 25296 -29042 25336 -28962
rect 25416 -29042 25456 -28962
rect 25536 -29042 25576 -28962
rect 25656 -29042 25696 -28962
rect 25776 -29042 25816 -28962
rect 25896 -29042 25936 -28962
rect 26016 -29042 26056 -28962
rect 26136 -29042 26176 -28962
rect 26256 -29042 26296 -28962
rect 26376 -29042 26416 -28962
rect 26496 -29042 26536 -28962
rect 26616 -29042 26656 -28962
rect 26736 -29042 26776 -28962
rect 26856 -29042 26896 -28962
rect 26976 -29042 27016 -28962
rect 27096 -29042 27136 -28962
rect 27216 -29042 27256 -28962
rect 27336 -29042 27376 -28962
rect 27456 -29042 27496 -28962
rect 27576 -29042 27616 -28962
rect 27696 -29042 27736 -28962
rect 27816 -29042 27856 -28962
rect 27936 -29042 27976 -28962
rect 28056 -29042 28096 -28962
rect 28176 -29042 28216 -28962
rect 28296 -29042 28336 -28962
rect 28416 -29042 28456 -28962
rect 28536 -29042 28576 -28962
rect 28656 -29042 28696 -28962
rect 28776 -29042 28816 -28962
rect 28896 -29042 28936 -28962
rect 29016 -29042 29056 -28962
rect 29136 -29042 29176 -28962
rect 29256 -29042 29296 -28962
rect 29376 -29042 29416 -28962
rect 29496 -29042 29536 -28962
rect 29616 -29042 29656 -28962
rect 29736 -29042 29776 -28962
rect 29856 -29042 29896 -28962
rect 29976 -29042 30016 -28962
rect 30096 -29042 30116 -28962
rect 23636 -29082 30116 -29042
rect 23636 -29162 23656 -29082
rect 23736 -29162 23776 -29082
rect 23856 -29162 23896 -29082
rect 23976 -29162 24016 -29082
rect 24096 -29162 24136 -29082
rect 24216 -29162 24256 -29082
rect 24336 -29162 24376 -29082
rect 24456 -29162 24496 -29082
rect 24576 -29162 24616 -29082
rect 24696 -29162 24736 -29082
rect 24816 -29162 24856 -29082
rect 24936 -29162 24976 -29082
rect 25056 -29162 25096 -29082
rect 25176 -29162 25216 -29082
rect 25296 -29162 25336 -29082
rect 25416 -29162 25456 -29082
rect 25536 -29162 25576 -29082
rect 25656 -29162 25696 -29082
rect 25776 -29162 25816 -29082
rect 25896 -29162 25936 -29082
rect 26016 -29162 26056 -29082
rect 26136 -29162 26176 -29082
rect 26256 -29162 26296 -29082
rect 26376 -29162 26416 -29082
rect 26496 -29162 26536 -29082
rect 26616 -29162 26656 -29082
rect 26736 -29162 26776 -29082
rect 26856 -29162 26896 -29082
rect 26976 -29162 27016 -29082
rect 27096 -29162 27136 -29082
rect 27216 -29162 27256 -29082
rect 27336 -29162 27376 -29082
rect 27456 -29162 27496 -29082
rect 27576 -29162 27616 -29082
rect 27696 -29162 27736 -29082
rect 27816 -29162 27856 -29082
rect 27936 -29162 27976 -29082
rect 28056 -29162 28096 -29082
rect 28176 -29162 28216 -29082
rect 28296 -29162 28336 -29082
rect 28416 -29162 28456 -29082
rect 28536 -29162 28576 -29082
rect 28656 -29162 28696 -29082
rect 28776 -29162 28816 -29082
rect 28896 -29162 28936 -29082
rect 29016 -29162 29056 -29082
rect 29136 -29162 29176 -29082
rect 29256 -29162 29296 -29082
rect 29376 -29162 29416 -29082
rect 29496 -29162 29536 -29082
rect 29616 -29162 29656 -29082
rect 29736 -29162 29776 -29082
rect 29856 -29162 29896 -29082
rect 29976 -29162 30016 -29082
rect 30096 -29162 30116 -29082
rect 23636 -29182 30116 -29162
rect 30156 -28242 33496 -28222
rect 30156 -29222 30196 -28242
rect 23556 -29242 30196 -29222
rect 23556 -29402 23596 -29242
rect 30156 -29402 30196 -29242
rect 30316 -28402 30356 -28242
rect 33276 -28402 33496 -28242
rect 30316 -28422 33496 -28402
rect 30316 -29402 30356 -28422
rect 23396 -29422 30356 -29402
<< viali >>
rect 23656 -19002 23736 -18922
rect 23776 -19002 23856 -18922
rect 23896 -19002 23976 -18922
rect 24016 -19002 24096 -18922
rect 24136 -19002 24216 -18922
rect 24256 -19002 24336 -18922
rect 24376 -19002 24456 -18922
rect 24496 -19002 24576 -18922
rect 24616 -19002 24696 -18922
rect 24736 -19002 24816 -18922
rect 24856 -19002 24936 -18922
rect 24976 -19002 25056 -18922
rect 25096 -19002 25176 -18922
rect 25216 -19002 25296 -18922
rect 25336 -19002 25416 -18922
rect 25456 -19002 25536 -18922
rect 25576 -19002 25656 -18922
rect 25696 -19002 25776 -18922
rect 25816 -19002 25896 -18922
rect 25936 -19002 26016 -18922
rect 26056 -19002 26136 -18922
rect 26176 -19002 26256 -18922
rect 26296 -19002 26376 -18922
rect 26416 -19002 26496 -18922
rect 26536 -19002 26616 -18922
rect 26656 -19002 26736 -18922
rect 26776 -19002 26856 -18922
rect 26896 -19002 26976 -18922
rect 27016 -19002 27096 -18922
rect 27136 -19002 27216 -18922
rect 27256 -19002 27336 -18922
rect 27376 -19002 27456 -18922
rect 27496 -19002 27576 -18922
rect 27616 -19002 27696 -18922
rect 27736 -19002 27816 -18922
rect 27856 -19002 27936 -18922
rect 27976 -19002 28056 -18922
rect 28096 -19002 28176 -18922
rect 28216 -19002 28296 -18922
rect 28336 -19002 28416 -18922
rect 28456 -19002 28536 -18922
rect 28576 -19002 28656 -18922
rect 28696 -19002 28776 -18922
rect 28816 -19002 28896 -18922
rect 28936 -19002 29016 -18922
rect 29056 -19002 29136 -18922
rect 29176 -19002 29256 -18922
rect 29296 -19002 29376 -18922
rect 29416 -19002 29496 -18922
rect 29536 -19002 29616 -18922
rect 29656 -19002 29736 -18922
rect 29776 -19002 29856 -18922
rect 29896 -19002 29976 -18922
rect 30016 -19002 30096 -18922
rect 23656 -19122 23736 -19042
rect 23776 -19122 23856 -19042
rect 23896 -19122 23976 -19042
rect 24016 -19122 24096 -19042
rect 24136 -19122 24216 -19042
rect 24256 -19122 24336 -19042
rect 24376 -19122 24456 -19042
rect 24496 -19122 24576 -19042
rect 24616 -19122 24696 -19042
rect 24736 -19122 24816 -19042
rect 24856 -19122 24936 -19042
rect 24976 -19122 25056 -19042
rect 25096 -19122 25176 -19042
rect 25216 -19122 25296 -19042
rect 25336 -19122 25416 -19042
rect 25456 -19122 25536 -19042
rect 25576 -19122 25656 -19042
rect 25696 -19122 25776 -19042
rect 25816 -19122 25896 -19042
rect 25936 -19122 26016 -19042
rect 26056 -19122 26136 -19042
rect 26176 -19122 26256 -19042
rect 26296 -19122 26376 -19042
rect 26416 -19122 26496 -19042
rect 26536 -19122 26616 -19042
rect 26656 -19122 26736 -19042
rect 26776 -19122 26856 -19042
rect 26896 -19122 26976 -19042
rect 27016 -19122 27096 -19042
rect 27136 -19122 27216 -19042
rect 27256 -19122 27336 -19042
rect 27376 -19122 27456 -19042
rect 27496 -19122 27576 -19042
rect 27616 -19122 27696 -19042
rect 27736 -19122 27816 -19042
rect 27856 -19122 27936 -19042
rect 27976 -19122 28056 -19042
rect 28096 -19122 28176 -19042
rect 28216 -19122 28296 -19042
rect 28336 -19122 28416 -19042
rect 28456 -19122 28536 -19042
rect 28576 -19122 28656 -19042
rect 28696 -19122 28776 -19042
rect 28816 -19122 28896 -19042
rect 28936 -19122 29016 -19042
rect 29056 -19122 29136 -19042
rect 29176 -19122 29256 -19042
rect 29296 -19122 29376 -19042
rect 29416 -19122 29496 -19042
rect 29536 -19122 29616 -19042
rect 29656 -19122 29736 -19042
rect 29776 -19122 29856 -19042
rect 29896 -19122 29976 -19042
rect 30016 -19122 30096 -19042
rect 23656 -19242 23736 -19162
rect 23776 -19242 23856 -19162
rect 23896 -19242 23976 -19162
rect 24016 -19242 24096 -19162
rect 24136 -19242 24216 -19162
rect 24256 -19242 24336 -19162
rect 24376 -19242 24456 -19162
rect 24496 -19242 24576 -19162
rect 24616 -19242 24696 -19162
rect 24736 -19242 24816 -19162
rect 24856 -19242 24936 -19162
rect 24976 -19242 25056 -19162
rect 25096 -19242 25176 -19162
rect 25216 -19242 25296 -19162
rect 25336 -19242 25416 -19162
rect 25456 -19242 25536 -19162
rect 25576 -19242 25656 -19162
rect 25696 -19242 25776 -19162
rect 25816 -19242 25896 -19162
rect 25936 -19242 26016 -19162
rect 26056 -19242 26136 -19162
rect 26176 -19242 26256 -19162
rect 26296 -19242 26376 -19162
rect 26416 -19242 26496 -19162
rect 26536 -19242 26616 -19162
rect 26656 -19242 26736 -19162
rect 26776 -19242 26856 -19162
rect 26896 -19242 26976 -19162
rect 27016 -19242 27096 -19162
rect 27136 -19242 27216 -19162
rect 27256 -19242 27336 -19162
rect 27376 -19242 27456 -19162
rect 27496 -19242 27576 -19162
rect 27616 -19242 27696 -19162
rect 27736 -19242 27816 -19162
rect 27856 -19242 27936 -19162
rect 27976 -19242 28056 -19162
rect 28096 -19242 28176 -19162
rect 28216 -19242 28296 -19162
rect 28336 -19242 28416 -19162
rect 28456 -19242 28536 -19162
rect 28576 -19242 28656 -19162
rect 28696 -19242 28776 -19162
rect 28816 -19242 28896 -19162
rect 28936 -19242 29016 -19162
rect 29056 -19242 29136 -19162
rect 29176 -19242 29256 -19162
rect 29296 -19242 29376 -19162
rect 29416 -19242 29496 -19162
rect 29536 -19242 29616 -19162
rect 29656 -19242 29736 -19162
rect 29776 -19242 29856 -19162
rect 29896 -19242 29976 -19162
rect 30016 -19242 30096 -19162
rect 23656 -19362 23736 -19282
rect 23776 -19362 23856 -19282
rect 23896 -19362 23976 -19282
rect 24016 -19362 24096 -19282
rect 24136 -19362 24216 -19282
rect 24256 -19362 24336 -19282
rect 24376 -19362 24456 -19282
rect 24496 -19362 24576 -19282
rect 24616 -19362 24696 -19282
rect 24736 -19362 24816 -19282
rect 24856 -19362 24936 -19282
rect 24976 -19362 25056 -19282
rect 25096 -19362 25176 -19282
rect 25216 -19362 25296 -19282
rect 25336 -19362 25416 -19282
rect 25456 -19362 25536 -19282
rect 25576 -19362 25656 -19282
rect 25696 -19362 25776 -19282
rect 25816 -19362 25896 -19282
rect 25936 -19362 26016 -19282
rect 26056 -19362 26136 -19282
rect 26176 -19362 26256 -19282
rect 26296 -19362 26376 -19282
rect 26416 -19362 26496 -19282
rect 26536 -19362 26616 -19282
rect 26656 -19362 26736 -19282
rect 26776 -19362 26856 -19282
rect 26896 -19362 26976 -19282
rect 27016 -19362 27096 -19282
rect 27136 -19362 27216 -19282
rect 27256 -19362 27336 -19282
rect 27376 -19362 27456 -19282
rect 27496 -19362 27576 -19282
rect 27616 -19362 27696 -19282
rect 27736 -19362 27816 -19282
rect 27856 -19362 27936 -19282
rect 27976 -19362 28056 -19282
rect 28096 -19362 28176 -19282
rect 28216 -19362 28296 -19282
rect 28336 -19362 28416 -19282
rect 28456 -19362 28536 -19282
rect 28576 -19362 28656 -19282
rect 28696 -19362 28776 -19282
rect 28816 -19362 28896 -19282
rect 28936 -19362 29016 -19282
rect 29056 -19362 29136 -19282
rect 29176 -19362 29256 -19282
rect 29296 -19362 29376 -19282
rect 29416 -19362 29496 -19282
rect 29536 -19362 29616 -19282
rect 29656 -19362 29736 -19282
rect 29776 -19362 29856 -19282
rect 29896 -19362 29976 -19282
rect 30016 -19362 30096 -19282
rect 23656 -19482 23736 -19402
rect 23776 -19482 23856 -19402
rect 23896 -19482 23976 -19402
rect 24016 -19482 24096 -19402
rect 24136 -19482 24216 -19402
rect 24256 -19482 24336 -19402
rect 24376 -19482 24456 -19402
rect 24496 -19482 24576 -19402
rect 24616 -19482 24696 -19402
rect 24736 -19482 24816 -19402
rect 24856 -19482 24936 -19402
rect 24976 -19482 25056 -19402
rect 25096 -19482 25176 -19402
rect 25216 -19482 25296 -19402
rect 25336 -19482 25416 -19402
rect 25456 -19482 25536 -19402
rect 25576 -19482 25656 -19402
rect 25696 -19482 25776 -19402
rect 25816 -19482 25896 -19402
rect 25936 -19482 26016 -19402
rect 26056 -19482 26136 -19402
rect 26176 -19482 26256 -19402
rect 26296 -19482 26376 -19402
rect 26416 -19482 26496 -19402
rect 26536 -19482 26616 -19402
rect 26656 -19482 26736 -19402
rect 26776 -19482 26856 -19402
rect 26896 -19482 26976 -19402
rect 27016 -19482 27096 -19402
rect 27136 -19482 27216 -19402
rect 27256 -19482 27336 -19402
rect 27376 -19482 27456 -19402
rect 27496 -19482 27576 -19402
rect 27616 -19482 27696 -19402
rect 27736 -19482 27816 -19402
rect 27856 -19482 27936 -19402
rect 27976 -19482 28056 -19402
rect 28096 -19482 28176 -19402
rect 28216 -19482 28296 -19402
rect 28336 -19482 28416 -19402
rect 28456 -19482 28536 -19402
rect 28576 -19482 28656 -19402
rect 28696 -19482 28776 -19402
rect 28816 -19482 28896 -19402
rect 28936 -19482 29016 -19402
rect 29056 -19482 29136 -19402
rect 29176 -19482 29256 -19402
rect 29296 -19482 29376 -19402
rect 29416 -19482 29496 -19402
rect 29536 -19482 29616 -19402
rect 29656 -19482 29736 -19402
rect 29776 -19482 29856 -19402
rect 29896 -19482 29976 -19402
rect 30016 -19482 30096 -19402
rect 23656 -19602 23736 -19522
rect 23776 -19602 23856 -19522
rect 23896 -19602 23976 -19522
rect 24016 -19602 24096 -19522
rect 24136 -19602 24216 -19522
rect 24256 -19602 24336 -19522
rect 24376 -19602 24456 -19522
rect 24496 -19602 24576 -19522
rect 24616 -19602 24696 -19522
rect 24736 -19602 24816 -19522
rect 24856 -19602 24936 -19522
rect 24976 -19602 25056 -19522
rect 25096 -19602 25176 -19522
rect 25216 -19602 25296 -19522
rect 25336 -19602 25416 -19522
rect 25456 -19602 25536 -19522
rect 25576 -19602 25656 -19522
rect 25696 -19602 25776 -19522
rect 25816 -19602 25896 -19522
rect 25936 -19602 26016 -19522
rect 26056 -19602 26136 -19522
rect 26176 -19602 26256 -19522
rect 26296 -19602 26376 -19522
rect 26416 -19602 26496 -19522
rect 26536 -19602 26616 -19522
rect 26656 -19602 26736 -19522
rect 26776 -19602 26856 -19522
rect 26896 -19602 26976 -19522
rect 27016 -19602 27096 -19522
rect 27136 -19602 27216 -19522
rect 27256 -19602 27336 -19522
rect 27376 -19602 27456 -19522
rect 27496 -19602 27576 -19522
rect 27616 -19602 27696 -19522
rect 27736 -19602 27816 -19522
rect 27856 -19602 27936 -19522
rect 27976 -19602 28056 -19522
rect 28096 -19602 28176 -19522
rect 28216 -19602 28296 -19522
rect 28336 -19602 28416 -19522
rect 28456 -19602 28536 -19522
rect 28576 -19602 28656 -19522
rect 28696 -19602 28776 -19522
rect 28816 -19602 28896 -19522
rect 28936 -19602 29016 -19522
rect 29056 -19602 29136 -19522
rect 29176 -19602 29256 -19522
rect 29296 -19602 29376 -19522
rect 29416 -19602 29496 -19522
rect 29536 -19602 29616 -19522
rect 29656 -19602 29736 -19522
rect 29776 -19602 29856 -19522
rect 29896 -19602 29976 -19522
rect 30016 -19602 30096 -19522
rect 20914 -22210 20948 -20234
rect 21222 -22210 21256 -20234
rect 21530 -22210 21564 -20234
rect 21838 -22210 21872 -20234
rect 22146 -22210 22180 -20234
rect 22454 -22210 22488 -20234
rect 22762 -22210 22796 -20234
rect 23070 -22210 23104 -20234
rect 23378 -22210 23412 -20234
rect 20976 -22303 21194 -22269
rect 21284 -22303 21502 -22269
rect 21592 -22303 21810 -22269
rect 21900 -22303 22118 -22269
rect 22208 -22303 22426 -22269
rect 22516 -22303 22734 -22269
rect 22824 -22303 23042 -22269
rect 23132 -22303 23350 -22269
rect 23914 -21730 23948 -19874
rect 24072 -21730 24106 -19874
rect 24230 -21730 24264 -19874
rect 24349 -21549 24383 -20065
rect 23976 -21823 24044 -21789
rect 24134 -21823 24202 -21789
rect 24657 -21549 24691 -20065
rect 24965 -21549 24999 -20065
rect 25273 -21549 25307 -20065
rect 25581 -21549 25615 -20065
rect 25889 -21549 25923 -20065
rect 26197 -21549 26231 -20065
rect 26505 -21549 26539 -20065
rect 26813 -21549 26847 -20065
rect 27121 -21549 27155 -20065
rect 27429 -21549 27463 -20065
rect 27737 -21549 27771 -20065
rect 28045 -21549 28079 -20065
rect 28353 -21549 28387 -20065
rect 28661 -21549 28695 -20065
rect 28969 -21549 29003 -20065
rect 29277 -21549 29311 -20065
rect 24411 -21828 24629 -21794
rect 24719 -21828 24937 -21794
rect 25027 -21828 25245 -21794
rect 25335 -21828 25553 -21794
rect 25643 -21828 25861 -21794
rect 25951 -21828 26169 -21794
rect 26259 -21828 26477 -21794
rect 26567 -21828 26785 -21794
rect 26875 -21828 27093 -21794
rect 27183 -21828 27401 -21794
rect 27491 -21828 27709 -21794
rect 27799 -21828 28017 -21794
rect 28107 -21828 28325 -21794
rect 28415 -21828 28633 -21794
rect 28723 -21828 28941 -21794
rect 29031 -21828 29249 -21794
rect 29454 -21730 29488 -19874
rect 29612 -21730 29646 -19874
rect 29770 -21730 29804 -19874
rect 29516 -21823 29584 -21789
rect 29674 -21823 29742 -21789
rect 30354 -22210 30388 -20234
rect 30662 -22210 30696 -20234
rect 30970 -22210 31004 -20234
rect 31278 -22210 31312 -20234
rect 31586 -22210 31620 -20234
rect 31894 -22210 31928 -20234
rect 32202 -22210 32236 -20234
rect 32510 -22210 32544 -20234
rect 32818 -22210 32852 -20234
rect 30416 -22303 30634 -22269
rect 30724 -22303 30942 -22269
rect 31032 -22303 31250 -22269
rect 31340 -22303 31558 -22269
rect 31648 -22303 31866 -22269
rect 31956 -22303 32174 -22269
rect 32264 -22303 32482 -22269
rect 32572 -22303 32790 -22269
rect 21874 -23910 21908 -22934
rect 22112 -23910 22146 -22934
rect 22350 -23910 22384 -22934
rect 21936 -24003 22084 -23969
rect 22174 -24003 22322 -23969
rect 21936 -24482 22016 -24402
rect 22076 -24482 22176 -24402
rect 22236 -24482 22316 -24402
rect 21428 -26242 21462 -24766
rect 21736 -26242 21770 -24766
rect 22044 -26242 22078 -24766
rect 22352 -26242 22386 -24766
rect 22660 -26242 22694 -24766
rect 21490 -26326 21708 -26292
rect 21798 -26326 22016 -26292
rect 22106 -26326 22324 -26292
rect 22414 -26326 22632 -26292
rect 26716 -23002 26796 -22922
rect 26856 -23002 26936 -22922
rect 26996 -23002 27076 -22922
rect 23368 -24082 23402 -23156
rect 23526 -24082 23560 -23156
rect 23684 -24082 23718 -23156
rect 23808 -24082 23842 -23156
rect 23966 -24082 24000 -23156
rect 24124 -24082 24158 -23156
rect 24248 -24082 24282 -23156
rect 24406 -24082 24440 -23156
rect 24564 -24082 24598 -23156
rect 23430 -24166 23498 -24132
rect 23588 -24166 23656 -24132
rect 23870 -24166 23938 -24132
rect 24028 -24166 24096 -24132
rect 24310 -24166 24378 -24132
rect 24468 -24166 24536 -24132
rect 24856 -23162 24936 -23082
rect 24856 -23282 24936 -23202
rect 24856 -23402 24936 -23322
rect 24856 -23522 24936 -23442
rect 24856 -23642 24936 -23562
rect 24856 -23762 24936 -23682
rect 24856 -23882 24936 -23802
rect 24856 -24002 24936 -23922
rect 24856 -24122 24936 -24042
rect 24856 -24242 24936 -24162
rect 25168 -24082 25202 -23156
rect 25326 -24082 25360 -23156
rect 25484 -24082 25518 -23156
rect 25608 -24082 25642 -23156
rect 25766 -24082 25800 -23156
rect 25924 -24082 25958 -23156
rect 26048 -24082 26082 -23156
rect 26206 -24082 26240 -23156
rect 26364 -24082 26398 -23156
rect 25230 -24166 25298 -24132
rect 25388 -24166 25456 -24132
rect 25670 -24166 25738 -24132
rect 25828 -24166 25896 -24132
rect 26110 -24166 26178 -24132
rect 26268 -24166 26336 -24132
rect 26716 -23122 26796 -23042
rect 26856 -23122 26936 -23042
rect 26996 -23122 27076 -23042
rect 26716 -23242 26796 -23162
rect 26856 -23242 26936 -23162
rect 26996 -23242 27076 -23162
rect 26716 -23362 26796 -23282
rect 26856 -23362 26936 -23282
rect 26996 -23362 27076 -23282
rect 26716 -23482 26796 -23402
rect 26856 -23482 26936 -23402
rect 26996 -23482 27076 -23402
rect 26716 -23602 26796 -23522
rect 26856 -23602 26936 -23522
rect 26996 -23602 27076 -23522
rect 26716 -23722 26796 -23642
rect 26856 -23722 26936 -23642
rect 26996 -23722 27076 -23642
rect 26716 -23842 26796 -23762
rect 26856 -23842 26936 -23762
rect 26996 -23842 27076 -23762
rect 26716 -23962 26796 -23882
rect 26856 -23962 26936 -23882
rect 26996 -23962 27076 -23882
rect 26716 -24082 26796 -24002
rect 26856 -24082 26936 -24002
rect 26996 -24082 27076 -24002
rect 24856 -24362 24936 -24282
rect 26716 -24202 26796 -24122
rect 26856 -24202 26936 -24122
rect 26996 -24202 27076 -24122
rect 27368 -24082 27402 -23156
rect 27526 -24082 27560 -23156
rect 27684 -24082 27718 -23156
rect 27808 -24082 27842 -23156
rect 27966 -24082 28000 -23156
rect 28124 -24082 28158 -23156
rect 28248 -24082 28282 -23156
rect 28406 -24082 28440 -23156
rect 28564 -24082 28598 -23156
rect 27430 -24166 27498 -24132
rect 27588 -24166 27656 -24132
rect 27870 -24166 27938 -24132
rect 28028 -24166 28096 -24132
rect 28310 -24166 28378 -24132
rect 28468 -24166 28536 -24132
rect 28856 -23162 28936 -23082
rect 28856 -23282 28936 -23202
rect 28856 -23402 28936 -23322
rect 28856 -23522 28936 -23442
rect 28856 -23642 28936 -23562
rect 28856 -23762 28936 -23682
rect 28856 -23882 28936 -23802
rect 28856 -24002 28936 -23922
rect 28856 -24122 28936 -24042
rect 26716 -24322 26796 -24242
rect 26856 -24322 26936 -24242
rect 26996 -24322 27076 -24242
rect 28856 -24242 28936 -24162
rect 29168 -24082 29202 -23156
rect 29326 -24082 29360 -23156
rect 29484 -24082 29518 -23156
rect 29608 -24082 29642 -23156
rect 29766 -24082 29800 -23156
rect 29924 -24082 29958 -23156
rect 30048 -24082 30082 -23156
rect 30206 -24082 30240 -23156
rect 30364 -24082 30398 -23156
rect 29230 -24166 29298 -24132
rect 29388 -24166 29456 -24132
rect 29670 -24166 29738 -24132
rect 29828 -24166 29896 -24132
rect 30110 -24166 30178 -24132
rect 30268 -24166 30336 -24132
rect 28856 -24362 28936 -24282
rect 23236 -24442 23316 -24362
rect 23356 -24442 23436 -24362
rect 23476 -24442 23556 -24362
rect 23596 -24442 23676 -24362
rect 23716 -24442 23796 -24362
rect 23836 -24442 23916 -24362
rect 23956 -24442 24036 -24362
rect 24076 -24442 24156 -24362
rect 24196 -24442 24276 -24362
rect 24316 -24442 24396 -24362
rect 24436 -24442 24516 -24362
rect 24556 -24442 24636 -24362
rect 24676 -24442 24756 -24362
rect 24856 -24482 24936 -24402
rect 25036 -24442 25116 -24362
rect 25156 -24442 25236 -24362
rect 25276 -24442 25356 -24362
rect 25396 -24442 25476 -24362
rect 25516 -24442 25596 -24362
rect 25636 -24442 25716 -24362
rect 25756 -24442 25836 -24362
rect 25876 -24442 25956 -24362
rect 25996 -24442 26076 -24362
rect 26116 -24442 26196 -24362
rect 26236 -24442 26316 -24362
rect 26356 -24442 26436 -24362
rect 26476 -24442 26556 -24362
rect 26596 -24442 26676 -24362
rect 26716 -24442 26796 -24362
rect 26856 -24442 26936 -24362
rect 26996 -24442 27076 -24362
rect 27116 -24442 27196 -24362
rect 27236 -24442 27316 -24362
rect 27356 -24442 27436 -24362
rect 27476 -24442 27556 -24362
rect 27596 -24442 27676 -24362
rect 27716 -24442 27796 -24362
rect 27836 -24442 27916 -24362
rect 27956 -24442 28036 -24362
rect 28076 -24442 28156 -24362
rect 28196 -24442 28276 -24362
rect 28316 -24442 28396 -24362
rect 28436 -24442 28516 -24362
rect 28556 -24442 28636 -24362
rect 28676 -24442 28756 -24362
rect 28856 -24482 28936 -24402
rect 29036 -24442 29116 -24362
rect 29156 -24442 29236 -24362
rect 29276 -24442 29356 -24362
rect 29396 -24442 29476 -24362
rect 29516 -24442 29596 -24362
rect 29636 -24442 29716 -24362
rect 29756 -24442 29836 -24362
rect 29876 -24442 29956 -24362
rect 29996 -24442 30076 -24362
rect 30116 -24442 30196 -24362
rect 30236 -24442 30316 -24362
rect 30356 -24442 30436 -24362
rect 30476 -24442 30556 -24362
rect 23236 -24582 23316 -24502
rect 23356 -24582 23436 -24502
rect 23476 -24582 23556 -24502
rect 23596 -24582 23676 -24502
rect 23716 -24582 23796 -24502
rect 23836 -24582 23916 -24502
rect 23956 -24582 24036 -24502
rect 24076 -24582 24156 -24502
rect 24196 -24582 24276 -24502
rect 24316 -24582 24396 -24502
rect 24436 -24582 24516 -24502
rect 24556 -24582 24636 -24502
rect 24676 -24582 24756 -24502
rect 24856 -24602 24936 -24522
rect 25036 -24582 25116 -24502
rect 25156 -24582 25236 -24502
rect 25276 -24582 25356 -24502
rect 25396 -24582 25476 -24502
rect 25516 -24582 25596 -24502
rect 25636 -24582 25716 -24502
rect 25756 -24582 25836 -24502
rect 25876 -24582 25956 -24502
rect 25996 -24582 26076 -24502
rect 26116 -24582 26196 -24502
rect 26236 -24582 26316 -24502
rect 26356 -24582 26436 -24502
rect 26476 -24582 26556 -24502
rect 26596 -24582 26676 -24502
rect 26716 -24562 26796 -24482
rect 26856 -24562 26936 -24482
rect 26996 -24562 27076 -24482
rect 27116 -24582 27196 -24502
rect 27236 -24582 27316 -24502
rect 27356 -24582 27436 -24502
rect 27476 -24582 27556 -24502
rect 27596 -24582 27676 -24502
rect 27716 -24582 27796 -24502
rect 27836 -24582 27916 -24502
rect 27956 -24582 28036 -24502
rect 28076 -24582 28156 -24502
rect 28196 -24582 28276 -24502
rect 28316 -24582 28396 -24502
rect 28436 -24582 28516 -24502
rect 28556 -24582 28636 -24502
rect 28676 -24582 28756 -24502
rect 28856 -24602 28936 -24522
rect 29036 -24582 29116 -24502
rect 29156 -24582 29236 -24502
rect 29276 -24582 29356 -24502
rect 29396 -24582 29476 -24502
rect 29516 -24582 29596 -24502
rect 29636 -24582 29716 -24502
rect 29756 -24582 29836 -24502
rect 29876 -24582 29956 -24502
rect 29996 -24582 30076 -24502
rect 30116 -24582 30196 -24502
rect 30236 -24582 30316 -24502
rect 30356 -24582 30436 -24502
rect 30476 -24582 30556 -24502
rect 24856 -24722 24936 -24642
rect 26716 -24682 26796 -24602
rect 26856 -24682 26936 -24602
rect 26996 -24682 27076 -24602
rect 23430 -24808 23498 -24774
rect 23588 -24808 23656 -24774
rect 23870 -24808 23938 -24774
rect 24028 -24808 24096 -24774
rect 24310 -24808 24378 -24774
rect 24468 -24808 24536 -24774
rect 23368 -25784 23402 -24858
rect 23526 -25784 23560 -24858
rect 23684 -25784 23718 -24858
rect 23808 -25784 23842 -24858
rect 23966 -25784 24000 -24858
rect 24124 -25784 24158 -24858
rect 24248 -25784 24282 -24858
rect 24406 -25784 24440 -24858
rect 24564 -25784 24598 -24858
rect 24856 -24842 24936 -24762
rect 24856 -24962 24936 -24882
rect 24856 -25082 24936 -25002
rect 24856 -25202 24936 -25122
rect 24856 -25322 24936 -25242
rect 24856 -25442 24936 -25362
rect 24856 -25562 24936 -25482
rect 24856 -25682 24936 -25602
rect 24856 -25802 24936 -25722
rect 25230 -24808 25298 -24774
rect 25388 -24808 25456 -24774
rect 25670 -24808 25738 -24774
rect 25828 -24808 25896 -24774
rect 26110 -24808 26178 -24774
rect 26268 -24808 26336 -24774
rect 25168 -25784 25202 -24858
rect 25326 -25784 25360 -24858
rect 25484 -25784 25518 -24858
rect 25608 -25784 25642 -24858
rect 25766 -25784 25800 -24858
rect 25924 -25784 25958 -24858
rect 26048 -25784 26082 -24858
rect 26206 -25784 26240 -24858
rect 26364 -25784 26398 -24858
rect 26716 -24802 26796 -24722
rect 26856 -24802 26936 -24722
rect 26996 -24802 27076 -24722
rect 28856 -24722 28936 -24642
rect 26716 -24922 26796 -24842
rect 26856 -24922 26936 -24842
rect 26996 -24922 27076 -24842
rect 26716 -25042 26796 -24962
rect 26856 -25042 26936 -24962
rect 26996 -25042 27076 -24962
rect 26716 -25162 26796 -25082
rect 26856 -25162 26936 -25082
rect 26996 -25162 27076 -25082
rect 26716 -25282 26796 -25202
rect 26856 -25282 26936 -25202
rect 26996 -25282 27076 -25202
rect 26716 -25402 26796 -25322
rect 26856 -25402 26936 -25322
rect 26996 -25402 27076 -25322
rect 26716 -25522 26796 -25442
rect 26856 -25522 26936 -25442
rect 26996 -25522 27076 -25442
rect 26716 -25642 26796 -25562
rect 26856 -25642 26936 -25562
rect 26996 -25642 27076 -25562
rect 26716 -25762 26796 -25682
rect 26856 -25762 26936 -25682
rect 26996 -25762 27076 -25682
rect 26716 -25882 26796 -25802
rect 26856 -25882 26936 -25802
rect 26996 -25882 27076 -25802
rect 27430 -24808 27498 -24774
rect 27588 -24808 27656 -24774
rect 27870 -24808 27938 -24774
rect 28028 -24808 28096 -24774
rect 28310 -24808 28378 -24774
rect 28468 -24808 28536 -24774
rect 27368 -25784 27402 -24858
rect 27526 -25784 27560 -24858
rect 27684 -25784 27718 -24858
rect 27808 -25784 27842 -24858
rect 27966 -25784 28000 -24858
rect 28124 -25784 28158 -24858
rect 28248 -25784 28282 -24858
rect 28406 -25784 28440 -24858
rect 28564 -25784 28598 -24858
rect 28856 -24842 28936 -24762
rect 28856 -24962 28936 -24882
rect 28856 -25082 28936 -25002
rect 28856 -25202 28936 -25122
rect 28856 -25322 28936 -25242
rect 28856 -25442 28936 -25362
rect 28856 -25562 28936 -25482
rect 28856 -25682 28936 -25602
rect 28856 -25802 28936 -25722
rect 29230 -24808 29298 -24774
rect 29388 -24808 29456 -24774
rect 29670 -24808 29738 -24774
rect 29828 -24808 29896 -24774
rect 30110 -24808 30178 -24774
rect 30268 -24808 30336 -24774
rect 29168 -25784 29202 -24858
rect 29326 -25784 29360 -24858
rect 29484 -25784 29518 -24858
rect 29608 -25784 29642 -24858
rect 29766 -25784 29800 -24858
rect 29924 -25784 29958 -24858
rect 30048 -25784 30082 -24858
rect 30206 -25784 30240 -24858
rect 30364 -25784 30398 -24858
rect 26716 -26002 26796 -25922
rect 26856 -26002 26936 -25922
rect 26996 -26002 27076 -25922
rect 31454 -23890 31488 -22914
rect 31692 -23890 31726 -22914
rect 31930 -23890 31964 -22914
rect 31516 -23983 31664 -23949
rect 31754 -23983 31902 -23949
rect 31516 -24482 31596 -24402
rect 31636 -24482 31776 -24402
rect 31816 -24482 31896 -24402
rect 24010 -26358 24078 -26324
rect 24168 -26358 24236 -26324
rect 23948 -27884 23982 -26408
rect 24106 -27884 24140 -26408
rect 24264 -27884 24298 -26408
rect 24450 -26358 24668 -26324
rect 24758 -26358 24976 -26324
rect 25066 -26358 25284 -26324
rect 25374 -26358 25592 -26324
rect 25682 -26358 25900 -26324
rect 25990 -26358 26208 -26324
rect 26298 -26358 26516 -26324
rect 26606 -26358 26824 -26324
rect 26914 -26358 27132 -26324
rect 27222 -26358 27440 -26324
rect 27530 -26358 27748 -26324
rect 27838 -26358 28056 -26324
rect 28146 -26358 28364 -26324
rect 28454 -26358 28672 -26324
rect 28762 -26358 28980 -26324
rect 29070 -26358 29288 -26324
rect 24388 -27884 24422 -26408
rect 24696 -27884 24730 -26408
rect 25004 -27884 25038 -26408
rect 25312 -27884 25346 -26408
rect 25620 -27884 25654 -26408
rect 25928 -27884 25962 -26408
rect 26236 -27884 26270 -26408
rect 26544 -27884 26578 -26408
rect 26852 -27884 26886 -26408
rect 27160 -27884 27194 -26408
rect 27468 -27884 27502 -26408
rect 27776 -27884 27810 -26408
rect 28084 -27884 28118 -26408
rect 28392 -27884 28426 -26408
rect 28700 -27884 28734 -26408
rect 29008 -27884 29042 -26408
rect 29316 -27884 29350 -26408
rect 29510 -26358 29578 -26324
rect 29668 -26358 29736 -26324
rect 29448 -27884 29482 -26408
rect 29606 -27884 29640 -26408
rect 29764 -27884 29798 -26408
rect 31088 -26262 31122 -24786
rect 31396 -26262 31430 -24786
rect 31704 -26262 31738 -24786
rect 32012 -26262 32046 -24786
rect 32320 -26262 32354 -24786
rect 31150 -26346 31368 -26312
rect 31458 -26346 31676 -26312
rect 31766 -26346 31984 -26312
rect 32074 -26346 32292 -26312
rect 23656 -28322 23736 -28242
rect 23776 -28322 23856 -28242
rect 23896 -28322 23976 -28242
rect 24016 -28322 24096 -28242
rect 24136 -28322 24216 -28242
rect 24256 -28322 24336 -28242
rect 24376 -28322 24456 -28242
rect 24496 -28322 24576 -28242
rect 24616 -28322 24696 -28242
rect 24736 -28322 24816 -28242
rect 24856 -28322 24936 -28242
rect 24976 -28322 25056 -28242
rect 25096 -28322 25176 -28242
rect 25216 -28322 25296 -28242
rect 25336 -28322 25416 -28242
rect 25456 -28322 25536 -28242
rect 25576 -28322 25656 -28242
rect 25696 -28322 25776 -28242
rect 25816 -28322 25896 -28242
rect 25936 -28322 26016 -28242
rect 26056 -28322 26136 -28242
rect 26176 -28322 26256 -28242
rect 26296 -28322 26376 -28242
rect 26416 -28322 26496 -28242
rect 26536 -28322 26616 -28242
rect 26656 -28322 26736 -28242
rect 26776 -28322 26856 -28242
rect 26896 -28322 26976 -28242
rect 27016 -28322 27096 -28242
rect 27136 -28322 27216 -28242
rect 27256 -28322 27336 -28242
rect 27376 -28322 27456 -28242
rect 27496 -28322 27576 -28242
rect 27616 -28322 27696 -28242
rect 27736 -28322 27816 -28242
rect 27856 -28322 27936 -28242
rect 27976 -28322 28056 -28242
rect 28096 -28322 28176 -28242
rect 28216 -28322 28296 -28242
rect 28336 -28322 28416 -28242
rect 28456 -28322 28536 -28242
rect 28576 -28322 28656 -28242
rect 28696 -28322 28776 -28242
rect 28816 -28322 28896 -28242
rect 28936 -28322 29016 -28242
rect 29056 -28322 29136 -28242
rect 29176 -28322 29256 -28242
rect 29296 -28322 29376 -28242
rect 29416 -28322 29496 -28242
rect 29536 -28322 29616 -28242
rect 29656 -28322 29736 -28242
rect 29776 -28322 29856 -28242
rect 29896 -28322 29976 -28242
rect 30016 -28322 30096 -28242
rect 23656 -28442 23736 -28362
rect 23776 -28442 23856 -28362
rect 23896 -28442 23976 -28362
rect 24016 -28442 24096 -28362
rect 24136 -28442 24216 -28362
rect 24256 -28442 24336 -28362
rect 24376 -28442 24456 -28362
rect 24496 -28442 24576 -28362
rect 24616 -28442 24696 -28362
rect 24736 -28442 24816 -28362
rect 24856 -28442 24936 -28362
rect 24976 -28442 25056 -28362
rect 25096 -28442 25176 -28362
rect 25216 -28442 25296 -28362
rect 25336 -28442 25416 -28362
rect 25456 -28442 25536 -28362
rect 25576 -28442 25656 -28362
rect 25696 -28442 25776 -28362
rect 25816 -28442 25896 -28362
rect 25936 -28442 26016 -28362
rect 26056 -28442 26136 -28362
rect 26176 -28442 26256 -28362
rect 26296 -28442 26376 -28362
rect 26416 -28442 26496 -28362
rect 26536 -28442 26616 -28362
rect 26656 -28442 26736 -28362
rect 26776 -28442 26856 -28362
rect 26896 -28442 26976 -28362
rect 27016 -28442 27096 -28362
rect 27136 -28442 27216 -28362
rect 27256 -28442 27336 -28362
rect 27376 -28442 27456 -28362
rect 27496 -28442 27576 -28362
rect 27616 -28442 27696 -28362
rect 27736 -28442 27816 -28362
rect 27856 -28442 27936 -28362
rect 27976 -28442 28056 -28362
rect 28096 -28442 28176 -28362
rect 28216 -28442 28296 -28362
rect 28336 -28442 28416 -28362
rect 28456 -28442 28536 -28362
rect 28576 -28442 28656 -28362
rect 28696 -28442 28776 -28362
rect 28816 -28442 28896 -28362
rect 28936 -28442 29016 -28362
rect 29056 -28442 29136 -28362
rect 29176 -28442 29256 -28362
rect 29296 -28442 29376 -28362
rect 29416 -28442 29496 -28362
rect 29536 -28442 29616 -28362
rect 29656 -28442 29736 -28362
rect 29776 -28442 29856 -28362
rect 29896 -28442 29976 -28362
rect 30016 -28442 30096 -28362
rect 23656 -28562 23736 -28482
rect 23776 -28562 23856 -28482
rect 23896 -28562 23976 -28482
rect 24016 -28562 24096 -28482
rect 24136 -28562 24216 -28482
rect 24256 -28562 24336 -28482
rect 24376 -28562 24456 -28482
rect 24496 -28562 24576 -28482
rect 24616 -28562 24696 -28482
rect 24736 -28562 24816 -28482
rect 24856 -28562 24936 -28482
rect 24976 -28562 25056 -28482
rect 25096 -28562 25176 -28482
rect 25216 -28562 25296 -28482
rect 25336 -28562 25416 -28482
rect 25456 -28562 25536 -28482
rect 25576 -28562 25656 -28482
rect 25696 -28562 25776 -28482
rect 25816 -28562 25896 -28482
rect 25936 -28562 26016 -28482
rect 26056 -28562 26136 -28482
rect 26176 -28562 26256 -28482
rect 26296 -28562 26376 -28482
rect 26416 -28562 26496 -28482
rect 26536 -28562 26616 -28482
rect 26656 -28562 26736 -28482
rect 26776 -28562 26856 -28482
rect 26896 -28562 26976 -28482
rect 27016 -28562 27096 -28482
rect 27136 -28562 27216 -28482
rect 27256 -28562 27336 -28482
rect 27376 -28562 27456 -28482
rect 27496 -28562 27576 -28482
rect 27616 -28562 27696 -28482
rect 27736 -28562 27816 -28482
rect 27856 -28562 27936 -28482
rect 27976 -28562 28056 -28482
rect 28096 -28562 28176 -28482
rect 28216 -28562 28296 -28482
rect 28336 -28562 28416 -28482
rect 28456 -28562 28536 -28482
rect 28576 -28562 28656 -28482
rect 28696 -28562 28776 -28482
rect 28816 -28562 28896 -28482
rect 28936 -28562 29016 -28482
rect 29056 -28562 29136 -28482
rect 29176 -28562 29256 -28482
rect 29296 -28562 29376 -28482
rect 29416 -28562 29496 -28482
rect 29536 -28562 29616 -28482
rect 29656 -28562 29736 -28482
rect 29776 -28562 29856 -28482
rect 29896 -28562 29976 -28482
rect 30016 -28562 30096 -28482
rect 23656 -28682 23736 -28602
rect 23776 -28682 23856 -28602
rect 23896 -28682 23976 -28602
rect 24016 -28682 24096 -28602
rect 24136 -28682 24216 -28602
rect 24256 -28682 24336 -28602
rect 24376 -28682 24456 -28602
rect 24496 -28682 24576 -28602
rect 24616 -28682 24696 -28602
rect 24736 -28682 24816 -28602
rect 24856 -28682 24936 -28602
rect 24976 -28682 25056 -28602
rect 25096 -28682 25176 -28602
rect 25216 -28682 25296 -28602
rect 25336 -28682 25416 -28602
rect 25456 -28682 25536 -28602
rect 25576 -28682 25656 -28602
rect 25696 -28682 25776 -28602
rect 25816 -28682 25896 -28602
rect 25936 -28682 26016 -28602
rect 26056 -28682 26136 -28602
rect 26176 -28682 26256 -28602
rect 26296 -28682 26376 -28602
rect 26416 -28682 26496 -28602
rect 26536 -28682 26616 -28602
rect 26656 -28682 26736 -28602
rect 26776 -28682 26856 -28602
rect 26896 -28682 26976 -28602
rect 27016 -28682 27096 -28602
rect 27136 -28682 27216 -28602
rect 27256 -28682 27336 -28602
rect 27376 -28682 27456 -28602
rect 27496 -28682 27576 -28602
rect 27616 -28682 27696 -28602
rect 27736 -28682 27816 -28602
rect 27856 -28682 27936 -28602
rect 27976 -28682 28056 -28602
rect 28096 -28682 28176 -28602
rect 28216 -28682 28296 -28602
rect 28336 -28682 28416 -28602
rect 28456 -28682 28536 -28602
rect 28576 -28682 28656 -28602
rect 28696 -28682 28776 -28602
rect 28816 -28682 28896 -28602
rect 28936 -28682 29016 -28602
rect 29056 -28682 29136 -28602
rect 29176 -28682 29256 -28602
rect 29296 -28682 29376 -28602
rect 29416 -28682 29496 -28602
rect 29536 -28682 29616 -28602
rect 29656 -28682 29736 -28602
rect 29776 -28682 29856 -28602
rect 29896 -28682 29976 -28602
rect 30016 -28682 30096 -28602
rect 23656 -28802 23736 -28722
rect 23776 -28802 23856 -28722
rect 23896 -28802 23976 -28722
rect 24016 -28802 24096 -28722
rect 24136 -28802 24216 -28722
rect 24256 -28802 24336 -28722
rect 24376 -28802 24456 -28722
rect 24496 -28802 24576 -28722
rect 24616 -28802 24696 -28722
rect 24736 -28802 24816 -28722
rect 24856 -28802 24936 -28722
rect 24976 -28802 25056 -28722
rect 25096 -28802 25176 -28722
rect 25216 -28802 25296 -28722
rect 25336 -28802 25416 -28722
rect 25456 -28802 25536 -28722
rect 25576 -28802 25656 -28722
rect 25696 -28802 25776 -28722
rect 25816 -28802 25896 -28722
rect 25936 -28802 26016 -28722
rect 26056 -28802 26136 -28722
rect 26176 -28802 26256 -28722
rect 26296 -28802 26376 -28722
rect 26416 -28802 26496 -28722
rect 26536 -28802 26616 -28722
rect 26656 -28802 26736 -28722
rect 26776 -28802 26856 -28722
rect 26896 -28802 26976 -28722
rect 27016 -28802 27096 -28722
rect 27136 -28802 27216 -28722
rect 27256 -28802 27336 -28722
rect 27376 -28802 27456 -28722
rect 27496 -28802 27576 -28722
rect 27616 -28802 27696 -28722
rect 27736 -28802 27816 -28722
rect 27856 -28802 27936 -28722
rect 27976 -28802 28056 -28722
rect 28096 -28802 28176 -28722
rect 28216 -28802 28296 -28722
rect 28336 -28802 28416 -28722
rect 28456 -28802 28536 -28722
rect 28576 -28802 28656 -28722
rect 28696 -28802 28776 -28722
rect 28816 -28802 28896 -28722
rect 28936 -28802 29016 -28722
rect 29056 -28802 29136 -28722
rect 29176 -28802 29256 -28722
rect 29296 -28802 29376 -28722
rect 29416 -28802 29496 -28722
rect 29536 -28802 29616 -28722
rect 29656 -28802 29736 -28722
rect 29776 -28802 29856 -28722
rect 29896 -28802 29976 -28722
rect 30016 -28802 30096 -28722
rect 23656 -28922 23736 -28842
rect 23776 -28922 23856 -28842
rect 23896 -28922 23976 -28842
rect 24016 -28922 24096 -28842
rect 24136 -28922 24216 -28842
rect 24256 -28922 24336 -28842
rect 24376 -28922 24456 -28842
rect 24496 -28922 24576 -28842
rect 24616 -28922 24696 -28842
rect 24736 -28922 24816 -28842
rect 24856 -28922 24936 -28842
rect 24976 -28922 25056 -28842
rect 25096 -28922 25176 -28842
rect 25216 -28922 25296 -28842
rect 25336 -28922 25416 -28842
rect 25456 -28922 25536 -28842
rect 25576 -28922 25656 -28842
rect 25696 -28922 25776 -28842
rect 25816 -28922 25896 -28842
rect 25936 -28922 26016 -28842
rect 26056 -28922 26136 -28842
rect 26176 -28922 26256 -28842
rect 26296 -28922 26376 -28842
rect 26416 -28922 26496 -28842
rect 26536 -28922 26616 -28842
rect 26656 -28922 26736 -28842
rect 26776 -28922 26856 -28842
rect 26896 -28922 26976 -28842
rect 27016 -28922 27096 -28842
rect 27136 -28922 27216 -28842
rect 27256 -28922 27336 -28842
rect 27376 -28922 27456 -28842
rect 27496 -28922 27576 -28842
rect 27616 -28922 27696 -28842
rect 27736 -28922 27816 -28842
rect 27856 -28922 27936 -28842
rect 27976 -28922 28056 -28842
rect 28096 -28922 28176 -28842
rect 28216 -28922 28296 -28842
rect 28336 -28922 28416 -28842
rect 28456 -28922 28536 -28842
rect 28576 -28922 28656 -28842
rect 28696 -28922 28776 -28842
rect 28816 -28922 28896 -28842
rect 28936 -28922 29016 -28842
rect 29056 -28922 29136 -28842
rect 29176 -28922 29256 -28842
rect 29296 -28922 29376 -28842
rect 29416 -28922 29496 -28842
rect 29536 -28922 29616 -28842
rect 29656 -28922 29736 -28842
rect 29776 -28922 29856 -28842
rect 29896 -28922 29976 -28842
rect 30016 -28922 30096 -28842
rect 23656 -29042 23736 -28962
rect 23776 -29042 23856 -28962
rect 23896 -29042 23976 -28962
rect 24016 -29042 24096 -28962
rect 24136 -29042 24216 -28962
rect 24256 -29042 24336 -28962
rect 24376 -29042 24456 -28962
rect 24496 -29042 24576 -28962
rect 24616 -29042 24696 -28962
rect 24736 -29042 24816 -28962
rect 24856 -29042 24936 -28962
rect 24976 -29042 25056 -28962
rect 25096 -29042 25176 -28962
rect 25216 -29042 25296 -28962
rect 25336 -29042 25416 -28962
rect 25456 -29042 25536 -28962
rect 25576 -29042 25656 -28962
rect 25696 -29042 25776 -28962
rect 25816 -29042 25896 -28962
rect 25936 -29042 26016 -28962
rect 26056 -29042 26136 -28962
rect 26176 -29042 26256 -28962
rect 26296 -29042 26376 -28962
rect 26416 -29042 26496 -28962
rect 26536 -29042 26616 -28962
rect 26656 -29042 26736 -28962
rect 26776 -29042 26856 -28962
rect 26896 -29042 26976 -28962
rect 27016 -29042 27096 -28962
rect 27136 -29042 27216 -28962
rect 27256 -29042 27336 -28962
rect 27376 -29042 27456 -28962
rect 27496 -29042 27576 -28962
rect 27616 -29042 27696 -28962
rect 27736 -29042 27816 -28962
rect 27856 -29042 27936 -28962
rect 27976 -29042 28056 -28962
rect 28096 -29042 28176 -28962
rect 28216 -29042 28296 -28962
rect 28336 -29042 28416 -28962
rect 28456 -29042 28536 -28962
rect 28576 -29042 28656 -28962
rect 28696 -29042 28776 -28962
rect 28816 -29042 28896 -28962
rect 28936 -29042 29016 -28962
rect 29056 -29042 29136 -28962
rect 29176 -29042 29256 -28962
rect 29296 -29042 29376 -28962
rect 29416 -29042 29496 -28962
rect 29536 -29042 29616 -28962
rect 29656 -29042 29736 -28962
rect 29776 -29042 29856 -28962
rect 29896 -29042 29976 -28962
rect 30016 -29042 30096 -28962
rect 23656 -29162 23736 -29082
rect 23776 -29162 23856 -29082
rect 23896 -29162 23976 -29082
rect 24016 -29162 24096 -29082
rect 24136 -29162 24216 -29082
rect 24256 -29162 24336 -29082
rect 24376 -29162 24456 -29082
rect 24496 -29162 24576 -29082
rect 24616 -29162 24696 -29082
rect 24736 -29162 24816 -29082
rect 24856 -29162 24936 -29082
rect 24976 -29162 25056 -29082
rect 25096 -29162 25176 -29082
rect 25216 -29162 25296 -29082
rect 25336 -29162 25416 -29082
rect 25456 -29162 25536 -29082
rect 25576 -29162 25656 -29082
rect 25696 -29162 25776 -29082
rect 25816 -29162 25896 -29082
rect 25936 -29162 26016 -29082
rect 26056 -29162 26136 -29082
rect 26176 -29162 26256 -29082
rect 26296 -29162 26376 -29082
rect 26416 -29162 26496 -29082
rect 26536 -29162 26616 -29082
rect 26656 -29162 26736 -29082
rect 26776 -29162 26856 -29082
rect 26896 -29162 26976 -29082
rect 27016 -29162 27096 -29082
rect 27136 -29162 27216 -29082
rect 27256 -29162 27336 -29082
rect 27376 -29162 27456 -29082
rect 27496 -29162 27576 -29082
rect 27616 -29162 27696 -29082
rect 27736 -29162 27816 -29082
rect 27856 -29162 27936 -29082
rect 27976 -29162 28056 -29082
rect 28096 -29162 28176 -29082
rect 28216 -29162 28296 -29082
rect 28336 -29162 28416 -29082
rect 28456 -29162 28536 -29082
rect 28576 -29162 28656 -29082
rect 28696 -29162 28776 -29082
rect 28816 -29162 28896 -29082
rect 28936 -29162 29016 -29082
rect 29056 -29162 29136 -29082
rect 29176 -29162 29256 -29082
rect 29296 -29162 29376 -29082
rect 29416 -29162 29496 -29082
rect 29536 -29162 29616 -29082
rect 29656 -29162 29736 -29082
rect 29776 -29162 29856 -29082
rect 29896 -29162 29976 -29082
rect 30016 -29162 30096 -29082
<< metal1 >>
rect 23636 -18922 30156 -18902
rect 23636 -19002 23656 -18922
rect 23736 -19002 23776 -18922
rect 23856 -19002 23896 -18922
rect 23976 -19002 24016 -18922
rect 24096 -19002 24136 -18922
rect 24216 -19002 24256 -18922
rect 24336 -19002 24376 -18922
rect 24456 -19002 24496 -18922
rect 24576 -19002 24616 -18922
rect 24696 -19002 24736 -18922
rect 24816 -19002 24856 -18922
rect 24936 -19002 24976 -18922
rect 25056 -19002 25096 -18922
rect 25176 -19002 25216 -18922
rect 25296 -19002 25336 -18922
rect 25416 -19002 25456 -18922
rect 25536 -19002 25576 -18922
rect 25656 -19002 25696 -18922
rect 25776 -19002 25816 -18922
rect 25896 -19002 25936 -18922
rect 26016 -19002 26056 -18922
rect 26136 -19002 26176 -18922
rect 26256 -19002 26296 -18922
rect 26376 -19002 26416 -18922
rect 26496 -19002 26536 -18922
rect 26616 -19002 26656 -18922
rect 26736 -19002 26776 -18922
rect 26856 -19002 26896 -18922
rect 26976 -19002 27016 -18922
rect 27096 -19002 27136 -18922
rect 27216 -19002 27256 -18922
rect 27336 -19002 27376 -18922
rect 27456 -19002 27496 -18922
rect 27576 -19002 27616 -18922
rect 27696 -19002 27736 -18922
rect 27816 -19002 27856 -18922
rect 27936 -19002 27976 -18922
rect 28056 -19002 28096 -18922
rect 28176 -19002 28216 -18922
rect 28296 -19002 28336 -18922
rect 28416 -19002 28456 -18922
rect 28536 -19002 28576 -18922
rect 28656 -19002 28696 -18922
rect 28776 -19002 28816 -18922
rect 28896 -19002 28936 -18922
rect 29016 -19002 29056 -18922
rect 29136 -19002 29176 -18922
rect 29256 -19002 29296 -18922
rect 29376 -19002 29416 -18922
rect 29496 -19002 29536 -18922
rect 29616 -19002 29656 -18922
rect 29736 -19002 29776 -18922
rect 29856 -19002 29896 -18922
rect 29976 -19002 30016 -18922
rect 30096 -19002 30156 -18922
rect 23636 -19042 30156 -19002
rect 23636 -19122 23656 -19042
rect 23736 -19122 23776 -19042
rect 23856 -19122 23896 -19042
rect 23976 -19122 24016 -19042
rect 24096 -19122 24136 -19042
rect 24216 -19122 24256 -19042
rect 24336 -19122 24376 -19042
rect 24456 -19122 24496 -19042
rect 24576 -19122 24616 -19042
rect 24696 -19122 24736 -19042
rect 24816 -19122 24856 -19042
rect 24936 -19122 24976 -19042
rect 25056 -19122 25096 -19042
rect 25176 -19122 25216 -19042
rect 25296 -19122 25336 -19042
rect 25416 -19122 25456 -19042
rect 25536 -19122 25576 -19042
rect 25656 -19122 25696 -19042
rect 25776 -19122 25816 -19042
rect 25896 -19122 25936 -19042
rect 26016 -19122 26056 -19042
rect 26136 -19122 26176 -19042
rect 26256 -19122 26296 -19042
rect 26376 -19122 26416 -19042
rect 26496 -19122 26536 -19042
rect 26616 -19122 26656 -19042
rect 26736 -19122 26776 -19042
rect 26856 -19122 26896 -19042
rect 26976 -19122 27016 -19042
rect 27096 -19122 27136 -19042
rect 27216 -19122 27256 -19042
rect 27336 -19122 27376 -19042
rect 27456 -19122 27496 -19042
rect 27576 -19122 27616 -19042
rect 27696 -19122 27736 -19042
rect 27816 -19122 27856 -19042
rect 27936 -19122 27976 -19042
rect 28056 -19122 28096 -19042
rect 28176 -19122 28216 -19042
rect 28296 -19122 28336 -19042
rect 28416 -19122 28456 -19042
rect 28536 -19122 28576 -19042
rect 28656 -19122 28696 -19042
rect 28776 -19122 28816 -19042
rect 28896 -19122 28936 -19042
rect 29016 -19122 29056 -19042
rect 29136 -19122 29176 -19042
rect 29256 -19122 29296 -19042
rect 29376 -19122 29416 -19042
rect 29496 -19122 29536 -19042
rect 29616 -19122 29656 -19042
rect 29736 -19122 29776 -19042
rect 29856 -19122 29896 -19042
rect 29976 -19122 30016 -19042
rect 30096 -19122 30156 -19042
rect 23636 -19162 30156 -19122
rect 23636 -19242 23656 -19162
rect 23736 -19242 23776 -19162
rect 23856 -19242 23896 -19162
rect 23976 -19242 24016 -19162
rect 24096 -19242 24136 -19162
rect 24216 -19242 24256 -19162
rect 24336 -19242 24376 -19162
rect 24456 -19242 24496 -19162
rect 24576 -19242 24616 -19162
rect 24696 -19242 24736 -19162
rect 24816 -19242 24856 -19162
rect 24936 -19242 24976 -19162
rect 25056 -19242 25096 -19162
rect 25176 -19242 25216 -19162
rect 25296 -19242 25336 -19162
rect 25416 -19242 25456 -19162
rect 25536 -19242 25576 -19162
rect 25656 -19242 25696 -19162
rect 25776 -19242 25816 -19162
rect 25896 -19242 25936 -19162
rect 26016 -19242 26056 -19162
rect 26136 -19242 26176 -19162
rect 26256 -19242 26296 -19162
rect 26376 -19242 26416 -19162
rect 26496 -19242 26536 -19162
rect 26616 -19242 26656 -19162
rect 26736 -19242 26776 -19162
rect 26856 -19242 26896 -19162
rect 26976 -19242 27016 -19162
rect 27096 -19242 27136 -19162
rect 27216 -19242 27256 -19162
rect 27336 -19242 27376 -19162
rect 27456 -19242 27496 -19162
rect 27576 -19242 27616 -19162
rect 27696 -19242 27736 -19162
rect 27816 -19242 27856 -19162
rect 27936 -19242 27976 -19162
rect 28056 -19242 28096 -19162
rect 28176 -19242 28216 -19162
rect 28296 -19242 28336 -19162
rect 28416 -19242 28456 -19162
rect 28536 -19242 28576 -19162
rect 28656 -19242 28696 -19162
rect 28776 -19242 28816 -19162
rect 28896 -19242 28936 -19162
rect 29016 -19242 29056 -19162
rect 29136 -19242 29176 -19162
rect 29256 -19242 29296 -19162
rect 29376 -19242 29416 -19162
rect 29496 -19242 29536 -19162
rect 29616 -19242 29656 -19162
rect 29736 -19242 29776 -19162
rect 29856 -19242 29896 -19162
rect 29976 -19242 30016 -19162
rect 30096 -19242 30156 -19162
rect 23636 -19282 30156 -19242
rect 23636 -19362 23656 -19282
rect 23736 -19362 23776 -19282
rect 23856 -19362 23896 -19282
rect 23976 -19362 24016 -19282
rect 24096 -19362 24136 -19282
rect 24216 -19362 24256 -19282
rect 24336 -19362 24376 -19282
rect 24456 -19362 24496 -19282
rect 24576 -19362 24616 -19282
rect 24696 -19362 24736 -19282
rect 24816 -19362 24856 -19282
rect 24936 -19362 24976 -19282
rect 25056 -19362 25096 -19282
rect 25176 -19362 25216 -19282
rect 25296 -19362 25336 -19282
rect 25416 -19362 25456 -19282
rect 25536 -19362 25576 -19282
rect 25656 -19362 25696 -19282
rect 25776 -19362 25816 -19282
rect 25896 -19362 25936 -19282
rect 26016 -19362 26056 -19282
rect 26136 -19362 26176 -19282
rect 26256 -19362 26296 -19282
rect 26376 -19362 26416 -19282
rect 26496 -19362 26536 -19282
rect 26616 -19362 26656 -19282
rect 26736 -19362 26776 -19282
rect 26856 -19362 26896 -19282
rect 26976 -19362 27016 -19282
rect 27096 -19362 27136 -19282
rect 27216 -19362 27256 -19282
rect 27336 -19362 27376 -19282
rect 27456 -19362 27496 -19282
rect 27576 -19362 27616 -19282
rect 27696 -19362 27736 -19282
rect 27816 -19362 27856 -19282
rect 27936 -19362 27976 -19282
rect 28056 -19362 28096 -19282
rect 28176 -19362 28216 -19282
rect 28296 -19362 28336 -19282
rect 28416 -19362 28456 -19282
rect 28536 -19362 28576 -19282
rect 28656 -19362 28696 -19282
rect 28776 -19362 28816 -19282
rect 28896 -19362 28936 -19282
rect 29016 -19362 29056 -19282
rect 29136 -19362 29176 -19282
rect 29256 -19362 29296 -19282
rect 29376 -19362 29416 -19282
rect 29496 -19362 29536 -19282
rect 29616 -19362 29656 -19282
rect 29736 -19362 29776 -19282
rect 29856 -19362 29896 -19282
rect 29976 -19362 30016 -19282
rect 30096 -19362 30156 -19282
rect 23636 -19402 30156 -19362
rect 23636 -19482 23656 -19402
rect 23736 -19482 23776 -19402
rect 23856 -19482 23896 -19402
rect 23976 -19482 24016 -19402
rect 24096 -19482 24136 -19402
rect 24216 -19482 24256 -19402
rect 24336 -19482 24376 -19402
rect 24456 -19482 24496 -19402
rect 24576 -19482 24616 -19402
rect 24696 -19482 24736 -19402
rect 24816 -19482 24856 -19402
rect 24936 -19482 24976 -19402
rect 25056 -19482 25096 -19402
rect 25176 -19482 25216 -19402
rect 25296 -19482 25336 -19402
rect 25416 -19482 25456 -19402
rect 25536 -19482 25576 -19402
rect 25656 -19482 25696 -19402
rect 25776 -19482 25816 -19402
rect 25896 -19482 25936 -19402
rect 26016 -19482 26056 -19402
rect 26136 -19482 26176 -19402
rect 26256 -19482 26296 -19402
rect 26376 -19482 26416 -19402
rect 26496 -19482 26536 -19402
rect 26616 -19482 26656 -19402
rect 26736 -19482 26776 -19402
rect 26856 -19482 26896 -19402
rect 26976 -19482 27016 -19402
rect 27096 -19482 27136 -19402
rect 27216 -19482 27256 -19402
rect 27336 -19482 27376 -19402
rect 27456 -19482 27496 -19402
rect 27576 -19482 27616 -19402
rect 27696 -19482 27736 -19402
rect 27816 -19482 27856 -19402
rect 27936 -19482 27976 -19402
rect 28056 -19482 28096 -19402
rect 28176 -19482 28216 -19402
rect 28296 -19482 28336 -19402
rect 28416 -19482 28456 -19402
rect 28536 -19482 28576 -19402
rect 28656 -19482 28696 -19402
rect 28776 -19482 28816 -19402
rect 28896 -19482 28936 -19402
rect 29016 -19482 29056 -19402
rect 29136 -19482 29176 -19402
rect 29256 -19482 29296 -19402
rect 29376 -19482 29416 -19402
rect 29496 -19482 29536 -19402
rect 29616 -19482 29656 -19402
rect 29736 -19482 29776 -19402
rect 29856 -19482 29896 -19402
rect 29976 -19482 30016 -19402
rect 30096 -19482 30156 -19402
rect 23636 -19522 30156 -19482
rect 23636 -19602 23656 -19522
rect 23736 -19602 23776 -19522
rect 23856 -19602 23896 -19522
rect 23976 -19602 24016 -19522
rect 24096 -19602 24136 -19522
rect 24216 -19602 24256 -19522
rect 24336 -19602 24376 -19522
rect 24456 -19602 24496 -19522
rect 24576 -19602 24616 -19522
rect 24696 -19602 24736 -19522
rect 24816 -19602 24856 -19522
rect 24936 -19602 24976 -19522
rect 25056 -19602 25096 -19522
rect 25176 -19602 25216 -19522
rect 25296 -19602 25336 -19522
rect 25416 -19602 25456 -19522
rect 25536 -19602 25576 -19522
rect 25656 -19602 25696 -19522
rect 25776 -19602 25816 -19522
rect 25896 -19602 25936 -19522
rect 26016 -19602 26056 -19522
rect 26136 -19602 26176 -19522
rect 26256 -19602 26296 -19522
rect 26376 -19602 26416 -19522
rect 26496 -19602 26536 -19522
rect 26616 -19602 26656 -19522
rect 26736 -19602 26776 -19522
rect 26856 -19602 26896 -19522
rect 26976 -19602 27016 -19522
rect 27096 -19602 27136 -19522
rect 27216 -19602 27256 -19522
rect 27336 -19602 27376 -19522
rect 27456 -19602 27496 -19522
rect 27576 -19602 27616 -19522
rect 27696 -19602 27736 -19522
rect 27816 -19602 27856 -19522
rect 27936 -19602 27976 -19522
rect 28056 -19602 28096 -19522
rect 28176 -19602 28216 -19522
rect 28296 -19602 28336 -19522
rect 28416 -19602 28456 -19522
rect 28536 -19602 28576 -19522
rect 28656 -19602 28696 -19522
rect 28776 -19602 28816 -19522
rect 28896 -19602 28936 -19522
rect 29016 -19602 29056 -19522
rect 29136 -19602 29176 -19522
rect 29256 -19602 29296 -19522
rect 29376 -19602 29416 -19522
rect 29496 -19602 29536 -19522
rect 29616 -19602 29656 -19522
rect 29736 -19602 29776 -19522
rect 29856 -19602 29896 -19522
rect 29976 -19602 30016 -19522
rect 30096 -19602 30156 -19522
rect 23636 -19622 30156 -19602
rect 23908 -19874 23954 -19862
rect 20908 -20234 20954 -20222
rect 20908 -21882 20914 -20234
rect 20876 -21902 20914 -21882
rect 20948 -21882 20954 -20234
rect 21216 -20234 21262 -20222
rect 20948 -21902 20996 -21882
rect 20876 -21962 20896 -21902
rect 20956 -21962 20996 -21902
rect 20876 -22082 20914 -21962
rect 20948 -22082 20996 -21962
rect 20876 -22142 20896 -22082
rect 20956 -22142 20996 -22082
rect 20876 -22162 20914 -22142
rect 20908 -22210 20914 -22162
rect 20948 -22162 20996 -22142
rect 20948 -22210 20954 -22162
rect 20908 -22222 20954 -22210
rect 21216 -22210 21222 -20234
rect 21256 -22210 21262 -20234
rect 21524 -20234 21570 -20222
rect 21524 -21882 21530 -20234
rect 21476 -21902 21530 -21882
rect 21564 -21882 21570 -20234
rect 21832 -20234 21878 -20222
rect 21476 -21962 21496 -21902
rect 21476 -22082 21530 -21962
rect 21476 -22142 21496 -22082
rect 21476 -22162 21530 -22142
rect 21216 -22222 21262 -22210
rect 21524 -22210 21530 -22162
rect 21564 -22162 21596 -21882
rect 21564 -22210 21570 -22162
rect 21524 -22222 21570 -22210
rect 21832 -22210 21838 -20234
rect 21872 -22210 21878 -20234
rect 22140 -20234 22186 -20222
rect 22140 -21882 22146 -20234
rect 22096 -21902 22146 -21882
rect 22180 -21882 22186 -20234
rect 22448 -20234 22494 -20222
rect 22180 -21902 22216 -21882
rect 22096 -21962 22136 -21902
rect 22196 -21962 22216 -21902
rect 22096 -22082 22146 -21962
rect 22180 -22082 22216 -21962
rect 22096 -22142 22136 -22082
rect 22196 -22142 22216 -22082
rect 22096 -22162 22146 -22142
rect 21832 -22222 21878 -22210
rect 22140 -22210 22146 -22162
rect 22180 -22162 22216 -22142
rect 22180 -22210 22186 -22162
rect 22140 -22222 22186 -22210
rect 22448 -22210 22454 -20234
rect 22488 -22210 22494 -20234
rect 22756 -20234 22802 -20222
rect 22756 -21882 22762 -20234
rect 22716 -21902 22762 -21882
rect 22796 -21882 22802 -20234
rect 23064 -20234 23110 -20222
rect 22716 -21962 22736 -21902
rect 22716 -22082 22762 -21962
rect 22716 -22142 22736 -22082
rect 22716 -22162 22762 -22142
rect 22448 -22222 22494 -22210
rect 22756 -22210 22762 -22162
rect 22796 -22162 22836 -21882
rect 22796 -22210 22802 -22162
rect 22756 -22222 22802 -22210
rect 23064 -22210 23070 -20234
rect 23104 -22210 23110 -20234
rect 23372 -20234 23418 -20222
rect 23372 -21882 23378 -20234
rect 23336 -21902 23378 -21882
rect 23412 -21882 23418 -20234
rect 23908 -21730 23914 -19874
rect 23948 -21730 23954 -19874
rect 23908 -21742 23954 -21730
rect 24066 -19874 24112 -19862
rect 24066 -21730 24072 -19874
rect 24106 -21730 24112 -19874
rect 24066 -21742 24112 -21730
rect 24224 -19874 24270 -19862
rect 24224 -21730 24230 -19874
rect 24264 -21730 24270 -19874
rect 29448 -19874 29494 -19862
rect 24343 -20065 24389 -20053
rect 24343 -21549 24349 -20065
rect 24383 -21549 24389 -20065
rect 24343 -21561 24389 -21549
rect 24651 -20065 24697 -20053
rect 24651 -21549 24657 -20065
rect 24691 -21549 24697 -20065
rect 24959 -20065 25005 -20053
rect 24959 -20982 24965 -20065
rect 24876 -21002 24965 -20982
rect 24999 -20982 25005 -20065
rect 25267 -20065 25313 -20053
rect 24999 -21002 25076 -20982
rect 24876 -21062 24896 -21002
rect 24956 -21062 24965 -21002
rect 25056 -21062 25076 -21002
rect 24876 -21082 24965 -21062
rect 24999 -21082 25076 -21062
rect 24876 -21142 24896 -21082
rect 24956 -21142 24965 -21082
rect 25056 -21142 25076 -21082
rect 24876 -21202 24965 -21142
rect 24999 -21202 25076 -21142
rect 24876 -21262 24896 -21202
rect 24956 -21262 24965 -21202
rect 25056 -21262 25076 -21202
rect 24876 -21282 24965 -21262
rect 24999 -21282 25076 -21262
rect 24876 -21342 24896 -21282
rect 24956 -21342 24965 -21282
rect 25056 -21342 25076 -21282
rect 24876 -21362 24965 -21342
rect 24651 -21561 24697 -21549
rect 24959 -21549 24965 -21362
rect 24999 -21362 25076 -21342
rect 24999 -21549 25005 -21362
rect 24959 -21561 25005 -21549
rect 25267 -21549 25273 -20065
rect 25307 -21549 25313 -20065
rect 25267 -21561 25313 -21549
rect 25575 -20065 25621 -20053
rect 25575 -21549 25581 -20065
rect 25615 -21549 25621 -20065
rect 25575 -21561 25621 -21549
rect 25883 -20065 25929 -20053
rect 25883 -21549 25889 -20065
rect 25923 -21549 25929 -20065
rect 26191 -20065 26237 -20053
rect 26191 -20982 26197 -20065
rect 26116 -21002 26197 -20982
rect 26116 -21062 26136 -21002
rect 26196 -21062 26197 -21002
rect 26116 -21082 26197 -21062
rect 26116 -21142 26136 -21082
rect 26196 -21142 26197 -21082
rect 26116 -21202 26197 -21142
rect 26116 -21262 26136 -21202
rect 26196 -21262 26197 -21202
rect 26116 -21282 26197 -21262
rect 26116 -21342 26136 -21282
rect 26196 -21342 26197 -21282
rect 26116 -21362 26197 -21342
rect 25883 -21561 25929 -21549
rect 26191 -21549 26197 -21362
rect 26231 -20982 26237 -20065
rect 26499 -20065 26545 -20053
rect 26231 -21002 26316 -20982
rect 26231 -21062 26236 -21002
rect 26296 -21062 26316 -21002
rect 26231 -21082 26316 -21062
rect 26231 -21142 26236 -21082
rect 26296 -21142 26316 -21082
rect 26231 -21202 26316 -21142
rect 26231 -21262 26236 -21202
rect 26296 -21262 26316 -21202
rect 26231 -21282 26316 -21262
rect 26231 -21342 26236 -21282
rect 26296 -21342 26316 -21282
rect 26231 -21362 26316 -21342
rect 26231 -21549 26237 -21362
rect 26191 -21561 26237 -21549
rect 26499 -21549 26505 -20065
rect 26539 -21549 26545 -20065
rect 26499 -21561 26545 -21549
rect 26807 -20065 26853 -20053
rect 26807 -21549 26813 -20065
rect 26847 -21549 26853 -20065
rect 26807 -21561 26853 -21549
rect 27115 -20065 27161 -20053
rect 27115 -21549 27121 -20065
rect 27155 -21549 27161 -20065
rect 27423 -20065 27469 -20053
rect 27423 -20982 27429 -20065
rect 27336 -21002 27429 -20982
rect 27463 -20982 27469 -20065
rect 27731 -20065 27777 -20053
rect 27463 -21002 27536 -20982
rect 27336 -21062 27356 -21002
rect 27416 -21062 27429 -21002
rect 27516 -21062 27536 -21002
rect 27336 -21082 27429 -21062
rect 27463 -21082 27536 -21062
rect 27336 -21142 27356 -21082
rect 27416 -21142 27429 -21082
rect 27516 -21142 27536 -21082
rect 27336 -21202 27429 -21142
rect 27463 -21202 27536 -21142
rect 27336 -21262 27356 -21202
rect 27416 -21262 27429 -21202
rect 27516 -21262 27536 -21202
rect 27336 -21282 27429 -21262
rect 27463 -21282 27536 -21262
rect 27336 -21342 27356 -21282
rect 27416 -21342 27429 -21282
rect 27516 -21342 27536 -21282
rect 27336 -21362 27429 -21342
rect 27115 -21561 27161 -21549
rect 27423 -21549 27429 -21362
rect 27463 -21362 27536 -21342
rect 27463 -21549 27469 -21362
rect 27423 -21561 27469 -21549
rect 27731 -21549 27737 -20065
rect 27771 -21549 27777 -20065
rect 27731 -21561 27777 -21549
rect 28039 -20065 28085 -20053
rect 28039 -21549 28045 -20065
rect 28079 -21549 28085 -20065
rect 28039 -21561 28085 -21549
rect 28347 -20065 28393 -20053
rect 28347 -21549 28353 -20065
rect 28387 -21549 28393 -20065
rect 28655 -20065 28701 -20053
rect 28655 -20982 28661 -20065
rect 28576 -21002 28661 -20982
rect 28576 -21062 28596 -21002
rect 28656 -21062 28661 -21002
rect 28576 -21082 28661 -21062
rect 28576 -21142 28596 -21082
rect 28656 -21142 28661 -21082
rect 28576 -21202 28661 -21142
rect 28576 -21262 28596 -21202
rect 28656 -21262 28661 -21202
rect 28576 -21282 28661 -21262
rect 28576 -21342 28596 -21282
rect 28656 -21342 28661 -21282
rect 28576 -21362 28661 -21342
rect 28347 -21561 28393 -21549
rect 28655 -21549 28661 -21362
rect 28695 -20982 28701 -20065
rect 28963 -20065 29009 -20053
rect 28695 -21002 28776 -20982
rect 28695 -21062 28696 -21002
rect 28756 -21062 28776 -21002
rect 28695 -21082 28776 -21062
rect 28695 -21142 28696 -21082
rect 28756 -21142 28776 -21082
rect 28695 -21202 28776 -21142
rect 28695 -21262 28696 -21202
rect 28756 -21262 28776 -21202
rect 28695 -21282 28776 -21262
rect 28695 -21342 28696 -21282
rect 28756 -21342 28776 -21282
rect 28695 -21362 28776 -21342
rect 28695 -21549 28701 -21362
rect 28655 -21561 28701 -21549
rect 28963 -21549 28969 -20065
rect 29003 -21549 29009 -20065
rect 28963 -21561 29009 -21549
rect 29271 -20065 29317 -20053
rect 29271 -21549 29277 -20065
rect 29311 -21549 29317 -20065
rect 29271 -21561 29317 -21549
rect 24224 -21742 24270 -21730
rect 23964 -21789 24056 -21783
rect 23964 -21823 23976 -21789
rect 24044 -21823 24056 -21789
rect 23964 -21829 24056 -21823
rect 24122 -21789 24214 -21783
rect 24122 -21823 24134 -21789
rect 24202 -21823 24214 -21789
rect 24122 -21829 24214 -21823
rect 24356 -21794 29356 -21642
rect 29448 -21730 29454 -19874
rect 29488 -21730 29494 -19874
rect 29448 -21742 29494 -21730
rect 29606 -19874 29652 -19862
rect 29606 -21730 29612 -19874
rect 29646 -21730 29652 -19874
rect 29606 -21742 29652 -21730
rect 29764 -19874 29810 -19862
rect 29764 -21730 29770 -19874
rect 29804 -21730 29810 -19874
rect 29764 -21742 29810 -21730
rect 30348 -20234 30394 -20222
rect 24356 -21828 24411 -21794
rect 24629 -21828 24719 -21794
rect 24937 -21828 25027 -21794
rect 25245 -21828 25335 -21794
rect 25553 -21828 25643 -21794
rect 25861 -21828 25951 -21794
rect 26169 -21828 26259 -21794
rect 26477 -21828 26567 -21794
rect 26785 -21828 26875 -21794
rect 27093 -21828 27183 -21794
rect 27401 -21828 27491 -21794
rect 27709 -21828 27799 -21794
rect 28017 -21828 28107 -21794
rect 28325 -21828 28415 -21794
rect 28633 -21828 28723 -21794
rect 28941 -21828 29031 -21794
rect 29249 -21828 29356 -21794
rect 24356 -21842 29356 -21828
rect 29504 -21789 29596 -21783
rect 29504 -21823 29516 -21789
rect 29584 -21823 29596 -21789
rect 29504 -21829 29596 -21823
rect 29662 -21789 29754 -21783
rect 29662 -21823 29674 -21789
rect 29742 -21823 29754 -21789
rect 29662 -21829 29754 -21823
rect 23412 -21902 23456 -21882
rect 23336 -21962 23376 -21902
rect 23436 -21962 23456 -21902
rect 23336 -22082 23378 -21962
rect 23412 -22082 23456 -21962
rect 23336 -22142 23376 -22082
rect 23436 -22142 23456 -22082
rect 23336 -22162 23378 -22142
rect 23064 -22222 23110 -22210
rect 23372 -22210 23378 -22162
rect 23412 -22162 23456 -22142
rect 24616 -21962 29176 -21842
rect 30348 -21882 30354 -20234
rect 24616 -22042 24636 -21962
rect 24716 -22042 24756 -21962
rect 24836 -22042 24876 -21962
rect 24956 -22042 24996 -21962
rect 25076 -22042 25116 -21962
rect 25196 -22042 25236 -21962
rect 25316 -22042 25356 -21962
rect 25436 -22042 25476 -21962
rect 25556 -22042 25596 -21962
rect 25676 -22042 25716 -21962
rect 25796 -22042 25836 -21962
rect 25916 -22042 25956 -21962
rect 26036 -22042 26076 -21962
rect 26156 -22042 26196 -21962
rect 26276 -22042 26316 -21962
rect 26396 -22042 26436 -21962
rect 26516 -22042 26556 -21962
rect 26636 -22042 26676 -21962
rect 26756 -22042 26796 -21962
rect 26876 -22042 26916 -21962
rect 26996 -22042 27036 -21962
rect 27116 -22042 27156 -21962
rect 27236 -22042 27276 -21962
rect 27356 -22042 27396 -21962
rect 27476 -22042 27516 -21962
rect 27596 -22042 27636 -21962
rect 27716 -22042 27756 -21962
rect 27836 -22042 27876 -21962
rect 27956 -22042 27996 -21962
rect 28076 -22042 28116 -21962
rect 28196 -22042 28236 -21962
rect 28316 -22042 28356 -21962
rect 28436 -22042 28476 -21962
rect 28556 -22042 28596 -21962
rect 28676 -22042 28716 -21962
rect 28796 -22042 28836 -21962
rect 28916 -22042 28956 -21962
rect 29036 -22042 29076 -21962
rect 29156 -22042 29176 -21962
rect 24616 -22102 29176 -22042
rect 23412 -22210 23418 -22162
rect 23372 -22222 23418 -22210
rect 24616 -22182 24636 -22102
rect 24716 -22182 24756 -22102
rect 24836 -22182 24876 -22102
rect 24956 -22182 24996 -22102
rect 25076 -22182 25116 -22102
rect 25196 -22182 25236 -22102
rect 25316 -22182 25356 -22102
rect 25436 -22182 25476 -22102
rect 25556 -22182 25596 -22102
rect 25676 -22182 25716 -22102
rect 25796 -22182 25836 -22102
rect 25916 -22182 25956 -22102
rect 26036 -22182 26076 -22102
rect 26156 -22182 26196 -22102
rect 26276 -22182 26316 -22102
rect 26396 -22182 26436 -22102
rect 26516 -22182 26556 -22102
rect 26636 -22182 26676 -22102
rect 26756 -22182 26796 -22102
rect 26876 -22182 26916 -22102
rect 26996 -22182 27036 -22102
rect 27116 -22182 27156 -22102
rect 27236 -22182 27276 -22102
rect 27356 -22182 27396 -22102
rect 27476 -22182 27516 -22102
rect 27596 -22182 27636 -22102
rect 27716 -22182 27756 -22102
rect 27836 -22182 27876 -22102
rect 27956 -22182 27996 -22102
rect 28076 -22182 28116 -22102
rect 28196 -22182 28236 -22102
rect 28316 -22182 28356 -22102
rect 28436 -22182 28476 -22102
rect 28556 -22182 28596 -22102
rect 28676 -22182 28716 -22102
rect 28796 -22182 28836 -22102
rect 28916 -22182 28956 -22102
rect 29036 -22182 29076 -22102
rect 29156 -22182 29176 -22102
rect 30316 -21902 30354 -21882
rect 30388 -21882 30394 -20234
rect 30656 -20234 30702 -20222
rect 30388 -21902 30436 -21882
rect 30316 -21962 30336 -21902
rect 30396 -21962 30436 -21902
rect 30316 -22082 30354 -21962
rect 30388 -22082 30436 -21962
rect 30316 -22142 30336 -22082
rect 30396 -22142 30436 -22082
rect 30316 -22162 30354 -22142
rect 24616 -22242 29176 -22182
rect 30348 -22210 30354 -22162
rect 30388 -22162 30436 -22142
rect 30388 -22210 30394 -22162
rect 30348 -22222 30394 -22210
rect 30656 -22210 30662 -20234
rect 30696 -22210 30702 -20234
rect 30964 -20234 31010 -20222
rect 30964 -21882 30970 -20234
rect 30916 -21902 30970 -21882
rect 31004 -21882 31010 -20234
rect 31272 -20234 31318 -20222
rect 30916 -21962 30936 -21902
rect 30916 -22082 30970 -21962
rect 30916 -22142 30936 -22082
rect 30916 -22162 30970 -22142
rect 30656 -22222 30702 -22210
rect 30964 -22210 30970 -22162
rect 31004 -22162 31036 -21882
rect 31004 -22210 31010 -22162
rect 30964 -22222 31010 -22210
rect 31272 -22210 31278 -20234
rect 31312 -22210 31318 -20234
rect 31580 -20234 31626 -20222
rect 31580 -21882 31586 -20234
rect 31536 -21902 31586 -21882
rect 31620 -21882 31626 -20234
rect 31888 -20234 31934 -20222
rect 31620 -21902 31656 -21882
rect 31536 -21962 31576 -21902
rect 31636 -21962 31656 -21902
rect 31536 -22082 31586 -21962
rect 31620 -22082 31656 -21962
rect 31536 -22142 31576 -22082
rect 31636 -22142 31656 -22082
rect 31536 -22162 31586 -22142
rect 31272 -22222 31318 -22210
rect 31580 -22210 31586 -22162
rect 31620 -22162 31656 -22142
rect 31620 -22210 31626 -22162
rect 31580 -22222 31626 -22210
rect 31888 -22210 31894 -20234
rect 31928 -22210 31934 -20234
rect 32196 -20234 32242 -20222
rect 32196 -21882 32202 -20234
rect 32156 -21902 32202 -21882
rect 32236 -21882 32242 -20234
rect 32504 -20234 32550 -20222
rect 32156 -21962 32176 -21902
rect 32156 -22082 32202 -21962
rect 32156 -22142 32176 -22082
rect 32156 -22162 32202 -22142
rect 31888 -22222 31934 -22210
rect 32196 -22210 32202 -22162
rect 32236 -22162 32276 -21882
rect 32236 -22210 32242 -22162
rect 32196 -22222 32242 -22210
rect 32504 -22210 32510 -20234
rect 32544 -22210 32550 -20234
rect 32812 -20234 32858 -20222
rect 32812 -21882 32818 -20234
rect 32776 -21902 32818 -21882
rect 32852 -21882 32858 -20234
rect 32852 -21902 32896 -21882
rect 32776 -21962 32796 -21902
rect 32856 -21962 32896 -21902
rect 32776 -22082 32818 -21962
rect 32852 -22082 32896 -21962
rect 32776 -22142 32796 -22082
rect 32856 -22142 32896 -22082
rect 32776 -22162 32818 -22142
rect 32504 -22222 32550 -22210
rect 32812 -22210 32818 -22162
rect 32852 -22162 32896 -22142
rect 32852 -22210 32858 -22162
rect 32812 -22222 32858 -22210
rect 20964 -22269 21206 -22263
rect 20964 -22282 20976 -22269
rect 20956 -22303 20976 -22282
rect 21194 -22282 21206 -22269
rect 21272 -22269 21514 -22263
rect 21272 -22282 21284 -22269
rect 21194 -22303 21284 -22282
rect 21502 -22282 21514 -22269
rect 21580 -22269 21822 -22263
rect 21580 -22282 21592 -22269
rect 21502 -22303 21592 -22282
rect 21810 -22282 21822 -22269
rect 21888 -22269 22130 -22263
rect 21888 -22282 21900 -22269
rect 21810 -22303 21900 -22282
rect 22118 -22282 22130 -22269
rect 22196 -22269 22438 -22263
rect 22196 -22282 22208 -22269
rect 22118 -22303 22208 -22282
rect 22426 -22282 22438 -22269
rect 22504 -22269 22746 -22263
rect 22504 -22282 22516 -22269
rect 22426 -22303 22516 -22282
rect 22734 -22282 22746 -22269
rect 22812 -22269 23054 -22263
rect 22812 -22282 22824 -22269
rect 22734 -22303 22824 -22282
rect 23042 -22282 23054 -22269
rect 23120 -22269 23362 -22263
rect 23120 -22282 23132 -22269
rect 23042 -22303 23132 -22282
rect 23350 -22282 23362 -22269
rect 23350 -22303 23376 -22282
rect 20956 -22442 23376 -22303
rect 24616 -22322 24636 -22242
rect 24716 -22322 24756 -22242
rect 24836 -22322 24876 -22242
rect 24956 -22322 24996 -22242
rect 25076 -22322 25116 -22242
rect 25196 -22322 25236 -22242
rect 25316 -22322 25356 -22242
rect 25436 -22322 25476 -22242
rect 25556 -22322 25596 -22242
rect 25676 -22322 25716 -22242
rect 25796 -22322 25836 -22242
rect 25916 -22322 25956 -22242
rect 26036 -22322 26076 -22242
rect 26156 -22322 26196 -22242
rect 26276 -22322 26316 -22242
rect 26396 -22322 26436 -22242
rect 26516 -22322 26556 -22242
rect 26636 -22322 26676 -22242
rect 26756 -22322 26796 -22242
rect 26876 -22322 26916 -22242
rect 26996 -22322 27036 -22242
rect 27116 -22322 27156 -22242
rect 27236 -22322 27276 -22242
rect 27356 -22322 27396 -22242
rect 27476 -22322 27516 -22242
rect 27596 -22322 27636 -22242
rect 27716 -22322 27756 -22242
rect 27836 -22322 27876 -22242
rect 27956 -22322 27996 -22242
rect 28076 -22322 28116 -22242
rect 28196 -22322 28236 -22242
rect 28316 -22322 28356 -22242
rect 28436 -22322 28476 -22242
rect 28556 -22322 28596 -22242
rect 28676 -22322 28716 -22242
rect 28796 -22322 28836 -22242
rect 28916 -22322 28956 -22242
rect 29036 -22322 29076 -22242
rect 29156 -22322 29176 -22242
rect 30404 -22269 30646 -22263
rect 30404 -22282 30416 -22269
rect 24616 -22342 29176 -22322
rect 30396 -22303 30416 -22282
rect 30634 -22282 30646 -22269
rect 30712 -22269 30954 -22263
rect 30712 -22282 30724 -22269
rect 30634 -22303 30724 -22282
rect 30942 -22282 30954 -22269
rect 31020 -22269 31262 -22263
rect 31020 -22282 31032 -22269
rect 30942 -22303 31032 -22282
rect 31250 -22282 31262 -22269
rect 31328 -22269 31570 -22263
rect 31328 -22282 31340 -22269
rect 31250 -22303 31340 -22282
rect 31558 -22282 31570 -22269
rect 31636 -22269 31878 -22263
rect 31636 -22282 31648 -22269
rect 31558 -22303 31648 -22282
rect 31866 -22282 31878 -22269
rect 31944 -22269 32186 -22263
rect 31944 -22282 31956 -22269
rect 31866 -22303 31956 -22282
rect 32174 -22282 32186 -22269
rect 32252 -22269 32494 -22263
rect 32252 -22282 32264 -22269
rect 32174 -22303 32264 -22282
rect 32482 -22282 32494 -22269
rect 32560 -22269 32802 -22263
rect 32560 -22282 32572 -22269
rect 32482 -22303 32572 -22282
rect 32790 -22282 32802 -22269
rect 32790 -22303 32816 -22282
rect 20956 -22522 20976 -22442
rect 21056 -22522 21076 -22442
rect 21156 -22522 21176 -22442
rect 21256 -22522 21276 -22442
rect 21356 -22522 21376 -22442
rect 21456 -22522 21476 -22442
rect 21556 -22522 21576 -22442
rect 21656 -22522 21676 -22442
rect 21756 -22522 21776 -22442
rect 21856 -22522 21876 -22442
rect 21956 -22522 21976 -22442
rect 22056 -22522 22076 -22442
rect 22156 -22522 22176 -22442
rect 22256 -22522 22276 -22442
rect 22356 -22522 22376 -22442
rect 22456 -22522 22476 -22442
rect 22556 -22522 22576 -22442
rect 22656 -22522 22676 -22442
rect 22756 -22522 22776 -22442
rect 22856 -22522 22876 -22442
rect 22956 -22522 22976 -22442
rect 23056 -22522 23076 -22442
rect 23156 -22522 23176 -22442
rect 23256 -22522 23276 -22442
rect 23356 -22522 23376 -22442
rect 20956 -22582 23376 -22522
rect 20956 -22662 20976 -22582
rect 21056 -22662 21076 -22582
rect 21156 -22662 21176 -22582
rect 21256 -22662 21276 -22582
rect 21356 -22662 21376 -22582
rect 21456 -22662 21476 -22582
rect 21556 -22662 21576 -22582
rect 21656 -22662 21676 -22582
rect 21756 -22662 21776 -22582
rect 21856 -22662 21876 -22582
rect 21956 -22662 21976 -22582
rect 22056 -22662 22076 -22582
rect 22156 -22662 22176 -22582
rect 22256 -22662 22276 -22582
rect 22356 -22662 22376 -22582
rect 22456 -22662 22476 -22582
rect 22556 -22662 22576 -22582
rect 22656 -22662 22676 -22582
rect 22756 -22662 22776 -22582
rect 22856 -22662 22876 -22582
rect 22956 -22662 22976 -22582
rect 23056 -22662 23076 -22582
rect 23156 -22662 23176 -22582
rect 23256 -22662 23276 -22582
rect 23356 -22662 23376 -22582
rect 20956 -22722 23376 -22662
rect 20956 -22802 20976 -22722
rect 21056 -22802 21076 -22722
rect 21156 -22802 21176 -22722
rect 21256 -22802 21276 -22722
rect 21356 -22802 21376 -22722
rect 21456 -22802 21476 -22722
rect 21556 -22802 21576 -22722
rect 21656 -22802 21676 -22722
rect 21756 -22802 21776 -22722
rect 21856 -22802 21876 -22722
rect 21956 -22802 21976 -22722
rect 22056 -22802 22076 -22722
rect 22156 -22802 22176 -22722
rect 22256 -22802 22276 -22722
rect 22356 -22802 22376 -22722
rect 22456 -22802 22476 -22722
rect 22556 -22802 22576 -22722
rect 22656 -22802 22676 -22722
rect 22756 -22802 22776 -22722
rect 22856 -22802 22876 -22722
rect 22956 -22802 22976 -22722
rect 23056 -22802 23076 -22722
rect 23156 -22802 23176 -22722
rect 23256 -22802 23276 -22722
rect 23356 -22802 23376 -22722
rect 20956 -22822 23376 -22802
rect 30396 -22442 32816 -22303
rect 30396 -22522 30416 -22442
rect 30496 -22522 30516 -22442
rect 30596 -22522 30616 -22442
rect 30696 -22522 30716 -22442
rect 30796 -22522 30816 -22442
rect 30896 -22522 30916 -22442
rect 30996 -22522 31016 -22442
rect 31096 -22522 31116 -22442
rect 31196 -22522 31216 -22442
rect 31296 -22522 31316 -22442
rect 31396 -22522 31416 -22442
rect 31496 -22522 31516 -22442
rect 31596 -22522 31616 -22442
rect 31696 -22522 31716 -22442
rect 31796 -22522 31816 -22442
rect 31896 -22522 31916 -22442
rect 31996 -22522 32016 -22442
rect 32096 -22522 32116 -22442
rect 32196 -22522 32216 -22442
rect 32296 -22522 32316 -22442
rect 32396 -22522 32416 -22442
rect 32496 -22522 32516 -22442
rect 32596 -22522 32616 -22442
rect 32696 -22522 32716 -22442
rect 32796 -22522 32816 -22442
rect 30396 -22582 32816 -22522
rect 30396 -22662 30416 -22582
rect 30496 -22662 30516 -22582
rect 30596 -22662 30616 -22582
rect 30696 -22662 30716 -22582
rect 30796 -22662 30816 -22582
rect 30896 -22662 30916 -22582
rect 30996 -22662 31016 -22582
rect 31096 -22662 31116 -22582
rect 31196 -22662 31216 -22582
rect 31296 -22662 31316 -22582
rect 31396 -22662 31416 -22582
rect 31496 -22662 31516 -22582
rect 31596 -22662 31616 -22582
rect 31696 -22662 31716 -22582
rect 31796 -22662 31816 -22582
rect 31896 -22662 31916 -22582
rect 31996 -22662 32016 -22582
rect 32096 -22662 32116 -22582
rect 32196 -22662 32216 -22582
rect 32296 -22662 32316 -22582
rect 32396 -22662 32416 -22582
rect 32496 -22662 32516 -22582
rect 32596 -22662 32616 -22582
rect 32696 -22662 32716 -22582
rect 32796 -22662 32816 -22582
rect 30396 -22722 32816 -22662
rect 30396 -22802 30416 -22722
rect 30496 -22802 30516 -22722
rect 30596 -22802 30616 -22722
rect 30696 -22802 30716 -22722
rect 30796 -22802 30816 -22722
rect 30896 -22802 30916 -22722
rect 30996 -22802 31016 -22722
rect 31096 -22802 31116 -22722
rect 31196 -22802 31216 -22722
rect 31296 -22802 31316 -22722
rect 31396 -22802 31416 -22722
rect 31496 -22802 31516 -22722
rect 31596 -22802 31616 -22722
rect 31696 -22802 31716 -22722
rect 31796 -22802 31816 -22722
rect 31896 -22802 31916 -22722
rect 31996 -22802 32016 -22722
rect 32096 -22802 32116 -22722
rect 32196 -22802 32216 -22722
rect 32296 -22802 32316 -22722
rect 32396 -22802 32416 -22722
rect 32496 -22802 32516 -22722
rect 32596 -22802 32616 -22722
rect 32696 -22802 32716 -22722
rect 32796 -22802 32816 -22722
rect 30396 -22822 32816 -22802
rect 26696 -22922 27096 -22902
rect 21868 -22934 21914 -22922
rect 21868 -22962 21874 -22934
rect 21816 -22982 21874 -22962
rect 21908 -22962 21914 -22934
rect 22106 -22934 22152 -22922
rect 21908 -22982 21956 -22962
rect 21816 -23042 21856 -22982
rect 21916 -23042 21956 -22982
rect 21816 -23162 21874 -23042
rect 21908 -23162 21956 -23042
rect 21816 -23222 21856 -23162
rect 21916 -23222 21956 -23162
rect 21816 -23242 21874 -23222
rect 21868 -23910 21874 -23242
rect 21908 -23242 21956 -23222
rect 21908 -23910 21914 -23242
rect 22106 -23442 22112 -22934
rect 22056 -23642 22112 -23442
rect 22146 -23442 22152 -22934
rect 22344 -22934 22390 -22922
rect 22344 -22962 22350 -22934
rect 22276 -22982 22350 -22962
rect 22384 -22962 22390 -22934
rect 22276 -23042 22316 -22982
rect 22276 -23162 22350 -23042
rect 22276 -23222 22316 -23162
rect 22276 -23242 22350 -23222
rect 22146 -23462 22196 -23442
rect 22176 -23522 22196 -23462
rect 22146 -23562 22196 -23522
rect 22176 -23622 22196 -23562
rect 21868 -23922 21914 -23910
rect 22106 -23910 22112 -23642
rect 22146 -23642 22196 -23622
rect 22146 -23910 22152 -23642
rect 22106 -23922 22152 -23910
rect 22344 -23910 22350 -23242
rect 22384 -23242 22416 -22962
rect 26696 -23002 26716 -22922
rect 26796 -23002 26856 -22922
rect 26936 -23002 26996 -22922
rect 27076 -23002 27096 -22922
rect 31448 -22914 31494 -22902
rect 31448 -22962 31454 -22914
rect 23916 -23082 25856 -23002
rect 23916 -23102 24856 -23082
rect 23362 -23156 23408 -23144
rect 22384 -23910 22390 -23242
rect 22344 -23922 22390 -23910
rect 21924 -23969 22096 -23963
rect 21924 -23982 21936 -23969
rect 21916 -24003 21936 -23982
rect 22084 -23982 22096 -23969
rect 22162 -23969 22334 -23963
rect 22162 -23982 22174 -23969
rect 22084 -24003 22174 -23982
rect 22322 -23982 22334 -23969
rect 22322 -24003 22336 -23982
rect 21916 -24402 22336 -24003
rect 23362 -24082 23368 -23156
rect 23402 -24082 23408 -23156
rect 23362 -24094 23408 -24082
rect 23520 -23156 23566 -23144
rect 23520 -24082 23526 -23156
rect 23560 -24082 23566 -23156
rect 23520 -24094 23566 -24082
rect 23678 -23156 23724 -23144
rect 23678 -24082 23684 -23156
rect 23718 -24082 23724 -23156
rect 23802 -23156 23848 -23144
rect 23802 -23442 23808 -23156
rect 23776 -23462 23808 -23442
rect 23842 -23442 23848 -23156
rect 23916 -23156 24056 -23102
rect 23842 -23462 23876 -23442
rect 23776 -23522 23796 -23462
rect 23856 -23522 23876 -23462
rect 23776 -23542 23808 -23522
rect 23842 -23542 23876 -23522
rect 23776 -23602 23796 -23542
rect 23856 -23602 23876 -23542
rect 23776 -23622 23808 -23602
rect 23842 -23622 23876 -23602
rect 23776 -23682 23796 -23622
rect 23856 -23682 23876 -23622
rect 23776 -23702 23808 -23682
rect 23678 -24094 23724 -24082
rect 23802 -24082 23808 -23702
rect 23842 -23702 23876 -23682
rect 23842 -24082 23848 -23702
rect 23916 -24082 23966 -23156
rect 24000 -24082 24056 -23156
rect 24118 -23156 24164 -23144
rect 24118 -23442 24124 -23156
rect 24096 -23462 24124 -23442
rect 24158 -23442 24164 -23156
rect 24242 -23156 24288 -23144
rect 24158 -23462 24196 -23442
rect 24096 -23522 24116 -23462
rect 24176 -23522 24196 -23462
rect 24096 -23542 24124 -23522
rect 24158 -23542 24196 -23522
rect 24096 -23602 24116 -23542
rect 24176 -23602 24196 -23542
rect 24096 -23622 24124 -23602
rect 24158 -23622 24196 -23602
rect 24096 -23682 24116 -23622
rect 24176 -23682 24196 -23622
rect 24096 -23702 24124 -23682
rect 24118 -24082 24124 -23702
rect 24158 -23702 24196 -23682
rect 24158 -24082 24164 -23702
rect 23802 -24094 23848 -24082
rect 23960 -24094 24006 -24082
rect 24118 -24094 24164 -24082
rect 24242 -24082 24248 -23156
rect 24282 -24082 24288 -23156
rect 24242 -24094 24288 -24082
rect 24400 -23156 24446 -23144
rect 24400 -24082 24406 -23156
rect 24440 -24082 24446 -23156
rect 24400 -24094 24446 -24082
rect 24558 -23156 24604 -23144
rect 24558 -24082 24564 -23156
rect 24598 -24082 24604 -23156
rect 24558 -24094 24604 -24082
rect 24816 -23162 24856 -23102
rect 24936 -23102 25856 -23082
rect 24936 -23162 24976 -23102
rect 24816 -23202 24976 -23162
rect 24816 -23282 24856 -23202
rect 24936 -23282 24976 -23202
rect 24816 -23322 24976 -23282
rect 24816 -23402 24856 -23322
rect 24936 -23402 24976 -23322
rect 24816 -23442 24976 -23402
rect 24816 -23522 24856 -23442
rect 24936 -23522 24976 -23442
rect 24816 -23562 24976 -23522
rect 24816 -23642 24856 -23562
rect 24936 -23642 24976 -23562
rect 24816 -23682 24976 -23642
rect 24816 -23762 24856 -23682
rect 24936 -23762 24976 -23682
rect 24816 -23802 24976 -23762
rect 24816 -23882 24856 -23802
rect 24936 -23882 24976 -23802
rect 24816 -23922 24976 -23882
rect 24816 -24002 24856 -23922
rect 24936 -24002 24976 -23922
rect 24816 -24042 24976 -24002
rect 24816 -24122 24856 -24042
rect 24936 -24122 24976 -24042
rect 25162 -23156 25208 -23144
rect 25162 -24082 25168 -23156
rect 25202 -24082 25208 -23156
rect 25162 -24094 25208 -24082
rect 25320 -23156 25366 -23144
rect 25320 -24082 25326 -23156
rect 25360 -24082 25366 -23156
rect 25320 -24094 25366 -24082
rect 25478 -23156 25524 -23144
rect 25478 -24082 25484 -23156
rect 25518 -24082 25524 -23156
rect 25602 -23156 25648 -23144
rect 25602 -23442 25608 -23156
rect 25576 -23462 25608 -23442
rect 25642 -23442 25648 -23156
rect 25716 -23156 25856 -23102
rect 26696 -23042 27096 -23002
rect 26696 -23122 26716 -23042
rect 26796 -23122 26856 -23042
rect 26936 -23122 26996 -23042
rect 27076 -23122 27096 -23042
rect 25642 -23462 25676 -23442
rect 25576 -23522 25596 -23462
rect 25656 -23522 25676 -23462
rect 25576 -23542 25608 -23522
rect 25642 -23542 25676 -23522
rect 25576 -23602 25596 -23542
rect 25656 -23602 25676 -23542
rect 25576 -23622 25608 -23602
rect 25642 -23622 25676 -23602
rect 25576 -23682 25596 -23622
rect 25656 -23682 25676 -23622
rect 25576 -23702 25608 -23682
rect 25478 -24094 25524 -24082
rect 25602 -24082 25608 -23702
rect 25642 -23702 25676 -23682
rect 25642 -24082 25648 -23702
rect 25716 -24082 25766 -23156
rect 25800 -24082 25856 -23156
rect 25918 -23156 25964 -23144
rect 25918 -23442 25924 -23156
rect 25896 -23462 25924 -23442
rect 25958 -23442 25964 -23156
rect 26042 -23156 26088 -23144
rect 25958 -23462 25996 -23442
rect 25896 -23522 25916 -23462
rect 25976 -23522 25996 -23462
rect 25896 -23542 25924 -23522
rect 25958 -23542 25996 -23522
rect 25896 -23602 25916 -23542
rect 25976 -23602 25996 -23542
rect 25896 -23622 25924 -23602
rect 25958 -23622 25996 -23602
rect 25896 -23682 25916 -23622
rect 25976 -23682 25996 -23622
rect 25896 -23702 25924 -23682
rect 25918 -24082 25924 -23702
rect 25958 -23702 25996 -23682
rect 25958 -24082 25964 -23702
rect 25602 -24094 25648 -24082
rect 25760 -24094 25806 -24082
rect 25918 -24094 25964 -24082
rect 26042 -24082 26048 -23156
rect 26082 -24082 26088 -23156
rect 26042 -24094 26088 -24082
rect 26200 -23156 26246 -23144
rect 26200 -24082 26206 -23156
rect 26240 -24082 26246 -23156
rect 26200 -24094 26246 -24082
rect 26358 -23156 26404 -23144
rect 26358 -24082 26364 -23156
rect 26398 -24082 26404 -23156
rect 26358 -24094 26404 -24082
rect 26696 -23162 27096 -23122
rect 27916 -23082 29856 -23002
rect 27916 -23102 28856 -23082
rect 26696 -23242 26716 -23162
rect 26796 -23242 26856 -23162
rect 26936 -23242 26996 -23162
rect 27076 -23242 27096 -23162
rect 26696 -23282 27096 -23242
rect 26696 -23362 26716 -23282
rect 26796 -23362 26856 -23282
rect 26936 -23362 26996 -23282
rect 27076 -23362 27096 -23282
rect 26696 -23402 27096 -23362
rect 26696 -23482 26716 -23402
rect 26796 -23482 26856 -23402
rect 26936 -23482 26996 -23402
rect 27076 -23482 27096 -23402
rect 26696 -23522 27096 -23482
rect 26696 -23602 26716 -23522
rect 26796 -23602 26856 -23522
rect 26936 -23602 26996 -23522
rect 27076 -23602 27096 -23522
rect 26696 -23642 27096 -23602
rect 26696 -23722 26716 -23642
rect 26796 -23722 26856 -23642
rect 26936 -23722 26996 -23642
rect 27076 -23722 27096 -23642
rect 26696 -23762 27096 -23722
rect 26696 -23842 26716 -23762
rect 26796 -23842 26856 -23762
rect 26936 -23842 26996 -23762
rect 27076 -23842 27096 -23762
rect 26696 -23882 27096 -23842
rect 26696 -23962 26716 -23882
rect 26796 -23962 26856 -23882
rect 26936 -23962 26996 -23882
rect 27076 -23962 27096 -23882
rect 26696 -24002 27096 -23962
rect 26696 -24082 26716 -24002
rect 26796 -24082 26856 -24002
rect 26936 -24082 26996 -24002
rect 27076 -24082 27096 -24002
rect 26696 -24122 27096 -24082
rect 27362 -23156 27408 -23144
rect 27362 -24082 27368 -23156
rect 27402 -24082 27408 -23156
rect 27362 -24094 27408 -24082
rect 27520 -23156 27566 -23144
rect 27520 -24082 27526 -23156
rect 27560 -24082 27566 -23156
rect 27520 -24094 27566 -24082
rect 27678 -23156 27724 -23144
rect 27678 -24082 27684 -23156
rect 27718 -24082 27724 -23156
rect 27802 -23156 27848 -23144
rect 27802 -23442 27808 -23156
rect 27776 -23462 27808 -23442
rect 27842 -23442 27848 -23156
rect 27916 -23156 28056 -23102
rect 27842 -23462 27876 -23442
rect 27776 -23522 27796 -23462
rect 27856 -23522 27876 -23462
rect 27776 -23542 27808 -23522
rect 27842 -23542 27876 -23522
rect 27776 -23602 27796 -23542
rect 27856 -23602 27876 -23542
rect 27776 -23622 27808 -23602
rect 27842 -23622 27876 -23602
rect 27776 -23682 27796 -23622
rect 27856 -23682 27876 -23622
rect 27776 -23702 27808 -23682
rect 27678 -24094 27724 -24082
rect 27802 -24082 27808 -23702
rect 27842 -23702 27876 -23682
rect 27842 -24082 27848 -23702
rect 27916 -24082 27966 -23156
rect 28000 -24082 28056 -23156
rect 28118 -23156 28164 -23144
rect 28118 -23442 28124 -23156
rect 28096 -23462 28124 -23442
rect 28158 -23442 28164 -23156
rect 28242 -23156 28288 -23144
rect 28158 -23462 28196 -23442
rect 28096 -23522 28116 -23462
rect 28176 -23522 28196 -23462
rect 28096 -23542 28124 -23522
rect 28158 -23542 28196 -23522
rect 28096 -23602 28116 -23542
rect 28176 -23602 28196 -23542
rect 28096 -23622 28124 -23602
rect 28158 -23622 28196 -23602
rect 28096 -23682 28116 -23622
rect 28176 -23682 28196 -23622
rect 28096 -23702 28124 -23682
rect 28118 -24082 28124 -23702
rect 28158 -23702 28196 -23682
rect 28158 -24082 28164 -23702
rect 27802 -24094 27848 -24082
rect 27960 -24094 28006 -24082
rect 28118 -24094 28164 -24082
rect 28242 -24082 28248 -23156
rect 28282 -24082 28288 -23156
rect 28242 -24094 28288 -24082
rect 28400 -23156 28446 -23144
rect 28400 -24082 28406 -23156
rect 28440 -24082 28446 -23156
rect 28400 -24094 28446 -24082
rect 28558 -23156 28604 -23144
rect 28558 -24082 28564 -23156
rect 28598 -24082 28604 -23156
rect 28558 -24094 28604 -24082
rect 28816 -23162 28856 -23102
rect 28936 -23102 29856 -23082
rect 28936 -23162 28976 -23102
rect 28816 -23202 28976 -23162
rect 28816 -23282 28856 -23202
rect 28936 -23282 28976 -23202
rect 28816 -23322 28976 -23282
rect 28816 -23402 28856 -23322
rect 28936 -23402 28976 -23322
rect 28816 -23442 28976 -23402
rect 28816 -23522 28856 -23442
rect 28936 -23522 28976 -23442
rect 28816 -23562 28976 -23522
rect 28816 -23642 28856 -23562
rect 28936 -23642 28976 -23562
rect 28816 -23682 28976 -23642
rect 28816 -23762 28856 -23682
rect 28936 -23762 28976 -23682
rect 28816 -23802 28976 -23762
rect 28816 -23882 28856 -23802
rect 28936 -23882 28976 -23802
rect 28816 -23922 28976 -23882
rect 28816 -24002 28856 -23922
rect 28936 -24002 28976 -23922
rect 28816 -24042 28976 -24002
rect 28816 -24122 28856 -24042
rect 28936 -24122 28976 -24042
rect 29162 -23156 29208 -23144
rect 29162 -24082 29168 -23156
rect 29202 -24082 29208 -23156
rect 29162 -24094 29208 -24082
rect 29320 -23156 29366 -23144
rect 29320 -24082 29326 -23156
rect 29360 -24082 29366 -23156
rect 29320 -24094 29366 -24082
rect 29478 -23156 29524 -23144
rect 29478 -24082 29484 -23156
rect 29518 -24082 29524 -23156
rect 29602 -23156 29648 -23144
rect 29602 -23442 29608 -23156
rect 29576 -23462 29608 -23442
rect 29642 -23442 29648 -23156
rect 29716 -23156 29856 -23102
rect 29642 -23462 29676 -23442
rect 29576 -23522 29596 -23462
rect 29656 -23522 29676 -23462
rect 29576 -23542 29608 -23522
rect 29642 -23542 29676 -23522
rect 29576 -23602 29596 -23542
rect 29656 -23602 29676 -23542
rect 29576 -23622 29608 -23602
rect 29642 -23622 29676 -23602
rect 29576 -23682 29596 -23622
rect 29656 -23682 29676 -23622
rect 29576 -23702 29608 -23682
rect 29478 -24094 29524 -24082
rect 29602 -24082 29608 -23702
rect 29642 -23702 29676 -23682
rect 29642 -24082 29648 -23702
rect 29716 -24082 29766 -23156
rect 29800 -24082 29856 -23156
rect 29918 -23156 29964 -23144
rect 29918 -23442 29924 -23156
rect 29896 -23462 29924 -23442
rect 29958 -23442 29964 -23156
rect 30042 -23156 30088 -23144
rect 29958 -23462 29996 -23442
rect 29896 -23522 29916 -23462
rect 29976 -23522 29996 -23462
rect 29896 -23542 29924 -23522
rect 29958 -23542 29996 -23522
rect 29896 -23602 29916 -23542
rect 29976 -23602 29996 -23542
rect 29896 -23622 29924 -23602
rect 29958 -23622 29996 -23602
rect 29896 -23682 29916 -23622
rect 29976 -23682 29996 -23622
rect 29896 -23702 29924 -23682
rect 29918 -24082 29924 -23702
rect 29958 -23702 29996 -23682
rect 29958 -24082 29964 -23702
rect 29602 -24094 29648 -24082
rect 29760 -24094 29806 -24082
rect 29918 -24094 29964 -24082
rect 30042 -24082 30048 -23156
rect 30082 -24082 30088 -23156
rect 30042 -24094 30088 -24082
rect 30200 -23156 30246 -23144
rect 30200 -24082 30206 -23156
rect 30240 -24082 30246 -23156
rect 30200 -24094 30246 -24082
rect 30358 -23156 30404 -23144
rect 30358 -24082 30364 -23156
rect 30398 -24082 30404 -23156
rect 31436 -23242 31454 -22962
rect 31488 -22962 31494 -22914
rect 31686 -22914 31732 -22902
rect 31488 -22982 31576 -22962
rect 31516 -23042 31576 -22982
rect 31488 -23162 31576 -23042
rect 31516 -23222 31576 -23162
rect 31448 -23890 31454 -23242
rect 31488 -23242 31576 -23222
rect 31488 -23890 31494 -23242
rect 31686 -23442 31692 -22914
rect 31616 -23462 31692 -23442
rect 31726 -23442 31732 -22914
rect 31924 -22914 31970 -22902
rect 31924 -22962 31930 -22914
rect 31876 -22982 31930 -22962
rect 31964 -22962 31970 -22914
rect 31964 -22982 32016 -22962
rect 31876 -23042 31916 -22982
rect 31976 -23042 32016 -22982
rect 31876 -23162 31930 -23042
rect 31964 -23162 32016 -23042
rect 31876 -23222 31916 -23162
rect 31976 -23222 32016 -23162
rect 31876 -23242 31930 -23222
rect 31616 -23522 31636 -23462
rect 31616 -23562 31692 -23522
rect 31616 -23622 31636 -23562
rect 31616 -23642 31692 -23622
rect 31448 -23902 31494 -23890
rect 31686 -23890 31692 -23642
rect 31726 -23642 31756 -23442
rect 31726 -23890 31732 -23642
rect 31686 -23902 31732 -23890
rect 31924 -23890 31930 -23242
rect 31964 -23242 32016 -23222
rect 31964 -23890 31970 -23242
rect 31924 -23902 31970 -23890
rect 31504 -23949 31676 -23943
rect 31504 -23982 31516 -23949
rect 30358 -24094 30404 -24082
rect 31496 -23983 31516 -23982
rect 31664 -23982 31676 -23949
rect 31742 -23949 31914 -23943
rect 31742 -23982 31754 -23949
rect 31664 -23983 31754 -23982
rect 31902 -23982 31914 -23949
rect 31902 -23983 31916 -23982
rect 23418 -24132 23510 -24126
rect 23418 -24166 23430 -24132
rect 23498 -24166 23510 -24132
rect 23418 -24172 23510 -24166
rect 23576 -24132 23668 -24126
rect 23576 -24166 23588 -24132
rect 23656 -24166 23668 -24132
rect 23576 -24172 23668 -24166
rect 23856 -24132 24116 -24122
rect 23856 -24166 23870 -24132
rect 23938 -24166 24028 -24132
rect 23856 -24202 23876 -24166
rect 23936 -24202 24036 -24166
rect 24096 -24202 24116 -24132
rect 24298 -24132 24390 -24126
rect 24298 -24166 24310 -24132
rect 24378 -24166 24390 -24132
rect 24298 -24172 24390 -24166
rect 24456 -24132 24548 -24126
rect 24456 -24166 24468 -24132
rect 24536 -24166 24548 -24132
rect 24456 -24172 24548 -24166
rect 24816 -24162 24976 -24122
rect 23856 -24262 24116 -24202
rect 24816 -24242 24856 -24162
rect 24936 -24242 24976 -24162
rect 25218 -24132 25310 -24126
rect 25218 -24166 25230 -24132
rect 25298 -24166 25310 -24132
rect 25218 -24172 25310 -24166
rect 25376 -24132 25468 -24126
rect 25376 -24166 25388 -24132
rect 25456 -24166 25468 -24132
rect 25376 -24172 25468 -24166
rect 25656 -24132 25916 -24122
rect 25656 -24166 25670 -24132
rect 25738 -24166 25828 -24132
rect 24816 -24282 24976 -24242
rect 25656 -24202 25676 -24166
rect 25736 -24202 25836 -24166
rect 25896 -24202 25916 -24132
rect 26098 -24132 26190 -24126
rect 26098 -24166 26110 -24132
rect 26178 -24166 26190 -24132
rect 26098 -24172 26190 -24166
rect 26256 -24132 26348 -24126
rect 26256 -24166 26268 -24132
rect 26336 -24166 26348 -24132
rect 26256 -24172 26348 -24166
rect 25656 -24262 25916 -24202
rect 26696 -24202 26716 -24122
rect 26796 -24202 26856 -24122
rect 26936 -24202 26996 -24122
rect 27076 -24202 27096 -24122
rect 27418 -24132 27510 -24126
rect 27418 -24166 27430 -24132
rect 27498 -24166 27510 -24132
rect 27418 -24172 27510 -24166
rect 27576 -24132 27668 -24126
rect 27576 -24166 27588 -24132
rect 27656 -24166 27668 -24132
rect 27576 -24172 27668 -24166
rect 27856 -24132 28116 -24122
rect 27856 -24166 27870 -24132
rect 27938 -24166 28028 -24132
rect 26696 -24242 27096 -24202
rect 24816 -24342 24856 -24282
rect 21916 -24482 21936 -24402
rect 22016 -24482 22076 -24402
rect 22176 -24482 22236 -24402
rect 22316 -24482 22336 -24402
rect 21916 -24522 22336 -24482
rect 23216 -24362 24856 -24342
rect 24936 -24342 24976 -24282
rect 26696 -24322 26716 -24242
rect 26796 -24322 26856 -24242
rect 26936 -24322 26996 -24242
rect 27076 -24322 27096 -24242
rect 27856 -24202 27876 -24166
rect 27936 -24202 28036 -24166
rect 28096 -24202 28116 -24132
rect 28298 -24132 28390 -24126
rect 28298 -24166 28310 -24132
rect 28378 -24166 28390 -24132
rect 28298 -24172 28390 -24166
rect 28456 -24132 28548 -24126
rect 28456 -24166 28468 -24132
rect 28536 -24166 28548 -24132
rect 28456 -24172 28548 -24166
rect 28816 -24162 28976 -24122
rect 27856 -24262 28116 -24202
rect 28816 -24242 28856 -24162
rect 28936 -24242 28976 -24162
rect 29218 -24132 29310 -24126
rect 29218 -24166 29230 -24132
rect 29298 -24166 29310 -24132
rect 29218 -24172 29310 -24166
rect 29376 -24132 29468 -24126
rect 29658 -24132 29750 -24126
rect 29816 -24132 29908 -24126
rect 30098 -24132 30190 -24126
rect 29376 -24166 29388 -24132
rect 29456 -24166 29468 -24132
rect 29376 -24172 29468 -24166
rect 29656 -24166 29670 -24132
rect 29738 -24166 29828 -24132
rect 26696 -24342 27096 -24322
rect 28816 -24282 28976 -24242
rect 29656 -24202 29676 -24166
rect 29736 -24202 29836 -24166
rect 29896 -24202 29916 -24132
rect 30098 -24166 30110 -24132
rect 30178 -24166 30190 -24132
rect 30098 -24172 30190 -24166
rect 30256 -24132 30348 -24126
rect 30256 -24166 30268 -24132
rect 30336 -24166 30348 -24132
rect 30256 -24172 30348 -24166
rect 29656 -24272 29916 -24202
rect 28816 -24342 28856 -24282
rect 24936 -24362 28856 -24342
rect 28936 -24342 28976 -24282
rect 28936 -24362 30576 -24342
rect 23216 -24442 23236 -24362
rect 23316 -24442 23356 -24362
rect 23436 -24442 23476 -24362
rect 23556 -24442 23596 -24362
rect 23676 -24442 23716 -24362
rect 23796 -24442 23836 -24362
rect 23916 -24442 23956 -24362
rect 24036 -24442 24076 -24362
rect 24156 -24442 24196 -24362
rect 24276 -24442 24316 -24362
rect 24396 -24442 24436 -24362
rect 24516 -24442 24556 -24362
rect 24636 -24442 24676 -24362
rect 24756 -24402 25036 -24362
rect 24756 -24442 24856 -24402
rect 23216 -24482 24856 -24442
rect 24936 -24442 25036 -24402
rect 25116 -24442 25156 -24362
rect 25236 -24442 25276 -24362
rect 25356 -24442 25396 -24362
rect 25476 -24442 25516 -24362
rect 25596 -24442 25636 -24362
rect 25716 -24442 25756 -24362
rect 25836 -24442 25876 -24362
rect 25956 -24442 25996 -24362
rect 26076 -24442 26116 -24362
rect 26196 -24442 26236 -24362
rect 26316 -24442 26356 -24362
rect 26436 -24442 26476 -24362
rect 26556 -24442 26596 -24362
rect 26676 -24442 26716 -24362
rect 26796 -24442 26856 -24362
rect 26936 -24442 26996 -24362
rect 27076 -24442 27116 -24362
rect 27196 -24442 27236 -24362
rect 27316 -24442 27356 -24362
rect 27436 -24442 27476 -24362
rect 27556 -24442 27596 -24362
rect 27676 -24442 27716 -24362
rect 27796 -24442 27836 -24362
rect 27916 -24442 27956 -24362
rect 28036 -24442 28076 -24362
rect 28156 -24442 28196 -24362
rect 28276 -24442 28316 -24362
rect 28396 -24442 28436 -24362
rect 28516 -24442 28556 -24362
rect 28636 -24442 28676 -24362
rect 28756 -24402 29036 -24362
rect 28756 -24442 28856 -24402
rect 24936 -24482 28856 -24442
rect 28936 -24442 29036 -24402
rect 29116 -24442 29156 -24362
rect 29236 -24442 29276 -24362
rect 29356 -24442 29396 -24362
rect 29476 -24442 29516 -24362
rect 29596 -24442 29636 -24362
rect 29716 -24442 29756 -24362
rect 29836 -24442 29876 -24362
rect 29956 -24442 29996 -24362
rect 30076 -24442 30116 -24362
rect 30196 -24442 30236 -24362
rect 30316 -24442 30356 -24362
rect 30436 -24442 30476 -24362
rect 30556 -24442 30576 -24362
rect 28936 -24482 30576 -24442
rect 23216 -24502 26716 -24482
rect 23216 -24582 23236 -24502
rect 23316 -24582 23356 -24502
rect 23436 -24582 23476 -24502
rect 23556 -24582 23596 -24502
rect 23676 -24582 23716 -24502
rect 23796 -24582 23836 -24502
rect 23916 -24582 23956 -24502
rect 24036 -24582 24076 -24502
rect 24156 -24582 24196 -24502
rect 24276 -24582 24316 -24502
rect 24396 -24582 24436 -24502
rect 24516 -24582 24556 -24502
rect 24636 -24582 24676 -24502
rect 24756 -24522 25036 -24502
rect 24756 -24582 24856 -24522
rect 23216 -24602 24856 -24582
rect 24936 -24582 25036 -24522
rect 25116 -24582 25156 -24502
rect 25236 -24582 25276 -24502
rect 25356 -24582 25396 -24502
rect 25476 -24582 25516 -24502
rect 25596 -24582 25636 -24502
rect 25716 -24582 25756 -24502
rect 25836 -24582 25876 -24502
rect 25956 -24582 25996 -24502
rect 26076 -24582 26116 -24502
rect 26196 -24582 26236 -24502
rect 26316 -24582 26356 -24502
rect 26436 -24582 26476 -24502
rect 26556 -24582 26596 -24502
rect 26676 -24562 26716 -24502
rect 26796 -24562 26856 -24482
rect 26936 -24562 26996 -24482
rect 27076 -24502 30576 -24482
rect 27076 -24562 27116 -24502
rect 26676 -24582 27116 -24562
rect 27196 -24582 27236 -24502
rect 27316 -24582 27356 -24502
rect 27436 -24582 27476 -24502
rect 27556 -24582 27596 -24502
rect 27676 -24582 27716 -24502
rect 27796 -24582 27836 -24502
rect 27916 -24582 27956 -24502
rect 28036 -24582 28076 -24502
rect 28156 -24582 28196 -24502
rect 28276 -24582 28316 -24502
rect 28396 -24582 28436 -24502
rect 28516 -24582 28556 -24502
rect 28636 -24582 28676 -24502
rect 28756 -24522 29036 -24502
rect 28756 -24582 28856 -24522
rect 24936 -24602 28856 -24582
rect 28936 -24582 29036 -24522
rect 29116 -24582 29156 -24502
rect 29236 -24582 29276 -24502
rect 29356 -24582 29396 -24502
rect 29476 -24582 29516 -24502
rect 29596 -24582 29636 -24502
rect 29716 -24582 29756 -24502
rect 29836 -24582 29876 -24502
rect 29956 -24582 29996 -24502
rect 30076 -24582 30116 -24502
rect 30196 -24582 30236 -24502
rect 30316 -24582 30356 -24502
rect 30436 -24582 30476 -24502
rect 30556 -24582 30576 -24502
rect 31496 -24402 31916 -23983
rect 31496 -24482 31516 -24402
rect 31596 -24482 31636 -24402
rect 31776 -24482 31816 -24402
rect 31896 -24482 31916 -24402
rect 31496 -24522 31916 -24482
rect 28936 -24602 30576 -24582
rect 24816 -24642 24976 -24602
rect 23856 -24742 24116 -24672
rect 21422 -24766 21468 -24754
rect 21422 -24962 21428 -24766
rect 21356 -24982 21428 -24962
rect 21462 -24962 21468 -24766
rect 21730 -24766 21776 -24754
rect 21462 -24982 21536 -24962
rect 21356 -25042 21416 -24982
rect 21476 -25042 21536 -24982
rect 21356 -25162 21428 -25042
rect 21462 -25162 21536 -25042
rect 21356 -25222 21416 -25162
rect 21476 -25222 21536 -25162
rect 21356 -25242 21428 -25222
rect 21422 -26242 21428 -25242
rect 21462 -25242 21536 -25222
rect 21462 -26242 21468 -25242
rect 21422 -26254 21468 -26242
rect 21730 -26242 21736 -24766
rect 21770 -26242 21776 -24766
rect 22038 -24766 22084 -24754
rect 22038 -24962 22044 -24766
rect 21976 -24982 22044 -24962
rect 22078 -24962 22084 -24766
rect 22346 -24766 22392 -24754
rect 22078 -24982 22156 -24962
rect 21976 -25042 22036 -24982
rect 22096 -25042 22156 -24982
rect 21976 -25162 22044 -25042
rect 22078 -25162 22156 -25042
rect 21976 -25222 22036 -25162
rect 22096 -25222 22156 -25162
rect 21976 -25242 22044 -25222
rect 21730 -26254 21776 -26242
rect 22038 -26242 22044 -25242
rect 22078 -25242 22156 -25222
rect 22078 -26242 22084 -25242
rect 22038 -26254 22084 -26242
rect 22346 -26242 22352 -24766
rect 22386 -26242 22392 -24766
rect 22654 -24766 22700 -24754
rect 22654 -24962 22660 -24766
rect 22596 -24982 22660 -24962
rect 22694 -24962 22700 -24766
rect 23418 -24774 23510 -24768
rect 23418 -24808 23430 -24774
rect 23498 -24808 23510 -24774
rect 23418 -24814 23510 -24808
rect 23576 -24774 23668 -24768
rect 23576 -24808 23588 -24774
rect 23656 -24808 23668 -24774
rect 23576 -24814 23668 -24808
rect 23856 -24774 23876 -24742
rect 23936 -24774 24036 -24742
rect 23856 -24808 23870 -24774
rect 23938 -24808 24028 -24774
rect 24096 -24808 24116 -24742
rect 24816 -24722 24856 -24642
rect 24936 -24722 24976 -24642
rect 24816 -24762 24976 -24722
rect 23856 -24812 24116 -24808
rect 24298 -24774 24390 -24768
rect 24298 -24808 24310 -24774
rect 24378 -24808 24390 -24774
rect 23858 -24814 23950 -24812
rect 24016 -24814 24108 -24812
rect 24298 -24814 24390 -24808
rect 24456 -24774 24548 -24768
rect 24456 -24808 24468 -24774
rect 24536 -24808 24548 -24774
rect 24456 -24814 24548 -24808
rect 24816 -24842 24856 -24762
rect 24936 -24842 24976 -24762
rect 25656 -24742 25916 -24672
rect 25218 -24774 25310 -24768
rect 25218 -24808 25230 -24774
rect 25298 -24808 25310 -24774
rect 25218 -24814 25310 -24808
rect 25376 -24774 25468 -24768
rect 25376 -24808 25388 -24774
rect 25456 -24808 25468 -24774
rect 25376 -24814 25468 -24808
rect 25656 -24774 25676 -24742
rect 25736 -24774 25836 -24742
rect 25656 -24808 25670 -24774
rect 25738 -24808 25828 -24774
rect 25896 -24808 25916 -24742
rect 26696 -24682 26716 -24602
rect 26796 -24682 26856 -24602
rect 26936 -24682 26996 -24602
rect 27076 -24682 27096 -24602
rect 28816 -24642 28976 -24602
rect 26696 -24722 27096 -24682
rect 25656 -24812 25916 -24808
rect 26098 -24774 26190 -24768
rect 26098 -24808 26110 -24774
rect 26178 -24808 26190 -24774
rect 25658 -24814 25750 -24812
rect 25816 -24814 25908 -24812
rect 26098 -24814 26190 -24808
rect 26256 -24774 26348 -24768
rect 26256 -24808 26268 -24774
rect 26336 -24808 26348 -24774
rect 26256 -24814 26348 -24808
rect 26696 -24802 26716 -24722
rect 26796 -24802 26856 -24722
rect 26936 -24802 26996 -24722
rect 27076 -24802 27096 -24722
rect 27856 -24742 28116 -24672
rect 23362 -24858 23408 -24846
rect 22694 -24982 22776 -24962
rect 22596 -25042 22636 -24982
rect 22696 -25042 22776 -24982
rect 22596 -25162 22660 -25042
rect 22694 -25162 22776 -25042
rect 22596 -25222 22636 -25162
rect 22696 -25222 22776 -25162
rect 22596 -25242 22660 -25222
rect 22346 -26254 22392 -26242
rect 22654 -26242 22660 -25242
rect 22694 -25242 22776 -25222
rect 22694 -26242 22700 -25242
rect 23362 -25784 23368 -24858
rect 23402 -25784 23408 -24858
rect 23362 -25796 23408 -25784
rect 23520 -24858 23566 -24846
rect 23520 -25784 23526 -24858
rect 23560 -25784 23566 -24858
rect 23520 -25796 23566 -25784
rect 23678 -24858 23724 -24846
rect 23678 -25784 23684 -24858
rect 23718 -25784 23724 -24858
rect 23802 -24858 23848 -24846
rect 23802 -24942 23808 -24858
rect 23776 -24962 23808 -24942
rect 23842 -24942 23848 -24858
rect 23960 -24858 24006 -24846
rect 23960 -24862 23966 -24858
rect 23842 -24962 23876 -24942
rect 23776 -25022 23796 -24962
rect 23856 -25022 23876 -24962
rect 23776 -25042 23808 -25022
rect 23842 -25042 23876 -25022
rect 23776 -25102 23796 -25042
rect 23856 -25102 23876 -25042
rect 23776 -25122 23808 -25102
rect 23842 -25122 23876 -25102
rect 23776 -25182 23796 -25122
rect 23856 -25182 23876 -25122
rect 23776 -25202 23808 -25182
rect 23678 -25796 23724 -25784
rect 23802 -25784 23808 -25202
rect 23842 -25202 23876 -25182
rect 23842 -25784 23848 -25202
rect 23802 -25796 23848 -25784
rect 23916 -25784 23966 -24862
rect 24000 -24862 24006 -24858
rect 24118 -24858 24164 -24846
rect 24000 -25784 24056 -24862
rect 24118 -24942 24124 -24858
rect 24096 -24962 24124 -24942
rect 24158 -24942 24164 -24858
rect 24242 -24858 24288 -24846
rect 24158 -24962 24196 -24942
rect 24096 -25022 24116 -24962
rect 24176 -25022 24196 -24962
rect 24096 -25042 24124 -25022
rect 24158 -25042 24196 -25022
rect 24096 -25102 24116 -25042
rect 24176 -25102 24196 -25042
rect 24096 -25122 24124 -25102
rect 24158 -25122 24196 -25102
rect 24096 -25182 24116 -25122
rect 24176 -25182 24196 -25122
rect 24096 -25202 24124 -25182
rect 23916 -25842 24056 -25784
rect 24118 -25784 24124 -25202
rect 24158 -25202 24196 -25182
rect 24158 -25784 24164 -25202
rect 24118 -25796 24164 -25784
rect 24242 -25784 24248 -24858
rect 24282 -25784 24288 -24858
rect 24242 -25796 24288 -25784
rect 24400 -24858 24446 -24846
rect 24400 -25784 24406 -24858
rect 24440 -25784 24446 -24858
rect 24400 -25796 24446 -25784
rect 24558 -24858 24604 -24846
rect 24558 -25784 24564 -24858
rect 24598 -25784 24604 -24858
rect 24558 -25796 24604 -25784
rect 24816 -24882 24976 -24842
rect 26696 -24842 27096 -24802
rect 27418 -24774 27510 -24768
rect 27418 -24808 27430 -24774
rect 27498 -24808 27510 -24774
rect 27418 -24814 27510 -24808
rect 27576 -24774 27668 -24768
rect 27576 -24808 27588 -24774
rect 27656 -24808 27668 -24774
rect 27576 -24814 27668 -24808
rect 27856 -24774 27876 -24742
rect 27936 -24774 28036 -24742
rect 27856 -24808 27870 -24774
rect 27938 -24808 28028 -24774
rect 28096 -24808 28116 -24742
rect 28816 -24722 28856 -24642
rect 28936 -24722 28976 -24642
rect 28816 -24762 28976 -24722
rect 27856 -24812 28116 -24808
rect 28298 -24774 28390 -24768
rect 28298 -24808 28310 -24774
rect 28378 -24808 28390 -24774
rect 27858 -24814 27950 -24812
rect 28016 -24814 28108 -24812
rect 28298 -24814 28390 -24808
rect 28456 -24774 28548 -24768
rect 28456 -24808 28468 -24774
rect 28536 -24808 28548 -24774
rect 28456 -24814 28548 -24808
rect 24816 -24962 24856 -24882
rect 24936 -24962 24976 -24882
rect 24816 -25002 24976 -24962
rect 24816 -25082 24856 -25002
rect 24936 -25082 24976 -25002
rect 24816 -25122 24976 -25082
rect 24816 -25202 24856 -25122
rect 24936 -25202 24976 -25122
rect 24816 -25242 24976 -25202
rect 24816 -25322 24856 -25242
rect 24936 -25322 24976 -25242
rect 24816 -25362 24976 -25322
rect 24816 -25442 24856 -25362
rect 24936 -25442 24976 -25362
rect 24816 -25482 24976 -25442
rect 24816 -25562 24856 -25482
rect 24936 -25562 24976 -25482
rect 24816 -25602 24976 -25562
rect 24816 -25682 24856 -25602
rect 24936 -25682 24976 -25602
rect 24816 -25722 24976 -25682
rect 24816 -25802 24856 -25722
rect 24936 -25802 24976 -25722
rect 25162 -24858 25208 -24846
rect 25162 -25784 25168 -24858
rect 25202 -25784 25208 -24858
rect 25162 -25796 25208 -25784
rect 25320 -24858 25366 -24846
rect 25320 -25784 25326 -24858
rect 25360 -25784 25366 -24858
rect 25320 -25796 25366 -25784
rect 25478 -24858 25524 -24846
rect 25478 -25784 25484 -24858
rect 25518 -25784 25524 -24858
rect 25602 -24858 25648 -24846
rect 25602 -25542 25608 -24858
rect 25478 -25796 25524 -25784
rect 25576 -25562 25608 -25542
rect 25642 -25542 25648 -24858
rect 25760 -24858 25806 -24846
rect 25760 -24862 25766 -24858
rect 25642 -25562 25676 -25542
rect 25576 -25622 25596 -25562
rect 25656 -25622 25676 -25562
rect 25576 -25642 25608 -25622
rect 25642 -25642 25676 -25622
rect 25576 -25702 25596 -25642
rect 25656 -25702 25676 -25642
rect 25576 -25722 25608 -25702
rect 25642 -25722 25676 -25702
rect 25576 -25782 25596 -25722
rect 25656 -25782 25676 -25722
rect 25576 -25784 25608 -25782
rect 25642 -25784 25676 -25782
rect 25576 -25802 25676 -25784
rect 25716 -25784 25766 -24862
rect 25800 -24862 25806 -24858
rect 25918 -24858 25964 -24846
rect 25800 -25784 25856 -24862
rect 25918 -25542 25924 -24858
rect 24816 -25842 24976 -25802
rect 25716 -25842 25856 -25784
rect 25896 -25562 25924 -25542
rect 25958 -25542 25964 -24858
rect 26042 -24858 26088 -24846
rect 25958 -25562 25996 -25542
rect 25896 -25622 25916 -25562
rect 25976 -25622 25996 -25562
rect 25896 -25642 25924 -25622
rect 25958 -25642 25996 -25622
rect 25896 -25702 25916 -25642
rect 25976 -25702 25996 -25642
rect 25896 -25722 25924 -25702
rect 25958 -25722 25996 -25702
rect 25896 -25782 25916 -25722
rect 25976 -25782 25996 -25722
rect 25896 -25784 25924 -25782
rect 25958 -25784 25996 -25782
rect 25896 -25802 25996 -25784
rect 26042 -25784 26048 -24858
rect 26082 -25784 26088 -24858
rect 26042 -25796 26088 -25784
rect 26200 -24858 26246 -24846
rect 26200 -25784 26206 -24858
rect 26240 -25784 26246 -24858
rect 26200 -25796 26246 -25784
rect 26358 -24858 26404 -24846
rect 26358 -25784 26364 -24858
rect 26398 -25784 26404 -24858
rect 26358 -25796 26404 -25784
rect 26696 -24922 26716 -24842
rect 26796 -24922 26856 -24842
rect 26936 -24922 26996 -24842
rect 27076 -24922 27096 -24842
rect 28816 -24842 28856 -24762
rect 28936 -24842 28976 -24762
rect 29656 -24742 29916 -24672
rect 29218 -24774 29310 -24768
rect 29218 -24808 29230 -24774
rect 29298 -24808 29310 -24774
rect 29218 -24814 29310 -24808
rect 29376 -24774 29468 -24768
rect 29376 -24808 29388 -24774
rect 29456 -24808 29468 -24774
rect 29376 -24814 29468 -24808
rect 29656 -24774 29676 -24742
rect 29736 -24774 29836 -24742
rect 29656 -24808 29670 -24774
rect 29738 -24808 29828 -24774
rect 29896 -24808 29916 -24742
rect 29656 -24812 29916 -24808
rect 30098 -24774 30190 -24768
rect 30098 -24808 30110 -24774
rect 30178 -24808 30190 -24774
rect 29658 -24814 29750 -24812
rect 29816 -24814 29908 -24812
rect 30098 -24814 30190 -24808
rect 30256 -24774 30348 -24768
rect 30256 -24808 30268 -24774
rect 30336 -24808 30348 -24774
rect 30256 -24814 30348 -24808
rect 31082 -24786 31128 -24774
rect 26696 -24962 27096 -24922
rect 26696 -25042 26716 -24962
rect 26796 -25042 26856 -24962
rect 26936 -25042 26996 -24962
rect 27076 -25042 27096 -24962
rect 26696 -25082 27096 -25042
rect 26696 -25162 26716 -25082
rect 26796 -25162 26856 -25082
rect 26936 -25162 26996 -25082
rect 27076 -25162 27096 -25082
rect 26696 -25202 27096 -25162
rect 26696 -25282 26716 -25202
rect 26796 -25282 26856 -25202
rect 26936 -25282 26996 -25202
rect 27076 -25282 27096 -25202
rect 26696 -25322 27096 -25282
rect 26696 -25402 26716 -25322
rect 26796 -25402 26856 -25322
rect 26936 -25402 26996 -25322
rect 27076 -25402 27096 -25322
rect 26696 -25442 27096 -25402
rect 26696 -25522 26716 -25442
rect 26796 -25522 26856 -25442
rect 26936 -25522 26996 -25442
rect 27076 -25522 27096 -25442
rect 26696 -25562 27096 -25522
rect 26696 -25642 26716 -25562
rect 26796 -25642 26856 -25562
rect 26936 -25642 26996 -25562
rect 27076 -25642 27096 -25562
rect 26696 -25682 27096 -25642
rect 26696 -25762 26716 -25682
rect 26796 -25762 26856 -25682
rect 26936 -25762 26996 -25682
rect 27076 -25762 27096 -25682
rect 26696 -25802 27096 -25762
rect 27362 -24858 27408 -24846
rect 27362 -25784 27368 -24858
rect 27402 -25784 27408 -24858
rect 27362 -25796 27408 -25784
rect 27520 -24858 27566 -24846
rect 27520 -25784 27526 -24858
rect 27560 -25784 27566 -24858
rect 27520 -25796 27566 -25784
rect 27678 -24858 27724 -24846
rect 27678 -25784 27684 -24858
rect 27718 -25784 27724 -24858
rect 27802 -24858 27848 -24846
rect 27802 -25542 27808 -24858
rect 27678 -25796 27724 -25784
rect 27776 -25562 27808 -25542
rect 27842 -25542 27848 -24858
rect 27960 -24858 28006 -24846
rect 27960 -24862 27966 -24858
rect 27842 -25562 27876 -25542
rect 27776 -25622 27796 -25562
rect 27856 -25622 27876 -25562
rect 27776 -25642 27808 -25622
rect 27842 -25642 27876 -25622
rect 27776 -25702 27796 -25642
rect 27856 -25702 27876 -25642
rect 27776 -25722 27808 -25702
rect 27842 -25722 27876 -25702
rect 27776 -25782 27796 -25722
rect 27856 -25782 27876 -25722
rect 27776 -25784 27808 -25782
rect 27842 -25784 27876 -25782
rect 27776 -25802 27876 -25784
rect 27916 -25784 27966 -24862
rect 28000 -24862 28006 -24858
rect 28118 -24858 28164 -24846
rect 28000 -25784 28056 -24862
rect 28118 -25542 28124 -24858
rect 23916 -25942 25856 -25842
rect 26696 -25882 26716 -25802
rect 26796 -25882 26856 -25802
rect 26936 -25882 26996 -25802
rect 27076 -25882 27096 -25802
rect 26696 -25922 27096 -25882
rect 26696 -26002 26716 -25922
rect 26796 -26002 26856 -25922
rect 26936 -26002 26996 -25922
rect 27076 -26002 27096 -25922
rect 27916 -25842 28056 -25784
rect 28096 -25562 28124 -25542
rect 28158 -25542 28164 -24858
rect 28242 -24858 28288 -24846
rect 28158 -25562 28196 -25542
rect 28096 -25622 28116 -25562
rect 28176 -25622 28196 -25562
rect 28096 -25642 28124 -25622
rect 28158 -25642 28196 -25622
rect 28096 -25702 28116 -25642
rect 28176 -25702 28196 -25642
rect 28096 -25722 28124 -25702
rect 28158 -25722 28196 -25702
rect 28096 -25782 28116 -25722
rect 28176 -25782 28196 -25722
rect 28096 -25784 28124 -25782
rect 28158 -25784 28196 -25782
rect 28096 -25802 28196 -25784
rect 28242 -25784 28248 -24858
rect 28282 -25784 28288 -24858
rect 28242 -25796 28288 -25784
rect 28400 -24858 28446 -24846
rect 28400 -25784 28406 -24858
rect 28440 -25784 28446 -24858
rect 28558 -24858 28604 -24846
rect 28558 -24942 28564 -24858
rect 28536 -25202 28564 -24942
rect 28400 -25796 28446 -25784
rect 28558 -25784 28564 -25202
rect 28598 -24942 28604 -24858
rect 28816 -24882 28976 -24842
rect 28598 -25202 28636 -24942
rect 28816 -24962 28856 -24882
rect 28936 -24962 28976 -24882
rect 28816 -25002 28976 -24962
rect 28816 -25082 28856 -25002
rect 28936 -25082 28976 -25002
rect 28816 -25122 28976 -25082
rect 28816 -25202 28856 -25122
rect 28936 -25202 28976 -25122
rect 28598 -25784 28604 -25202
rect 28558 -25796 28604 -25784
rect 28816 -25242 28976 -25202
rect 28816 -25322 28856 -25242
rect 28936 -25322 28976 -25242
rect 28816 -25362 28976 -25322
rect 28816 -25442 28856 -25362
rect 28936 -25442 28976 -25362
rect 28816 -25482 28976 -25442
rect 28816 -25562 28856 -25482
rect 28936 -25562 28976 -25482
rect 28816 -25602 28976 -25562
rect 28816 -25682 28856 -25602
rect 28936 -25682 28976 -25602
rect 28816 -25722 28976 -25682
rect 28816 -25802 28856 -25722
rect 28936 -25802 28976 -25722
rect 29162 -24858 29208 -24846
rect 29162 -25784 29168 -24858
rect 29202 -25784 29208 -24858
rect 29162 -25796 29208 -25784
rect 29320 -24858 29366 -24846
rect 29320 -25784 29326 -24858
rect 29360 -25784 29366 -24858
rect 29320 -25796 29366 -25784
rect 29478 -24858 29524 -24846
rect 29478 -25784 29484 -24858
rect 29518 -25784 29524 -24858
rect 29602 -24858 29648 -24846
rect 29602 -24942 29608 -24858
rect 29576 -24962 29608 -24942
rect 29642 -24942 29648 -24858
rect 29760 -24858 29806 -24846
rect 29760 -24862 29766 -24858
rect 29642 -24962 29676 -24942
rect 29576 -25022 29596 -24962
rect 29656 -25022 29676 -24962
rect 29576 -25042 29608 -25022
rect 29642 -25042 29676 -25022
rect 29576 -25102 29596 -25042
rect 29656 -25102 29676 -25042
rect 29576 -25122 29608 -25102
rect 29642 -25122 29676 -25102
rect 29576 -25182 29596 -25122
rect 29656 -25182 29676 -25122
rect 29576 -25202 29608 -25182
rect 29478 -25796 29524 -25784
rect 29602 -25784 29608 -25202
rect 29642 -25202 29676 -25182
rect 29642 -25784 29648 -25202
rect 29602 -25796 29648 -25784
rect 29716 -25784 29766 -24862
rect 29800 -24862 29806 -24858
rect 29918 -24858 29964 -24846
rect 29800 -25784 29856 -24862
rect 29918 -24942 29924 -24858
rect 29896 -24962 29924 -24942
rect 29958 -24942 29964 -24858
rect 30042 -24858 30088 -24846
rect 29958 -24962 29996 -24942
rect 29896 -25022 29916 -24962
rect 29976 -25022 29996 -24962
rect 29896 -25042 29924 -25022
rect 29958 -25042 29996 -25022
rect 29896 -25102 29916 -25042
rect 29976 -25102 29996 -25042
rect 29896 -25122 29924 -25102
rect 29958 -25122 29996 -25102
rect 29896 -25182 29916 -25122
rect 29976 -25182 29996 -25122
rect 29896 -25202 29924 -25182
rect 28816 -25842 28976 -25802
rect 29716 -25842 29856 -25784
rect 29918 -25784 29924 -25202
rect 29958 -25202 29996 -25182
rect 29958 -25784 29964 -25202
rect 29918 -25796 29964 -25784
rect 30042 -25784 30048 -24858
rect 30082 -25784 30088 -24858
rect 30042 -25796 30088 -25784
rect 30200 -24858 30246 -24846
rect 30200 -25784 30206 -24858
rect 30240 -25784 30246 -24858
rect 30200 -25796 30246 -25784
rect 30358 -24858 30404 -24846
rect 30358 -25784 30364 -24858
rect 30398 -25784 30404 -24858
rect 31082 -24962 31088 -24786
rect 31016 -24982 31088 -24962
rect 31122 -24962 31128 -24786
rect 31390 -24786 31436 -24774
rect 31122 -24982 31196 -24962
rect 31016 -25042 31076 -24982
rect 31136 -25042 31196 -24982
rect 31016 -25162 31088 -25042
rect 31122 -25162 31196 -25042
rect 31016 -25222 31076 -25162
rect 31136 -25222 31196 -25162
rect 31016 -25242 31088 -25222
rect 30358 -25796 30404 -25784
rect 27916 -25942 29856 -25842
rect 26696 -26042 27096 -26002
rect 22654 -26254 22700 -26242
rect 31082 -26262 31088 -25242
rect 31122 -25242 31196 -25222
rect 31122 -26262 31128 -25242
rect 31082 -26274 31128 -26262
rect 31390 -26262 31396 -24786
rect 31430 -26262 31436 -24786
rect 31698 -24786 31744 -24774
rect 31698 -24962 31704 -24786
rect 31656 -24982 31704 -24962
rect 31738 -24962 31744 -24786
rect 32006 -24786 32052 -24774
rect 31738 -24982 31836 -24962
rect 31656 -25042 31696 -24982
rect 31756 -25042 31836 -24982
rect 31656 -25162 31704 -25042
rect 31738 -25162 31836 -25042
rect 31656 -25222 31696 -25162
rect 31756 -25222 31836 -25162
rect 31656 -25242 31704 -25222
rect 31390 -26274 31436 -26262
rect 31698 -26262 31704 -25242
rect 31738 -25242 31836 -25222
rect 31738 -26262 31744 -25242
rect 31698 -26274 31744 -26262
rect 32006 -26262 32012 -24786
rect 32046 -26262 32052 -24786
rect 32314 -24786 32360 -24774
rect 32314 -24962 32320 -24786
rect 32236 -24982 32320 -24962
rect 32354 -24962 32360 -24786
rect 32354 -24982 32416 -24962
rect 32236 -25042 32296 -24982
rect 32356 -25042 32416 -24982
rect 32236 -25162 32320 -25042
rect 32354 -25162 32416 -25042
rect 32236 -25222 32296 -25162
rect 32356 -25222 32416 -25162
rect 32236 -25242 32320 -25222
rect 32006 -26274 32052 -26262
rect 32314 -26262 32320 -25242
rect 32354 -25242 32416 -25222
rect 32354 -26262 32360 -25242
rect 32314 -26274 32360 -26262
rect 21478 -26292 21720 -26286
rect 21478 -26302 21490 -26292
rect 21476 -26326 21490 -26302
rect 21708 -26302 21720 -26292
rect 21786 -26292 22028 -26286
rect 21786 -26302 21798 -26292
rect 21708 -26326 21798 -26302
rect 22016 -26302 22028 -26292
rect 22094 -26292 22336 -26286
rect 22094 -26302 22106 -26292
rect 22016 -26326 22106 -26302
rect 22324 -26302 22336 -26292
rect 22402 -26292 22644 -26286
rect 22402 -26302 22414 -26292
rect 22324 -26326 22414 -26302
rect 22632 -26302 22644 -26292
rect 22632 -26326 22656 -26302
rect 31138 -26312 31380 -26306
rect 21476 -26502 22656 -26326
rect 23998 -26324 24090 -26318
rect 23998 -26358 24010 -26324
rect 24078 -26358 24090 -26324
rect 23998 -26364 24090 -26358
rect 24156 -26324 24248 -26318
rect 24156 -26358 24168 -26324
rect 24236 -26358 24248 -26324
rect 24156 -26364 24248 -26358
rect 24438 -26324 24680 -26318
rect 24438 -26358 24450 -26324
rect 24668 -26358 24680 -26324
rect 24438 -26364 24680 -26358
rect 24746 -26324 24988 -26318
rect 24746 -26358 24758 -26324
rect 24976 -26358 24988 -26324
rect 24746 -26364 24988 -26358
rect 25054 -26324 25296 -26318
rect 25054 -26358 25066 -26324
rect 25284 -26358 25296 -26324
rect 25054 -26364 25296 -26358
rect 25362 -26324 25604 -26318
rect 25362 -26358 25374 -26324
rect 25592 -26358 25604 -26324
rect 25362 -26364 25604 -26358
rect 25670 -26324 25912 -26318
rect 25670 -26358 25682 -26324
rect 25900 -26358 25912 -26324
rect 25670 -26364 25912 -26358
rect 25978 -26324 26220 -26318
rect 25978 -26358 25990 -26324
rect 26208 -26358 26220 -26324
rect 25978 -26364 26220 -26358
rect 26286 -26324 26528 -26318
rect 26286 -26358 26298 -26324
rect 26516 -26358 26528 -26324
rect 26286 -26364 26528 -26358
rect 26594 -26324 26836 -26318
rect 26594 -26358 26606 -26324
rect 26824 -26358 26836 -26324
rect 26594 -26364 26836 -26358
rect 26902 -26324 27144 -26318
rect 26902 -26358 26914 -26324
rect 27132 -26358 27144 -26324
rect 26902 -26364 27144 -26358
rect 27210 -26324 27452 -26318
rect 27210 -26358 27222 -26324
rect 27440 -26358 27452 -26324
rect 27210 -26364 27452 -26358
rect 27518 -26324 27760 -26318
rect 27518 -26358 27530 -26324
rect 27748 -26358 27760 -26324
rect 27518 -26364 27760 -26358
rect 27826 -26324 28068 -26318
rect 27826 -26358 27838 -26324
rect 28056 -26358 28068 -26324
rect 27826 -26364 28068 -26358
rect 28134 -26324 28376 -26318
rect 28134 -26358 28146 -26324
rect 28364 -26358 28376 -26324
rect 28134 -26364 28376 -26358
rect 28442 -26324 28684 -26318
rect 28442 -26358 28454 -26324
rect 28672 -26358 28684 -26324
rect 28442 -26364 28684 -26358
rect 28750 -26324 28992 -26318
rect 28750 -26358 28762 -26324
rect 28980 -26358 28992 -26324
rect 28750 -26364 28992 -26358
rect 29058 -26324 29300 -26318
rect 29058 -26358 29070 -26324
rect 29288 -26358 29300 -26324
rect 29058 -26364 29300 -26358
rect 29498 -26324 29590 -26318
rect 29498 -26358 29510 -26324
rect 29578 -26358 29590 -26324
rect 29498 -26364 29590 -26358
rect 29656 -26324 29748 -26318
rect 31138 -26322 31150 -26312
rect 29656 -26358 29668 -26324
rect 29736 -26358 29748 -26324
rect 29656 -26364 29748 -26358
rect 31136 -26346 31150 -26322
rect 31368 -26322 31380 -26312
rect 31446 -26312 31688 -26306
rect 31446 -26322 31458 -26312
rect 31368 -26346 31458 -26322
rect 31676 -26322 31688 -26312
rect 31754 -26312 31996 -26306
rect 31754 -26322 31766 -26312
rect 31676 -26346 31766 -26322
rect 31984 -26322 31996 -26312
rect 32062 -26312 32304 -26306
rect 32062 -26322 32074 -26312
rect 31984 -26346 32074 -26322
rect 32292 -26322 32304 -26312
rect 32292 -26346 32316 -26322
rect 21476 -26562 21496 -26502
rect 21556 -26562 21576 -26502
rect 21636 -26562 21656 -26502
rect 21716 -26562 21736 -26502
rect 21796 -26562 21816 -26502
rect 21876 -26562 21896 -26502
rect 21956 -26562 21976 -26502
rect 22036 -26562 22056 -26502
rect 22116 -26562 22136 -26502
rect 22196 -26562 22216 -26502
rect 22276 -26562 22296 -26502
rect 22356 -26562 22376 -26502
rect 22436 -26562 22456 -26502
rect 22556 -26562 22576 -26502
rect 22636 -26562 22656 -26502
rect 21476 -26602 22656 -26562
rect 21476 -26662 21496 -26602
rect 21556 -26662 21576 -26602
rect 21636 -26662 21656 -26602
rect 21716 -26662 21736 -26602
rect 21796 -26662 21816 -26602
rect 21876 -26662 21896 -26602
rect 21956 -26662 21976 -26602
rect 22036 -26662 22056 -26602
rect 22116 -26662 22136 -26602
rect 22196 -26662 22216 -26602
rect 22276 -26662 22296 -26602
rect 22356 -26662 22376 -26602
rect 22436 -26662 22456 -26602
rect 22556 -26662 22576 -26602
rect 22636 -26662 22656 -26602
rect 21476 -26682 22656 -26662
rect 23942 -26408 23988 -26396
rect 23942 -27884 23948 -26408
rect 23982 -27884 23988 -26408
rect 23942 -27896 23988 -27884
rect 24100 -26408 24146 -26396
rect 24100 -27884 24106 -26408
rect 24140 -27884 24146 -26408
rect 24100 -27896 24146 -27884
rect 24258 -26408 24304 -26396
rect 24258 -27884 24264 -26408
rect 24298 -27884 24304 -26408
rect 24382 -26408 24428 -26396
rect 24382 -26482 24388 -26408
rect 24376 -26502 24388 -26482
rect 24422 -26482 24428 -26408
rect 24690 -26408 24736 -26396
rect 24422 -26502 24536 -26482
rect 24436 -26562 24476 -26502
rect 24376 -26582 24388 -26562
rect 24422 -26582 24536 -26562
rect 24436 -26642 24476 -26582
rect 24376 -26762 24388 -26642
rect 24422 -26762 24536 -26642
rect 24436 -26822 24476 -26762
rect 24376 -26842 24388 -26822
rect 24422 -26842 24536 -26822
rect 24436 -26902 24476 -26842
rect 24376 -26922 24388 -26902
rect 24382 -27102 24388 -26922
rect 24376 -27122 24388 -27102
rect 24422 -26922 24536 -26902
rect 24422 -27102 24428 -26922
rect 24422 -27122 24536 -27102
rect 24436 -27182 24476 -27122
rect 24376 -27202 24388 -27182
rect 24422 -27202 24536 -27182
rect 24436 -27262 24476 -27202
rect 24376 -27342 24388 -27262
rect 24422 -27342 24536 -27262
rect 24436 -27402 24476 -27342
rect 24376 -27422 24388 -27402
rect 24422 -27422 24536 -27402
rect 24436 -27482 24476 -27422
rect 24376 -27502 24388 -27482
rect 24258 -27896 24304 -27884
rect 24382 -27884 24388 -27502
rect 24422 -27502 24536 -27482
rect 24422 -27884 24428 -27502
rect 24382 -27896 24428 -27884
rect 24690 -27884 24696 -26408
rect 24730 -27884 24736 -26408
rect 24998 -26408 25044 -26396
rect 24998 -26482 25004 -26408
rect 24936 -26522 25004 -26482
rect 25038 -26482 25044 -26408
rect 25306 -26408 25352 -26396
rect 25038 -26522 25116 -26482
rect 24936 -26582 24956 -26522
rect 25096 -26582 25116 -26522
rect 24936 -26602 25004 -26582
rect 25038 -26602 25116 -26582
rect 24936 -26662 24956 -26602
rect 25096 -26662 25116 -26602
rect 24936 -26682 25004 -26662
rect 25038 -26682 25116 -26662
rect 24936 -26742 24956 -26682
rect 25096 -26742 25116 -26682
rect 24936 -26762 25004 -26742
rect 25038 -26762 25116 -26742
rect 24936 -26822 24956 -26762
rect 25096 -26822 25116 -26762
rect 24936 -26842 25004 -26822
rect 25038 -26842 25116 -26822
rect 24936 -26902 24956 -26842
rect 25096 -26902 25116 -26842
rect 24936 -26922 25004 -26902
rect 24690 -27896 24736 -27884
rect 24998 -27884 25004 -26922
rect 25038 -26922 25116 -26902
rect 25038 -27884 25044 -26922
rect 24998 -27896 25044 -27884
rect 25306 -27884 25312 -26408
rect 25346 -27884 25352 -26408
rect 25614 -26408 25660 -26396
rect 25614 -27102 25620 -26408
rect 25556 -27122 25620 -27102
rect 25616 -27182 25620 -27122
rect 25556 -27202 25620 -27182
rect 25616 -27262 25620 -27202
rect 25556 -27342 25620 -27262
rect 25616 -27402 25620 -27342
rect 25556 -27422 25620 -27402
rect 25616 -27482 25620 -27422
rect 25556 -27502 25620 -27482
rect 25306 -27896 25352 -27884
rect 25614 -27884 25620 -27502
rect 25654 -27102 25660 -26408
rect 25922 -26408 25968 -26396
rect 25654 -27122 25716 -27102
rect 25654 -27182 25656 -27122
rect 25654 -27202 25716 -27182
rect 25654 -27262 25656 -27202
rect 25654 -27342 25716 -27262
rect 25654 -27402 25656 -27342
rect 25654 -27422 25716 -27402
rect 25654 -27482 25656 -27422
rect 25654 -27502 25716 -27482
rect 25654 -27884 25660 -27502
rect 25614 -27896 25660 -27884
rect 25922 -27884 25928 -26408
rect 25962 -27884 25968 -26408
rect 26230 -26408 26276 -26396
rect 26230 -26482 26236 -26408
rect 26156 -26522 26236 -26482
rect 26270 -26482 26276 -26408
rect 26538 -26408 26584 -26396
rect 26270 -26522 26336 -26482
rect 26156 -26582 26176 -26522
rect 26316 -26582 26336 -26522
rect 26156 -26602 26236 -26582
rect 26270 -26602 26336 -26582
rect 26156 -26662 26176 -26602
rect 26316 -26662 26336 -26602
rect 26156 -26682 26236 -26662
rect 26270 -26682 26336 -26662
rect 26156 -26742 26176 -26682
rect 26316 -26742 26336 -26682
rect 26156 -26762 26236 -26742
rect 26270 -26762 26336 -26742
rect 26156 -26822 26176 -26762
rect 26316 -26822 26336 -26762
rect 26156 -26842 26236 -26822
rect 26270 -26842 26336 -26822
rect 26156 -26902 26176 -26842
rect 26316 -26902 26336 -26842
rect 26156 -26922 26236 -26902
rect 25922 -27896 25968 -27884
rect 26230 -27884 26236 -26922
rect 26270 -26922 26336 -26902
rect 26270 -27884 26276 -26922
rect 26230 -27896 26276 -27884
rect 26538 -27884 26544 -26408
rect 26578 -27884 26584 -26408
rect 26846 -26408 26892 -26396
rect 26846 -27102 26852 -26408
rect 26796 -27122 26852 -27102
rect 26886 -27102 26892 -26408
rect 27154 -26408 27200 -26396
rect 26886 -27122 26956 -27102
rect 26886 -27182 26896 -27122
rect 26796 -27202 26852 -27182
rect 26886 -27202 26956 -27182
rect 26886 -27262 26896 -27202
rect 26796 -27342 26852 -27262
rect 26886 -27342 26956 -27262
rect 26886 -27402 26896 -27342
rect 26796 -27422 26852 -27402
rect 26886 -27422 26956 -27402
rect 26886 -27482 26896 -27422
rect 26796 -27502 26852 -27482
rect 26538 -27896 26584 -27884
rect 26846 -27884 26852 -27502
rect 26886 -27502 26956 -27482
rect 26886 -27884 26892 -27502
rect 26846 -27896 26892 -27884
rect 27154 -27884 27160 -26408
rect 27194 -27884 27200 -26408
rect 27462 -26408 27508 -26396
rect 27462 -26482 27468 -26408
rect 27396 -26522 27468 -26482
rect 27502 -26482 27508 -26408
rect 27770 -26408 27816 -26396
rect 27502 -26522 27576 -26482
rect 27396 -26582 27416 -26522
rect 27556 -26582 27576 -26522
rect 27396 -26602 27468 -26582
rect 27502 -26602 27576 -26582
rect 27396 -26662 27416 -26602
rect 27556 -26662 27576 -26602
rect 27396 -26682 27468 -26662
rect 27502 -26682 27576 -26662
rect 27396 -26742 27416 -26682
rect 27556 -26742 27576 -26682
rect 27396 -26762 27468 -26742
rect 27502 -26762 27576 -26742
rect 27396 -26822 27416 -26762
rect 27556 -26822 27576 -26762
rect 27396 -26842 27468 -26822
rect 27502 -26842 27576 -26822
rect 27396 -26902 27416 -26842
rect 27556 -26902 27576 -26842
rect 27396 -26922 27468 -26902
rect 27154 -27896 27200 -27884
rect 27462 -27884 27468 -26922
rect 27502 -26922 27576 -26902
rect 27502 -27884 27508 -26922
rect 27462 -27896 27508 -27884
rect 27770 -27884 27776 -26408
rect 27810 -27884 27816 -26408
rect 28078 -26408 28124 -26396
rect 28078 -27102 28084 -26408
rect 28016 -27122 28084 -27102
rect 28118 -27102 28124 -26408
rect 28386 -26408 28432 -26396
rect 28118 -27122 28176 -27102
rect 28076 -27182 28084 -27122
rect 28016 -27202 28084 -27182
rect 28118 -27202 28176 -27182
rect 28076 -27262 28084 -27202
rect 28016 -27342 28084 -27262
rect 28118 -27342 28176 -27262
rect 28076 -27402 28084 -27342
rect 28016 -27422 28084 -27402
rect 28118 -27422 28176 -27402
rect 28076 -27482 28084 -27422
rect 28016 -27502 28084 -27482
rect 27770 -27896 27816 -27884
rect 28078 -27884 28084 -27502
rect 28118 -27502 28176 -27482
rect 28118 -27884 28124 -27502
rect 28078 -27896 28124 -27884
rect 28386 -27884 28392 -26408
rect 28426 -27884 28432 -26408
rect 28694 -26408 28740 -26396
rect 28694 -26482 28700 -26408
rect 28616 -26522 28700 -26482
rect 28734 -26482 28740 -26408
rect 29002 -26408 29048 -26396
rect 28734 -26522 28796 -26482
rect 28616 -26582 28636 -26522
rect 28696 -26582 28700 -26522
rect 28776 -26582 28796 -26522
rect 28616 -26602 28700 -26582
rect 28734 -26602 28796 -26582
rect 28616 -26662 28636 -26602
rect 28696 -26662 28700 -26602
rect 28776 -26662 28796 -26602
rect 28616 -26682 28700 -26662
rect 28734 -26682 28796 -26662
rect 28616 -26742 28636 -26682
rect 28696 -26742 28700 -26682
rect 28776 -26742 28796 -26682
rect 28616 -26762 28700 -26742
rect 28734 -26762 28796 -26742
rect 28616 -26822 28636 -26762
rect 28696 -26822 28700 -26762
rect 28776 -26822 28796 -26762
rect 28616 -26842 28700 -26822
rect 28734 -26842 28796 -26822
rect 28616 -26902 28636 -26842
rect 28696 -26902 28700 -26842
rect 28776 -26902 28796 -26842
rect 28616 -26922 28700 -26902
rect 28386 -27896 28432 -27884
rect 28694 -27884 28700 -26922
rect 28734 -26922 28796 -26902
rect 28734 -27884 28740 -26922
rect 28694 -27896 28740 -27884
rect 29002 -27884 29008 -26408
rect 29042 -27884 29048 -26408
rect 29310 -26408 29356 -26396
rect 29310 -26482 29316 -26408
rect 29216 -26502 29316 -26482
rect 29350 -26482 29356 -26408
rect 29442 -26408 29488 -26396
rect 29350 -26502 29376 -26482
rect 29276 -26562 29316 -26502
rect 29216 -26582 29316 -26562
rect 29350 -26582 29376 -26562
rect 29276 -26642 29316 -26582
rect 29216 -26762 29316 -26642
rect 29350 -26762 29376 -26642
rect 29276 -26822 29316 -26762
rect 29216 -26842 29316 -26822
rect 29350 -26842 29376 -26822
rect 29276 -26902 29316 -26842
rect 29216 -26922 29316 -26902
rect 29310 -27102 29316 -26922
rect 29216 -27122 29316 -27102
rect 29350 -26922 29376 -26902
rect 29350 -27102 29356 -26922
rect 29350 -27122 29376 -27102
rect 29276 -27182 29316 -27122
rect 29216 -27202 29316 -27182
rect 29350 -27202 29376 -27182
rect 29276 -27262 29316 -27202
rect 29216 -27342 29316 -27262
rect 29350 -27342 29376 -27262
rect 29276 -27402 29316 -27342
rect 29216 -27422 29316 -27402
rect 29350 -27422 29376 -27402
rect 29276 -27482 29316 -27422
rect 29216 -27502 29316 -27482
rect 29002 -27896 29048 -27884
rect 29310 -27884 29316 -27502
rect 29350 -27502 29376 -27482
rect 29350 -27884 29356 -27502
rect 29310 -27896 29356 -27884
rect 29442 -27884 29448 -26408
rect 29482 -27884 29488 -26408
rect 29442 -27896 29488 -27884
rect 29600 -26408 29646 -26396
rect 29600 -27884 29606 -26408
rect 29640 -27884 29646 -26408
rect 29600 -27896 29646 -27884
rect 29758 -26408 29804 -26396
rect 29758 -27884 29764 -26408
rect 29798 -27884 29804 -26408
rect 31136 -26502 32316 -26346
rect 31136 -26562 31156 -26502
rect 31216 -26562 31236 -26502
rect 31336 -26562 31356 -26502
rect 31416 -26562 31436 -26502
rect 31496 -26562 31516 -26502
rect 31576 -26562 31596 -26502
rect 31656 -26562 31676 -26502
rect 31736 -26562 31756 -26502
rect 31816 -26562 31836 -26502
rect 31896 -26562 31916 -26502
rect 31976 -26562 31996 -26502
rect 32056 -26562 32076 -26502
rect 32136 -26562 32156 -26502
rect 32216 -26562 32236 -26502
rect 32296 -26562 32316 -26502
rect 31136 -26602 32316 -26562
rect 31136 -26662 31156 -26602
rect 31216 -26662 31236 -26602
rect 31336 -26662 31356 -26602
rect 31416 -26662 31436 -26602
rect 31496 -26662 31516 -26602
rect 31576 -26662 31596 -26602
rect 31656 -26662 31676 -26602
rect 31736 -26662 31756 -26602
rect 31816 -26662 31836 -26602
rect 31896 -26662 31916 -26602
rect 31976 -26662 31996 -26602
rect 32056 -26662 32076 -26602
rect 32136 -26662 32156 -26602
rect 32216 -26662 32236 -26602
rect 32296 -26662 32316 -26602
rect 31136 -26682 32316 -26662
rect 29758 -27896 29804 -27884
rect 23636 -28242 30116 -28182
rect 23636 -28322 23656 -28242
rect 23736 -28322 23776 -28242
rect 23856 -28322 23896 -28242
rect 23976 -28322 24016 -28242
rect 24096 -28322 24136 -28242
rect 24216 -28322 24256 -28242
rect 24336 -28322 24376 -28242
rect 24456 -28322 24496 -28242
rect 24576 -28322 24616 -28242
rect 24696 -28322 24736 -28242
rect 24816 -28322 24856 -28242
rect 24936 -28322 24976 -28242
rect 25056 -28322 25096 -28242
rect 25176 -28322 25216 -28242
rect 25296 -28322 25336 -28242
rect 25416 -28322 25456 -28242
rect 25536 -28322 25576 -28242
rect 25656 -28322 25696 -28242
rect 25776 -28322 25816 -28242
rect 25896 -28322 25936 -28242
rect 26016 -28322 26056 -28242
rect 26136 -28322 26176 -28242
rect 26256 -28322 26296 -28242
rect 26376 -28322 26416 -28242
rect 26496 -28322 26536 -28242
rect 26616 -28322 26656 -28242
rect 26736 -28322 26776 -28242
rect 26856 -28322 26896 -28242
rect 26976 -28322 27016 -28242
rect 27096 -28322 27136 -28242
rect 27216 -28322 27256 -28242
rect 27336 -28322 27376 -28242
rect 27456 -28322 27496 -28242
rect 27576 -28322 27616 -28242
rect 27696 -28322 27736 -28242
rect 27816 -28322 27856 -28242
rect 27936 -28322 27976 -28242
rect 28056 -28322 28096 -28242
rect 28176 -28322 28216 -28242
rect 28296 -28322 28336 -28242
rect 28416 -28322 28456 -28242
rect 28536 -28322 28576 -28242
rect 28656 -28322 28696 -28242
rect 28776 -28322 28816 -28242
rect 28896 -28322 28936 -28242
rect 29016 -28322 29056 -28242
rect 29136 -28322 29176 -28242
rect 29256 -28322 29296 -28242
rect 29376 -28322 29416 -28242
rect 29496 -28322 29536 -28242
rect 29616 -28322 29656 -28242
rect 29736 -28322 29776 -28242
rect 29856 -28322 29896 -28242
rect 29976 -28322 30016 -28242
rect 30096 -28322 30116 -28242
rect 23636 -28362 30116 -28322
rect 23636 -28442 23656 -28362
rect 23736 -28442 23776 -28362
rect 23856 -28442 23896 -28362
rect 23976 -28442 24016 -28362
rect 24096 -28442 24136 -28362
rect 24216 -28442 24256 -28362
rect 24336 -28442 24376 -28362
rect 24456 -28442 24496 -28362
rect 24576 -28442 24616 -28362
rect 24696 -28442 24736 -28362
rect 24816 -28442 24856 -28362
rect 24936 -28442 24976 -28362
rect 25056 -28442 25096 -28362
rect 25176 -28442 25216 -28362
rect 25296 -28442 25336 -28362
rect 25416 -28442 25456 -28362
rect 25536 -28442 25576 -28362
rect 25656 -28442 25696 -28362
rect 25776 -28442 25816 -28362
rect 25896 -28442 25936 -28362
rect 26016 -28442 26056 -28362
rect 26136 -28442 26176 -28362
rect 26256 -28442 26296 -28362
rect 26376 -28442 26416 -28362
rect 26496 -28442 26536 -28362
rect 26616 -28442 26656 -28362
rect 26736 -28442 26776 -28362
rect 26856 -28442 26896 -28362
rect 26976 -28442 27016 -28362
rect 27096 -28442 27136 -28362
rect 27216 -28442 27256 -28362
rect 27336 -28442 27376 -28362
rect 27456 -28442 27496 -28362
rect 27576 -28442 27616 -28362
rect 27696 -28442 27736 -28362
rect 27816 -28442 27856 -28362
rect 27936 -28442 27976 -28362
rect 28056 -28442 28096 -28362
rect 28176 -28442 28216 -28362
rect 28296 -28442 28336 -28362
rect 28416 -28442 28456 -28362
rect 28536 -28442 28576 -28362
rect 28656 -28442 28696 -28362
rect 28776 -28442 28816 -28362
rect 28896 -28442 28936 -28362
rect 29016 -28442 29056 -28362
rect 29136 -28442 29176 -28362
rect 29256 -28442 29296 -28362
rect 29376 -28442 29416 -28362
rect 29496 -28442 29536 -28362
rect 29616 -28442 29656 -28362
rect 29736 -28442 29776 -28362
rect 29856 -28442 29896 -28362
rect 29976 -28442 30016 -28362
rect 30096 -28442 30116 -28362
rect 23636 -28482 30116 -28442
rect 23636 -28562 23656 -28482
rect 23736 -28562 23776 -28482
rect 23856 -28562 23896 -28482
rect 23976 -28562 24016 -28482
rect 24096 -28562 24136 -28482
rect 24216 -28562 24256 -28482
rect 24336 -28562 24376 -28482
rect 24456 -28562 24496 -28482
rect 24576 -28562 24616 -28482
rect 24696 -28562 24736 -28482
rect 24816 -28562 24856 -28482
rect 24936 -28562 24976 -28482
rect 25056 -28562 25096 -28482
rect 25176 -28562 25216 -28482
rect 25296 -28562 25336 -28482
rect 25416 -28562 25456 -28482
rect 25536 -28562 25576 -28482
rect 25656 -28562 25696 -28482
rect 25776 -28562 25816 -28482
rect 25896 -28562 25936 -28482
rect 26016 -28562 26056 -28482
rect 26136 -28562 26176 -28482
rect 26256 -28562 26296 -28482
rect 26376 -28562 26416 -28482
rect 26496 -28562 26536 -28482
rect 26616 -28562 26656 -28482
rect 26736 -28562 26776 -28482
rect 26856 -28562 26896 -28482
rect 26976 -28562 27016 -28482
rect 27096 -28562 27136 -28482
rect 27216 -28562 27256 -28482
rect 27336 -28562 27376 -28482
rect 27456 -28562 27496 -28482
rect 27576 -28562 27616 -28482
rect 27696 -28562 27736 -28482
rect 27816 -28562 27856 -28482
rect 27936 -28562 27976 -28482
rect 28056 -28562 28096 -28482
rect 28176 -28562 28216 -28482
rect 28296 -28562 28336 -28482
rect 28416 -28562 28456 -28482
rect 28536 -28562 28576 -28482
rect 28656 -28562 28696 -28482
rect 28776 -28562 28816 -28482
rect 28896 -28562 28936 -28482
rect 29016 -28562 29056 -28482
rect 29136 -28562 29176 -28482
rect 29256 -28562 29296 -28482
rect 29376 -28562 29416 -28482
rect 29496 -28562 29536 -28482
rect 29616 -28562 29656 -28482
rect 29736 -28562 29776 -28482
rect 29856 -28562 29896 -28482
rect 29976 -28562 30016 -28482
rect 30096 -28562 30116 -28482
rect 23636 -28602 30116 -28562
rect 23636 -28682 23656 -28602
rect 23736 -28682 23776 -28602
rect 23856 -28682 23896 -28602
rect 23976 -28682 24016 -28602
rect 24096 -28682 24136 -28602
rect 24216 -28682 24256 -28602
rect 24336 -28682 24376 -28602
rect 24456 -28682 24496 -28602
rect 24576 -28682 24616 -28602
rect 24696 -28682 24736 -28602
rect 24816 -28682 24856 -28602
rect 24936 -28682 24976 -28602
rect 25056 -28682 25096 -28602
rect 25176 -28682 25216 -28602
rect 25296 -28682 25336 -28602
rect 25416 -28682 25456 -28602
rect 25536 -28682 25576 -28602
rect 25656 -28682 25696 -28602
rect 25776 -28682 25816 -28602
rect 25896 -28682 25936 -28602
rect 26016 -28682 26056 -28602
rect 26136 -28682 26176 -28602
rect 26256 -28682 26296 -28602
rect 26376 -28682 26416 -28602
rect 26496 -28682 26536 -28602
rect 26616 -28682 26656 -28602
rect 26736 -28682 26776 -28602
rect 26856 -28682 26896 -28602
rect 26976 -28682 27016 -28602
rect 27096 -28682 27136 -28602
rect 27216 -28682 27256 -28602
rect 27336 -28682 27376 -28602
rect 27456 -28682 27496 -28602
rect 27576 -28682 27616 -28602
rect 27696 -28682 27736 -28602
rect 27816 -28682 27856 -28602
rect 27936 -28682 27976 -28602
rect 28056 -28682 28096 -28602
rect 28176 -28682 28216 -28602
rect 28296 -28682 28336 -28602
rect 28416 -28682 28456 -28602
rect 28536 -28682 28576 -28602
rect 28656 -28682 28696 -28602
rect 28776 -28682 28816 -28602
rect 28896 -28682 28936 -28602
rect 29016 -28682 29056 -28602
rect 29136 -28682 29176 -28602
rect 29256 -28682 29296 -28602
rect 29376 -28682 29416 -28602
rect 29496 -28682 29536 -28602
rect 29616 -28682 29656 -28602
rect 29736 -28682 29776 -28602
rect 29856 -28682 29896 -28602
rect 29976 -28682 30016 -28602
rect 30096 -28682 30116 -28602
rect 23636 -28722 30116 -28682
rect 23636 -28802 23656 -28722
rect 23736 -28802 23776 -28722
rect 23856 -28802 23896 -28722
rect 23976 -28802 24016 -28722
rect 24096 -28802 24136 -28722
rect 24216 -28802 24256 -28722
rect 24336 -28802 24376 -28722
rect 24456 -28802 24496 -28722
rect 24576 -28802 24616 -28722
rect 24696 -28802 24736 -28722
rect 24816 -28802 24856 -28722
rect 24936 -28802 24976 -28722
rect 25056 -28802 25096 -28722
rect 25176 -28802 25216 -28722
rect 25296 -28802 25336 -28722
rect 25416 -28802 25456 -28722
rect 25536 -28802 25576 -28722
rect 25656 -28802 25696 -28722
rect 25776 -28802 25816 -28722
rect 25896 -28802 25936 -28722
rect 26016 -28802 26056 -28722
rect 26136 -28802 26176 -28722
rect 26256 -28802 26296 -28722
rect 26376 -28802 26416 -28722
rect 26496 -28802 26536 -28722
rect 26616 -28802 26656 -28722
rect 26736 -28802 26776 -28722
rect 26856 -28802 26896 -28722
rect 26976 -28802 27016 -28722
rect 27096 -28802 27136 -28722
rect 27216 -28802 27256 -28722
rect 27336 -28802 27376 -28722
rect 27456 -28802 27496 -28722
rect 27576 -28802 27616 -28722
rect 27696 -28802 27736 -28722
rect 27816 -28802 27856 -28722
rect 27936 -28802 27976 -28722
rect 28056 -28802 28096 -28722
rect 28176 -28802 28216 -28722
rect 28296 -28802 28336 -28722
rect 28416 -28802 28456 -28722
rect 28536 -28802 28576 -28722
rect 28656 -28802 28696 -28722
rect 28776 -28802 28816 -28722
rect 28896 -28802 28936 -28722
rect 29016 -28802 29056 -28722
rect 29136 -28802 29176 -28722
rect 29256 -28802 29296 -28722
rect 29376 -28802 29416 -28722
rect 29496 -28802 29536 -28722
rect 29616 -28802 29656 -28722
rect 29736 -28802 29776 -28722
rect 29856 -28802 29896 -28722
rect 29976 -28802 30016 -28722
rect 30096 -28802 30116 -28722
rect 23636 -28842 30116 -28802
rect 23636 -28922 23656 -28842
rect 23736 -28922 23776 -28842
rect 23856 -28922 23896 -28842
rect 23976 -28922 24016 -28842
rect 24096 -28922 24136 -28842
rect 24216 -28922 24256 -28842
rect 24336 -28922 24376 -28842
rect 24456 -28922 24496 -28842
rect 24576 -28922 24616 -28842
rect 24696 -28922 24736 -28842
rect 24816 -28922 24856 -28842
rect 24936 -28922 24976 -28842
rect 25056 -28922 25096 -28842
rect 25176 -28922 25216 -28842
rect 25296 -28922 25336 -28842
rect 25416 -28922 25456 -28842
rect 25536 -28922 25576 -28842
rect 25656 -28922 25696 -28842
rect 25776 -28922 25816 -28842
rect 25896 -28922 25936 -28842
rect 26016 -28922 26056 -28842
rect 26136 -28922 26176 -28842
rect 26256 -28922 26296 -28842
rect 26376 -28922 26416 -28842
rect 26496 -28922 26536 -28842
rect 26616 -28922 26656 -28842
rect 26736 -28922 26776 -28842
rect 26856 -28922 26896 -28842
rect 26976 -28922 27016 -28842
rect 27096 -28922 27136 -28842
rect 27216 -28922 27256 -28842
rect 27336 -28922 27376 -28842
rect 27456 -28922 27496 -28842
rect 27576 -28922 27616 -28842
rect 27696 -28922 27736 -28842
rect 27816 -28922 27856 -28842
rect 27936 -28922 27976 -28842
rect 28056 -28922 28096 -28842
rect 28176 -28922 28216 -28842
rect 28296 -28922 28336 -28842
rect 28416 -28922 28456 -28842
rect 28536 -28922 28576 -28842
rect 28656 -28922 28696 -28842
rect 28776 -28922 28816 -28842
rect 28896 -28922 28936 -28842
rect 29016 -28922 29056 -28842
rect 29136 -28922 29176 -28842
rect 29256 -28922 29296 -28842
rect 29376 -28922 29416 -28842
rect 29496 -28922 29536 -28842
rect 29616 -28922 29656 -28842
rect 29736 -28922 29776 -28842
rect 29856 -28922 29896 -28842
rect 29976 -28922 30016 -28842
rect 30096 -28922 30116 -28842
rect 23636 -28962 30116 -28922
rect 22796 -29042 23196 -29022
rect 22796 -29122 22816 -29042
rect 22896 -29122 22956 -29042
rect 23036 -29122 23096 -29042
rect 23176 -29122 23196 -29042
rect 22796 -29182 23196 -29122
rect 23636 -29042 23656 -28962
rect 23736 -29042 23776 -28962
rect 23856 -29042 23896 -28962
rect 23976 -29042 24016 -28962
rect 24096 -29042 24136 -28962
rect 24216 -29042 24256 -28962
rect 24336 -29042 24376 -28962
rect 24456 -29042 24496 -28962
rect 24576 -29042 24616 -28962
rect 24696 -29042 24736 -28962
rect 24816 -29042 24856 -28962
rect 24936 -29042 24976 -28962
rect 25056 -29042 25096 -28962
rect 25176 -29042 25216 -28962
rect 25296 -29042 25336 -28962
rect 25416 -29042 25456 -28962
rect 25536 -29042 25576 -28962
rect 25656 -29042 25696 -28962
rect 25776 -29042 25816 -28962
rect 25896 -29042 25936 -28962
rect 26016 -29042 26056 -28962
rect 26136 -29042 26176 -28962
rect 26256 -29042 26296 -28962
rect 26376 -29042 26416 -28962
rect 26496 -29042 26536 -28962
rect 26616 -29042 26656 -28962
rect 26736 -29042 26776 -28962
rect 26856 -29042 26896 -28962
rect 26976 -29042 27016 -28962
rect 27096 -29042 27136 -28962
rect 27216 -29042 27256 -28962
rect 27336 -29042 27376 -28962
rect 27456 -29042 27496 -28962
rect 27576 -29042 27616 -28962
rect 27696 -29042 27736 -28962
rect 27816 -29042 27856 -28962
rect 27936 -29042 27976 -28962
rect 28056 -29042 28096 -28962
rect 28176 -29042 28216 -28962
rect 28296 -29042 28336 -28962
rect 28416 -29042 28456 -28962
rect 28536 -29042 28576 -28962
rect 28656 -29042 28696 -28962
rect 28776 -29042 28816 -28962
rect 28896 -29042 28936 -28962
rect 29016 -29042 29056 -28962
rect 29136 -29042 29176 -28962
rect 29256 -29042 29296 -28962
rect 29376 -29042 29416 -28962
rect 29496 -29042 29536 -28962
rect 29616 -29042 29656 -28962
rect 29736 -29042 29776 -28962
rect 29856 -29042 29896 -28962
rect 29976 -29042 30016 -28962
rect 30096 -29042 30116 -28962
rect 23636 -29082 30116 -29042
rect 23636 -29162 23656 -29082
rect 23736 -29162 23776 -29082
rect 23856 -29162 23896 -29082
rect 23976 -29162 24016 -29082
rect 24096 -29162 24136 -29082
rect 24216 -29162 24256 -29082
rect 24336 -29162 24376 -29082
rect 24456 -29162 24496 -29082
rect 24576 -29162 24616 -29082
rect 24696 -29162 24736 -29082
rect 24816 -29162 24856 -29082
rect 24936 -29162 24976 -29082
rect 25056 -29162 25096 -29082
rect 25176 -29162 25216 -29082
rect 25296 -29162 25336 -29082
rect 25416 -29162 25456 -29082
rect 25536 -29162 25576 -29082
rect 25656 -29162 25696 -29082
rect 25776 -29162 25816 -29082
rect 25896 -29162 25936 -29082
rect 26016 -29162 26056 -29082
rect 26136 -29162 26176 -29082
rect 26256 -29162 26296 -29082
rect 26376 -29162 26416 -29082
rect 26496 -29162 26536 -29082
rect 26616 -29162 26656 -29082
rect 26736 -29162 26776 -29082
rect 26856 -29162 26896 -29082
rect 26976 -29162 27016 -29082
rect 27096 -29162 27136 -29082
rect 27216 -29162 27256 -29082
rect 27336 -29162 27376 -29082
rect 27456 -29162 27496 -29082
rect 27576 -29162 27616 -29082
rect 27696 -29162 27736 -29082
rect 27816 -29162 27856 -29082
rect 27936 -29162 27976 -29082
rect 28056 -29162 28096 -29082
rect 28176 -29162 28216 -29082
rect 28296 -29162 28336 -29082
rect 28416 -29162 28456 -29082
rect 28536 -29162 28576 -29082
rect 28656 -29162 28696 -29082
rect 28776 -29162 28816 -29082
rect 28896 -29162 28936 -29082
rect 29016 -29162 29056 -29082
rect 29136 -29162 29176 -29082
rect 29256 -29162 29296 -29082
rect 29376 -29162 29416 -29082
rect 29496 -29162 29536 -29082
rect 29616 -29162 29656 -29082
rect 29736 -29162 29776 -29082
rect 29856 -29162 29896 -29082
rect 29976 -29162 30016 -29082
rect 30096 -29162 30116 -29082
rect 23636 -29182 30116 -29162
rect 30596 -29042 30996 -29022
rect 30596 -29122 30616 -29042
rect 30696 -29122 30756 -29042
rect 30836 -29122 30896 -29042
rect 30976 -29122 30996 -29042
rect 30596 -29182 30996 -29122
rect 22796 -29262 22816 -29182
rect 22896 -29262 22956 -29182
rect 23036 -29262 23096 -29182
rect 23176 -29262 23196 -29182
rect 22796 -29322 23196 -29262
rect 22796 -29402 22816 -29322
rect 22896 -29402 22956 -29322
rect 23036 -29402 23096 -29322
rect 23176 -29402 23196 -29322
rect 22796 -29422 23196 -29402
rect 30596 -29262 30616 -29182
rect 30696 -29262 30756 -29182
rect 30836 -29262 30896 -29182
rect 30976 -29262 30996 -29182
rect 30596 -29322 30996 -29262
rect 30596 -29402 30616 -29322
rect 30696 -29402 30756 -29322
rect 30836 -29402 30896 -29322
rect 30976 -29402 30996 -29322
rect 30596 -29422 30996 -29402
rect 26696 -29642 27096 -29622
rect 26696 -29702 26716 -29642
rect 26776 -29702 26816 -29642
rect 26876 -29702 26916 -29642
rect 26976 -29702 27016 -29642
rect 27076 -29702 27096 -29642
rect 26696 -29742 27096 -29702
rect 26696 -29802 26716 -29742
rect 26776 -29802 26816 -29742
rect 26876 -29802 26916 -29742
rect 26976 -29802 27016 -29742
rect 27076 -29802 27096 -29742
rect 26696 -29842 27096 -29802
rect 26696 -29902 26716 -29842
rect 26776 -29902 26816 -29842
rect 26876 -29902 26916 -29842
rect 26976 -29902 27016 -29842
rect 27076 -29902 27096 -29842
rect 26696 -29942 27096 -29902
rect 26696 -30002 26716 -29942
rect 26776 -30002 26816 -29942
rect 26876 -30002 26916 -29942
rect 26976 -30002 27016 -29942
rect 27076 -30002 27096 -29942
rect 26696 -30022 27096 -30002
rect 21736 -30442 22136 -30422
rect 21736 -30502 21756 -30442
rect 21816 -30502 21856 -30442
rect 21916 -30502 21956 -30442
rect 22016 -30502 22056 -30442
rect 22116 -30502 22136 -30442
rect 21736 -30522 22136 -30502
rect 21736 -30582 21756 -30522
rect 21816 -30582 21856 -30522
rect 21916 -30582 21956 -30522
rect 22016 -30582 22056 -30522
rect 22116 -30582 22136 -30522
rect 21736 -30622 22136 -30582
rect 21736 -30682 21756 -30622
rect 21816 -30682 21856 -30622
rect 21916 -30682 21956 -30622
rect 22016 -30682 22056 -30622
rect 22116 -30682 22136 -30622
rect 21736 -30722 22136 -30682
rect 21736 -30782 21756 -30722
rect 21816 -30782 21856 -30722
rect 21916 -30782 21956 -30722
rect 22016 -30782 22056 -30722
rect 22116 -30782 22136 -30722
rect 21736 -30802 22136 -30782
rect 31656 -30442 32056 -30422
rect 31656 -30502 31676 -30442
rect 31736 -30502 31776 -30442
rect 31836 -30502 31876 -30442
rect 31936 -30502 31976 -30442
rect 32036 -30502 32056 -30442
rect 31656 -30522 32056 -30502
rect 31656 -30582 31676 -30522
rect 31736 -30582 31776 -30522
rect 31836 -30582 31876 -30522
rect 31936 -30582 31976 -30522
rect 32036 -30582 32056 -30522
rect 31656 -30622 32056 -30582
rect 31656 -30682 31676 -30622
rect 31736 -30682 31776 -30622
rect 31836 -30682 31876 -30622
rect 31936 -30682 31976 -30622
rect 32036 -30682 32056 -30622
rect 31656 -30722 32056 -30682
rect 31656 -30782 31676 -30722
rect 31736 -30782 31776 -30722
rect 31836 -30782 31876 -30722
rect 31936 -30782 31976 -30722
rect 32036 -30782 32056 -30722
rect 31656 -30802 32056 -30782
<< via1 >>
rect 20896 -21962 20914 -21902
rect 20914 -21962 20948 -21902
rect 20948 -21962 20956 -21902
rect 20896 -22142 20914 -22082
rect 20914 -22142 20948 -22082
rect 20948 -22142 20956 -22082
rect 21496 -21962 21530 -21902
rect 21530 -21962 21556 -21902
rect 21496 -22142 21530 -22082
rect 21530 -22142 21556 -22082
rect 22136 -21962 22146 -21902
rect 22146 -21962 22180 -21902
rect 22180 -21962 22196 -21902
rect 22136 -22142 22146 -22082
rect 22146 -22142 22180 -22082
rect 22180 -22142 22196 -22082
rect 22736 -21962 22762 -21902
rect 22762 -21962 22796 -21902
rect 22736 -22142 22762 -22082
rect 22762 -22142 22796 -22082
rect 24896 -21062 24956 -21002
rect 24996 -21062 24999 -21002
rect 24999 -21062 25056 -21002
rect 24896 -21142 24956 -21082
rect 24996 -21142 24999 -21082
rect 24999 -21142 25056 -21082
rect 24896 -21262 24956 -21202
rect 24996 -21262 24999 -21202
rect 24999 -21262 25056 -21202
rect 24896 -21342 24956 -21282
rect 24996 -21342 24999 -21282
rect 24999 -21342 25056 -21282
rect 26136 -21062 26196 -21002
rect 26136 -21142 26196 -21082
rect 26136 -21262 26196 -21202
rect 26136 -21342 26196 -21282
rect 26236 -21062 26296 -21002
rect 26236 -21142 26296 -21082
rect 26236 -21262 26296 -21202
rect 26236 -21342 26296 -21282
rect 27356 -21062 27416 -21002
rect 27456 -21062 27463 -21002
rect 27463 -21062 27516 -21002
rect 27356 -21142 27416 -21082
rect 27456 -21142 27463 -21082
rect 27463 -21142 27516 -21082
rect 27356 -21262 27416 -21202
rect 27456 -21262 27463 -21202
rect 27463 -21262 27516 -21202
rect 27356 -21342 27416 -21282
rect 27456 -21342 27463 -21282
rect 27463 -21342 27516 -21282
rect 28596 -21062 28656 -21002
rect 28596 -21142 28656 -21082
rect 28596 -21262 28656 -21202
rect 28596 -21342 28656 -21282
rect 28696 -21062 28756 -21002
rect 28696 -21142 28756 -21082
rect 28696 -21262 28756 -21202
rect 28696 -21342 28756 -21282
rect 23376 -21962 23378 -21902
rect 23378 -21962 23412 -21902
rect 23412 -21962 23436 -21902
rect 23376 -22142 23378 -22082
rect 23378 -22142 23412 -22082
rect 23412 -22142 23436 -22082
rect 24636 -22042 24716 -21962
rect 24756 -22042 24836 -21962
rect 24876 -22042 24956 -21962
rect 24996 -22042 25076 -21962
rect 25116 -22042 25196 -21962
rect 25236 -22042 25316 -21962
rect 25356 -22042 25436 -21962
rect 25476 -22042 25556 -21962
rect 25596 -22042 25676 -21962
rect 25716 -22042 25796 -21962
rect 25836 -22042 25916 -21962
rect 25956 -22042 26036 -21962
rect 26076 -22042 26156 -21962
rect 26196 -22042 26276 -21962
rect 26316 -22042 26396 -21962
rect 26436 -22042 26516 -21962
rect 26556 -22042 26636 -21962
rect 26676 -22042 26756 -21962
rect 26796 -22042 26876 -21962
rect 26916 -22042 26996 -21962
rect 27036 -22042 27116 -21962
rect 27156 -22042 27236 -21962
rect 27276 -22042 27356 -21962
rect 27396 -22042 27476 -21962
rect 27516 -22042 27596 -21962
rect 27636 -22042 27716 -21962
rect 27756 -22042 27836 -21962
rect 27876 -22042 27956 -21962
rect 27996 -22042 28076 -21962
rect 28116 -22042 28196 -21962
rect 28236 -22042 28316 -21962
rect 28356 -22042 28436 -21962
rect 28476 -22042 28556 -21962
rect 28596 -22042 28676 -21962
rect 28716 -22042 28796 -21962
rect 28836 -22042 28916 -21962
rect 28956 -22042 29036 -21962
rect 29076 -22042 29156 -21962
rect 24636 -22182 24716 -22102
rect 24756 -22182 24836 -22102
rect 24876 -22182 24956 -22102
rect 24996 -22182 25076 -22102
rect 25116 -22182 25196 -22102
rect 25236 -22182 25316 -22102
rect 25356 -22182 25436 -22102
rect 25476 -22182 25556 -22102
rect 25596 -22182 25676 -22102
rect 25716 -22182 25796 -22102
rect 25836 -22182 25916 -22102
rect 25956 -22182 26036 -22102
rect 26076 -22182 26156 -22102
rect 26196 -22182 26276 -22102
rect 26316 -22182 26396 -22102
rect 26436 -22182 26516 -22102
rect 26556 -22182 26636 -22102
rect 26676 -22182 26756 -22102
rect 26796 -22182 26876 -22102
rect 26916 -22182 26996 -22102
rect 27036 -22182 27116 -22102
rect 27156 -22182 27236 -22102
rect 27276 -22182 27356 -22102
rect 27396 -22182 27476 -22102
rect 27516 -22182 27596 -22102
rect 27636 -22182 27716 -22102
rect 27756 -22182 27836 -22102
rect 27876 -22182 27956 -22102
rect 27996 -22182 28076 -22102
rect 28116 -22182 28196 -22102
rect 28236 -22182 28316 -22102
rect 28356 -22182 28436 -22102
rect 28476 -22182 28556 -22102
rect 28596 -22182 28676 -22102
rect 28716 -22182 28796 -22102
rect 28836 -22182 28916 -22102
rect 28956 -22182 29036 -22102
rect 29076 -22182 29156 -22102
rect 30336 -21962 30354 -21902
rect 30354 -21962 30388 -21902
rect 30388 -21962 30396 -21902
rect 30336 -22142 30354 -22082
rect 30354 -22142 30388 -22082
rect 30388 -22142 30396 -22082
rect 30936 -21962 30970 -21902
rect 30970 -21962 30996 -21902
rect 30936 -22142 30970 -22082
rect 30970 -22142 30996 -22082
rect 31576 -21962 31586 -21902
rect 31586 -21962 31620 -21902
rect 31620 -21962 31636 -21902
rect 31576 -22142 31586 -22082
rect 31586 -22142 31620 -22082
rect 31620 -22142 31636 -22082
rect 32176 -21962 32202 -21902
rect 32202 -21962 32236 -21902
rect 32176 -22142 32202 -22082
rect 32202 -22142 32236 -22082
rect 32796 -21962 32818 -21902
rect 32818 -21962 32852 -21902
rect 32852 -21962 32856 -21902
rect 32796 -22142 32818 -22082
rect 32818 -22142 32852 -22082
rect 32852 -22142 32856 -22082
rect 24636 -22322 24716 -22242
rect 24756 -22322 24836 -22242
rect 24876 -22322 24956 -22242
rect 24996 -22322 25076 -22242
rect 25116 -22322 25196 -22242
rect 25236 -22322 25316 -22242
rect 25356 -22322 25436 -22242
rect 25476 -22322 25556 -22242
rect 25596 -22322 25676 -22242
rect 25716 -22322 25796 -22242
rect 25836 -22322 25916 -22242
rect 25956 -22322 26036 -22242
rect 26076 -22322 26156 -22242
rect 26196 -22322 26276 -22242
rect 26316 -22322 26396 -22242
rect 26436 -22322 26516 -22242
rect 26556 -22322 26636 -22242
rect 26676 -22322 26756 -22242
rect 26796 -22322 26876 -22242
rect 26916 -22322 26996 -22242
rect 27036 -22322 27116 -22242
rect 27156 -22322 27236 -22242
rect 27276 -22322 27356 -22242
rect 27396 -22322 27476 -22242
rect 27516 -22322 27596 -22242
rect 27636 -22322 27716 -22242
rect 27756 -22322 27836 -22242
rect 27876 -22322 27956 -22242
rect 27996 -22322 28076 -22242
rect 28116 -22322 28196 -22242
rect 28236 -22322 28316 -22242
rect 28356 -22322 28436 -22242
rect 28476 -22322 28556 -22242
rect 28596 -22322 28676 -22242
rect 28716 -22322 28796 -22242
rect 28836 -22322 28916 -22242
rect 28956 -22322 29036 -22242
rect 29076 -22322 29156 -22242
rect 20976 -22522 21056 -22442
rect 21076 -22522 21156 -22442
rect 21176 -22522 21256 -22442
rect 21276 -22522 21356 -22442
rect 21376 -22522 21456 -22442
rect 21476 -22522 21556 -22442
rect 21576 -22522 21656 -22442
rect 21676 -22522 21756 -22442
rect 21776 -22522 21856 -22442
rect 21876 -22522 21956 -22442
rect 21976 -22522 22056 -22442
rect 22076 -22522 22156 -22442
rect 22176 -22522 22256 -22442
rect 22276 -22522 22356 -22442
rect 22376 -22522 22456 -22442
rect 22476 -22522 22556 -22442
rect 22576 -22522 22656 -22442
rect 22676 -22522 22756 -22442
rect 22776 -22522 22856 -22442
rect 22876 -22522 22956 -22442
rect 22976 -22522 23056 -22442
rect 23076 -22522 23156 -22442
rect 23176 -22522 23256 -22442
rect 23276 -22522 23356 -22442
rect 20976 -22662 21056 -22582
rect 21076 -22662 21156 -22582
rect 21176 -22662 21256 -22582
rect 21276 -22662 21356 -22582
rect 21376 -22662 21456 -22582
rect 21476 -22662 21556 -22582
rect 21576 -22662 21656 -22582
rect 21676 -22662 21756 -22582
rect 21776 -22662 21856 -22582
rect 21876 -22662 21956 -22582
rect 21976 -22662 22056 -22582
rect 22076 -22662 22156 -22582
rect 22176 -22662 22256 -22582
rect 22276 -22662 22356 -22582
rect 22376 -22662 22456 -22582
rect 22476 -22662 22556 -22582
rect 22576 -22662 22656 -22582
rect 22676 -22662 22756 -22582
rect 22776 -22662 22856 -22582
rect 22876 -22662 22956 -22582
rect 22976 -22662 23056 -22582
rect 23076 -22662 23156 -22582
rect 23176 -22662 23256 -22582
rect 23276 -22662 23356 -22582
rect 20976 -22802 21056 -22722
rect 21076 -22802 21156 -22722
rect 21176 -22802 21256 -22722
rect 21276 -22802 21356 -22722
rect 21376 -22802 21456 -22722
rect 21476 -22802 21556 -22722
rect 21576 -22802 21656 -22722
rect 21676 -22802 21756 -22722
rect 21776 -22802 21856 -22722
rect 21876 -22802 21956 -22722
rect 21976 -22802 22056 -22722
rect 22076 -22802 22156 -22722
rect 22176 -22802 22256 -22722
rect 22276 -22802 22356 -22722
rect 22376 -22802 22456 -22722
rect 22476 -22802 22556 -22722
rect 22576 -22802 22656 -22722
rect 22676 -22802 22756 -22722
rect 22776 -22802 22856 -22722
rect 22876 -22802 22956 -22722
rect 22976 -22802 23056 -22722
rect 23076 -22802 23156 -22722
rect 23176 -22802 23256 -22722
rect 23276 -22802 23356 -22722
rect 30416 -22522 30496 -22442
rect 30516 -22522 30596 -22442
rect 30616 -22522 30696 -22442
rect 30716 -22522 30796 -22442
rect 30816 -22522 30896 -22442
rect 30916 -22522 30996 -22442
rect 31016 -22522 31096 -22442
rect 31116 -22522 31196 -22442
rect 31216 -22522 31296 -22442
rect 31316 -22522 31396 -22442
rect 31416 -22522 31496 -22442
rect 31516 -22522 31596 -22442
rect 31616 -22522 31696 -22442
rect 31716 -22522 31796 -22442
rect 31816 -22522 31896 -22442
rect 31916 -22522 31996 -22442
rect 32016 -22522 32096 -22442
rect 32116 -22522 32196 -22442
rect 32216 -22522 32296 -22442
rect 32316 -22522 32396 -22442
rect 32416 -22522 32496 -22442
rect 32516 -22522 32596 -22442
rect 32616 -22522 32696 -22442
rect 32716 -22522 32796 -22442
rect 30416 -22662 30496 -22582
rect 30516 -22662 30596 -22582
rect 30616 -22662 30696 -22582
rect 30716 -22662 30796 -22582
rect 30816 -22662 30896 -22582
rect 30916 -22662 30996 -22582
rect 31016 -22662 31096 -22582
rect 31116 -22662 31196 -22582
rect 31216 -22662 31296 -22582
rect 31316 -22662 31396 -22582
rect 31416 -22662 31496 -22582
rect 31516 -22662 31596 -22582
rect 31616 -22662 31696 -22582
rect 31716 -22662 31796 -22582
rect 31816 -22662 31896 -22582
rect 31916 -22662 31996 -22582
rect 32016 -22662 32096 -22582
rect 32116 -22662 32196 -22582
rect 32216 -22662 32296 -22582
rect 32316 -22662 32396 -22582
rect 32416 -22662 32496 -22582
rect 32516 -22662 32596 -22582
rect 32616 -22662 32696 -22582
rect 32716 -22662 32796 -22582
rect 30416 -22802 30496 -22722
rect 30516 -22802 30596 -22722
rect 30616 -22802 30696 -22722
rect 30716 -22802 30796 -22722
rect 30816 -22802 30896 -22722
rect 30916 -22802 30996 -22722
rect 31016 -22802 31096 -22722
rect 31116 -22802 31196 -22722
rect 31216 -22802 31296 -22722
rect 31316 -22802 31396 -22722
rect 31416 -22802 31496 -22722
rect 31516 -22802 31596 -22722
rect 31616 -22802 31696 -22722
rect 31716 -22802 31796 -22722
rect 31816 -22802 31896 -22722
rect 31916 -22802 31996 -22722
rect 32016 -22802 32096 -22722
rect 32116 -22802 32196 -22722
rect 32216 -22802 32296 -22722
rect 32316 -22802 32396 -22722
rect 32416 -22802 32496 -22722
rect 32516 -22802 32596 -22722
rect 32616 -22802 32696 -22722
rect 32716 -22802 32796 -22722
rect 21856 -23042 21874 -22982
rect 21874 -23042 21908 -22982
rect 21908 -23042 21916 -22982
rect 21856 -23222 21874 -23162
rect 21874 -23222 21908 -23162
rect 21908 -23222 21916 -23162
rect 22316 -23042 22350 -22982
rect 22350 -23042 22376 -22982
rect 22316 -23222 22350 -23162
rect 22350 -23222 22376 -23162
rect 22116 -23522 22146 -23462
rect 22146 -23522 22176 -23462
rect 22116 -23622 22146 -23562
rect 22146 -23622 22176 -23562
rect 26716 -23002 26796 -22922
rect 26856 -23002 26936 -22922
rect 26996 -23002 27076 -22922
rect 23796 -23522 23808 -23462
rect 23808 -23522 23842 -23462
rect 23842 -23522 23856 -23462
rect 23796 -23602 23808 -23542
rect 23808 -23602 23842 -23542
rect 23842 -23602 23856 -23542
rect 23796 -23682 23808 -23622
rect 23808 -23682 23842 -23622
rect 23842 -23682 23856 -23622
rect 24116 -23522 24124 -23462
rect 24124 -23522 24158 -23462
rect 24158 -23522 24176 -23462
rect 24116 -23602 24124 -23542
rect 24124 -23602 24158 -23542
rect 24158 -23602 24176 -23542
rect 24116 -23682 24124 -23622
rect 24124 -23682 24158 -23622
rect 24158 -23682 24176 -23622
rect 26716 -23122 26796 -23042
rect 26856 -23122 26936 -23042
rect 26996 -23122 27076 -23042
rect 25596 -23522 25608 -23462
rect 25608 -23522 25642 -23462
rect 25642 -23522 25656 -23462
rect 25596 -23602 25608 -23542
rect 25608 -23602 25642 -23542
rect 25642 -23602 25656 -23542
rect 25596 -23682 25608 -23622
rect 25608 -23682 25642 -23622
rect 25642 -23682 25656 -23622
rect 25916 -23522 25924 -23462
rect 25924 -23522 25958 -23462
rect 25958 -23522 25976 -23462
rect 25916 -23602 25924 -23542
rect 25924 -23602 25958 -23542
rect 25958 -23602 25976 -23542
rect 25916 -23682 25924 -23622
rect 25924 -23682 25958 -23622
rect 25958 -23682 25976 -23622
rect 26716 -23242 26796 -23162
rect 26856 -23242 26936 -23162
rect 26996 -23242 27076 -23162
rect 26716 -23362 26796 -23282
rect 26856 -23362 26936 -23282
rect 26996 -23362 27076 -23282
rect 26716 -23482 26796 -23402
rect 26856 -23482 26936 -23402
rect 26996 -23482 27076 -23402
rect 26716 -23602 26796 -23522
rect 26856 -23602 26936 -23522
rect 26996 -23602 27076 -23522
rect 26716 -23722 26796 -23642
rect 26856 -23722 26936 -23642
rect 26996 -23722 27076 -23642
rect 26716 -23842 26796 -23762
rect 26856 -23842 26936 -23762
rect 26996 -23842 27076 -23762
rect 26716 -23962 26796 -23882
rect 26856 -23962 26936 -23882
rect 26996 -23962 27076 -23882
rect 26716 -24082 26796 -24002
rect 26856 -24082 26936 -24002
rect 26996 -24082 27076 -24002
rect 27796 -23522 27808 -23462
rect 27808 -23522 27842 -23462
rect 27842 -23522 27856 -23462
rect 27796 -23602 27808 -23542
rect 27808 -23602 27842 -23542
rect 27842 -23602 27856 -23542
rect 27796 -23682 27808 -23622
rect 27808 -23682 27842 -23622
rect 27842 -23682 27856 -23622
rect 28116 -23522 28124 -23462
rect 28124 -23522 28158 -23462
rect 28158 -23522 28176 -23462
rect 28116 -23602 28124 -23542
rect 28124 -23602 28158 -23542
rect 28158 -23602 28176 -23542
rect 28116 -23682 28124 -23622
rect 28124 -23682 28158 -23622
rect 28158 -23682 28176 -23622
rect 29596 -23522 29608 -23462
rect 29608 -23522 29642 -23462
rect 29642 -23522 29656 -23462
rect 29596 -23602 29608 -23542
rect 29608 -23602 29642 -23542
rect 29642 -23602 29656 -23542
rect 29596 -23682 29608 -23622
rect 29608 -23682 29642 -23622
rect 29642 -23682 29656 -23622
rect 29916 -23522 29924 -23462
rect 29924 -23522 29958 -23462
rect 29958 -23522 29976 -23462
rect 29916 -23602 29924 -23542
rect 29924 -23602 29958 -23542
rect 29958 -23602 29976 -23542
rect 29916 -23682 29924 -23622
rect 29924 -23682 29958 -23622
rect 29958 -23682 29976 -23622
rect 31456 -23042 31488 -22982
rect 31488 -23042 31516 -22982
rect 31456 -23222 31488 -23162
rect 31488 -23222 31516 -23162
rect 31916 -23042 31930 -22982
rect 31930 -23042 31964 -22982
rect 31964 -23042 31976 -22982
rect 31916 -23222 31930 -23162
rect 31930 -23222 31964 -23162
rect 31964 -23222 31976 -23162
rect 31636 -23522 31692 -23462
rect 31692 -23522 31696 -23462
rect 31636 -23622 31692 -23562
rect 31692 -23622 31696 -23562
rect 23876 -24166 23936 -24142
rect 24036 -24166 24096 -24142
rect 23876 -24202 23936 -24166
rect 24036 -24202 24096 -24166
rect 25676 -24166 25736 -24142
rect 25836 -24166 25896 -24142
rect 25676 -24202 25736 -24166
rect 25836 -24202 25896 -24166
rect 26716 -24202 26796 -24122
rect 26856 -24202 26936 -24122
rect 26996 -24202 27076 -24122
rect 27876 -24166 27936 -24142
rect 28036 -24166 28096 -24142
rect 26716 -24322 26796 -24242
rect 26856 -24322 26936 -24242
rect 26996 -24322 27076 -24242
rect 27876 -24202 27936 -24166
rect 28036 -24202 28096 -24166
rect 29676 -24166 29736 -24142
rect 29836 -24166 29896 -24142
rect 29676 -24202 29736 -24166
rect 29836 -24202 29896 -24166
rect 26716 -24442 26796 -24362
rect 26856 -24442 26936 -24362
rect 26996 -24442 27076 -24362
rect 26716 -24562 26796 -24482
rect 26856 -24562 26936 -24482
rect 26996 -24562 27076 -24482
rect 21416 -25042 21428 -24982
rect 21428 -25042 21462 -24982
rect 21462 -25042 21476 -24982
rect 21416 -25222 21428 -25162
rect 21428 -25222 21462 -25162
rect 21462 -25222 21476 -25162
rect 22036 -25042 22044 -24982
rect 22044 -25042 22078 -24982
rect 22078 -25042 22096 -24982
rect 22036 -25222 22044 -25162
rect 22044 -25222 22078 -25162
rect 22078 -25222 22096 -25162
rect 23876 -24774 23936 -24742
rect 24036 -24774 24096 -24742
rect 23876 -24802 23936 -24774
rect 24036 -24802 24096 -24774
rect 25676 -24774 25736 -24742
rect 25836 -24774 25896 -24742
rect 25676 -24802 25736 -24774
rect 25836 -24802 25896 -24774
rect 26716 -24682 26796 -24602
rect 26856 -24682 26936 -24602
rect 26996 -24682 27076 -24602
rect 26716 -24802 26796 -24722
rect 26856 -24802 26936 -24722
rect 26996 -24802 27076 -24722
rect 22636 -25042 22660 -24982
rect 22660 -25042 22694 -24982
rect 22694 -25042 22696 -24982
rect 22636 -25222 22660 -25162
rect 22660 -25222 22694 -25162
rect 22694 -25222 22696 -25162
rect 23796 -25022 23808 -24962
rect 23808 -25022 23842 -24962
rect 23842 -25022 23856 -24962
rect 23796 -25102 23808 -25042
rect 23808 -25102 23842 -25042
rect 23842 -25102 23856 -25042
rect 23796 -25182 23808 -25122
rect 23808 -25182 23842 -25122
rect 23842 -25182 23856 -25122
rect 24116 -25022 24124 -24962
rect 24124 -25022 24158 -24962
rect 24158 -25022 24176 -24962
rect 24116 -25102 24124 -25042
rect 24124 -25102 24158 -25042
rect 24158 -25102 24176 -25042
rect 24116 -25182 24124 -25122
rect 24124 -25182 24158 -25122
rect 24158 -25182 24176 -25122
rect 27876 -24774 27936 -24742
rect 28036 -24774 28096 -24742
rect 27876 -24802 27936 -24774
rect 28036 -24802 28096 -24774
rect 25596 -25622 25608 -25562
rect 25608 -25622 25642 -25562
rect 25642 -25622 25656 -25562
rect 25596 -25702 25608 -25642
rect 25608 -25702 25642 -25642
rect 25642 -25702 25656 -25642
rect 25596 -25782 25608 -25722
rect 25608 -25782 25642 -25722
rect 25642 -25782 25656 -25722
rect 25916 -25622 25924 -25562
rect 25924 -25622 25958 -25562
rect 25958 -25622 25976 -25562
rect 25916 -25702 25924 -25642
rect 25924 -25702 25958 -25642
rect 25958 -25702 25976 -25642
rect 25916 -25782 25924 -25722
rect 25924 -25782 25958 -25722
rect 25958 -25782 25976 -25722
rect 26716 -24922 26796 -24842
rect 26856 -24922 26936 -24842
rect 26996 -24922 27076 -24842
rect 29676 -24774 29736 -24742
rect 29836 -24774 29896 -24742
rect 29676 -24802 29736 -24774
rect 29836 -24802 29896 -24774
rect 26716 -25042 26796 -24962
rect 26856 -25042 26936 -24962
rect 26996 -25042 27076 -24962
rect 26716 -25162 26796 -25082
rect 26856 -25162 26936 -25082
rect 26996 -25162 27076 -25082
rect 26716 -25282 26796 -25202
rect 26856 -25282 26936 -25202
rect 26996 -25282 27076 -25202
rect 26716 -25402 26796 -25322
rect 26856 -25402 26936 -25322
rect 26996 -25402 27076 -25322
rect 26716 -25522 26796 -25442
rect 26856 -25522 26936 -25442
rect 26996 -25522 27076 -25442
rect 26716 -25642 26796 -25562
rect 26856 -25642 26936 -25562
rect 26996 -25642 27076 -25562
rect 26716 -25762 26796 -25682
rect 26856 -25762 26936 -25682
rect 26996 -25762 27076 -25682
rect 27796 -25622 27808 -25562
rect 27808 -25622 27842 -25562
rect 27842 -25622 27856 -25562
rect 27796 -25702 27808 -25642
rect 27808 -25702 27842 -25642
rect 27842 -25702 27856 -25642
rect 27796 -25782 27808 -25722
rect 27808 -25782 27842 -25722
rect 27842 -25782 27856 -25722
rect 26716 -25882 26796 -25802
rect 26856 -25882 26936 -25802
rect 26996 -25882 27076 -25802
rect 26716 -26002 26796 -25922
rect 26856 -26002 26936 -25922
rect 26996 -26002 27076 -25922
rect 28116 -25622 28124 -25562
rect 28124 -25622 28158 -25562
rect 28158 -25622 28176 -25562
rect 28116 -25702 28124 -25642
rect 28124 -25702 28158 -25642
rect 28158 -25702 28176 -25642
rect 28116 -25782 28124 -25722
rect 28124 -25782 28158 -25722
rect 28158 -25782 28176 -25722
rect 29596 -25022 29608 -24962
rect 29608 -25022 29642 -24962
rect 29642 -25022 29656 -24962
rect 29596 -25102 29608 -25042
rect 29608 -25102 29642 -25042
rect 29642 -25102 29656 -25042
rect 29596 -25182 29608 -25122
rect 29608 -25182 29642 -25122
rect 29642 -25182 29656 -25122
rect 29916 -25022 29924 -24962
rect 29924 -25022 29958 -24962
rect 29958 -25022 29976 -24962
rect 29916 -25102 29924 -25042
rect 29924 -25102 29958 -25042
rect 29958 -25102 29976 -25042
rect 29916 -25182 29924 -25122
rect 29924 -25182 29958 -25122
rect 29958 -25182 29976 -25122
rect 31076 -25042 31088 -24982
rect 31088 -25042 31122 -24982
rect 31122 -25042 31136 -24982
rect 31076 -25222 31088 -25162
rect 31088 -25222 31122 -25162
rect 31122 -25222 31136 -25162
rect 31696 -25042 31704 -24982
rect 31704 -25042 31738 -24982
rect 31738 -25042 31756 -24982
rect 31696 -25222 31704 -25162
rect 31704 -25222 31738 -25162
rect 31738 -25222 31756 -25162
rect 32296 -25042 32320 -24982
rect 32320 -25042 32354 -24982
rect 32354 -25042 32356 -24982
rect 32296 -25222 32320 -25162
rect 32320 -25222 32354 -25162
rect 32354 -25222 32356 -25162
rect 21496 -26562 21556 -26502
rect 21576 -26562 21636 -26502
rect 21656 -26562 21716 -26502
rect 21736 -26562 21796 -26502
rect 21816 -26562 21876 -26502
rect 21896 -26562 21956 -26502
rect 21976 -26562 22036 -26502
rect 22056 -26562 22116 -26502
rect 22136 -26562 22196 -26502
rect 22216 -26562 22276 -26502
rect 22296 -26562 22356 -26502
rect 22376 -26562 22436 -26502
rect 22456 -26562 22556 -26502
rect 22576 -26562 22636 -26502
rect 21496 -26662 21556 -26602
rect 21576 -26662 21636 -26602
rect 21656 -26662 21716 -26602
rect 21736 -26662 21796 -26602
rect 21816 -26662 21876 -26602
rect 21896 -26662 21956 -26602
rect 21976 -26662 22036 -26602
rect 22056 -26662 22116 -26602
rect 22136 -26662 22196 -26602
rect 22216 -26662 22276 -26602
rect 22296 -26662 22356 -26602
rect 22376 -26662 22436 -26602
rect 22456 -26662 22556 -26602
rect 22576 -26662 22636 -26602
rect 24376 -26562 24388 -26502
rect 24388 -26562 24422 -26502
rect 24422 -26562 24436 -26502
rect 24476 -26562 24536 -26502
rect 24376 -26642 24388 -26582
rect 24388 -26642 24422 -26582
rect 24422 -26642 24436 -26582
rect 24476 -26642 24536 -26582
rect 24376 -26822 24388 -26762
rect 24388 -26822 24422 -26762
rect 24422 -26822 24436 -26762
rect 24476 -26822 24536 -26762
rect 24376 -26902 24388 -26842
rect 24388 -26902 24422 -26842
rect 24422 -26902 24436 -26842
rect 24476 -26902 24536 -26842
rect 24376 -27182 24388 -27122
rect 24388 -27182 24422 -27122
rect 24422 -27182 24436 -27122
rect 24476 -27182 24536 -27122
rect 24376 -27262 24388 -27202
rect 24388 -27262 24422 -27202
rect 24422 -27262 24436 -27202
rect 24476 -27262 24536 -27202
rect 24376 -27402 24388 -27342
rect 24388 -27402 24422 -27342
rect 24422 -27402 24436 -27342
rect 24476 -27402 24536 -27342
rect 24376 -27482 24388 -27422
rect 24388 -27482 24422 -27422
rect 24422 -27482 24436 -27422
rect 24476 -27482 24536 -27422
rect 24956 -26582 25004 -26522
rect 25004 -26582 25016 -26522
rect 25036 -26582 25038 -26522
rect 25038 -26582 25096 -26522
rect 24956 -26662 25004 -26602
rect 25004 -26662 25016 -26602
rect 25036 -26662 25038 -26602
rect 25038 -26662 25096 -26602
rect 24956 -26742 25004 -26682
rect 25004 -26742 25016 -26682
rect 25036 -26742 25038 -26682
rect 25038 -26742 25096 -26682
rect 24956 -26822 25004 -26762
rect 25004 -26822 25016 -26762
rect 25036 -26822 25038 -26762
rect 25038 -26822 25096 -26762
rect 24956 -26902 25004 -26842
rect 25004 -26902 25016 -26842
rect 25036 -26902 25038 -26842
rect 25038 -26902 25096 -26842
rect 25556 -27182 25616 -27122
rect 25556 -27262 25616 -27202
rect 25556 -27402 25616 -27342
rect 25556 -27482 25616 -27422
rect 25656 -27182 25716 -27122
rect 25656 -27262 25716 -27202
rect 25656 -27402 25716 -27342
rect 25656 -27482 25716 -27422
rect 26176 -26582 26236 -26522
rect 26256 -26582 26270 -26522
rect 26270 -26582 26316 -26522
rect 26176 -26662 26236 -26602
rect 26256 -26662 26270 -26602
rect 26270 -26662 26316 -26602
rect 26176 -26742 26236 -26682
rect 26256 -26742 26270 -26682
rect 26270 -26742 26316 -26682
rect 26176 -26822 26236 -26762
rect 26256 -26822 26270 -26762
rect 26270 -26822 26316 -26762
rect 26176 -26902 26236 -26842
rect 26256 -26902 26270 -26842
rect 26270 -26902 26316 -26842
rect 26796 -27182 26852 -27122
rect 26852 -27182 26856 -27122
rect 26896 -27182 26956 -27122
rect 26796 -27262 26852 -27202
rect 26852 -27262 26856 -27202
rect 26896 -27262 26956 -27202
rect 26796 -27402 26852 -27342
rect 26852 -27402 26856 -27342
rect 26896 -27402 26956 -27342
rect 26796 -27482 26852 -27422
rect 26852 -27482 26856 -27422
rect 26896 -27482 26956 -27422
rect 27416 -26582 27468 -26522
rect 27468 -26582 27476 -26522
rect 27496 -26582 27502 -26522
rect 27502 -26582 27556 -26522
rect 27416 -26662 27468 -26602
rect 27468 -26662 27476 -26602
rect 27496 -26662 27502 -26602
rect 27502 -26662 27556 -26602
rect 27416 -26742 27468 -26682
rect 27468 -26742 27476 -26682
rect 27496 -26742 27502 -26682
rect 27502 -26742 27556 -26682
rect 27416 -26822 27468 -26762
rect 27468 -26822 27476 -26762
rect 27496 -26822 27502 -26762
rect 27502 -26822 27556 -26762
rect 27416 -26902 27468 -26842
rect 27468 -26902 27476 -26842
rect 27496 -26902 27502 -26842
rect 27502 -26902 27556 -26842
rect 28016 -27182 28076 -27122
rect 28116 -27182 28118 -27122
rect 28118 -27182 28176 -27122
rect 28016 -27262 28076 -27202
rect 28116 -27262 28118 -27202
rect 28118 -27262 28176 -27202
rect 28016 -27402 28076 -27342
rect 28116 -27402 28118 -27342
rect 28118 -27402 28176 -27342
rect 28016 -27482 28076 -27422
rect 28116 -27482 28118 -27422
rect 28118 -27482 28176 -27422
rect 28636 -26582 28696 -26522
rect 28716 -26582 28734 -26522
rect 28734 -26582 28776 -26522
rect 28636 -26662 28696 -26602
rect 28716 -26662 28734 -26602
rect 28734 -26662 28776 -26602
rect 28636 -26742 28696 -26682
rect 28716 -26742 28734 -26682
rect 28734 -26742 28776 -26682
rect 28636 -26822 28696 -26762
rect 28716 -26822 28734 -26762
rect 28734 -26822 28776 -26762
rect 28636 -26902 28696 -26842
rect 28716 -26902 28734 -26842
rect 28734 -26902 28776 -26842
rect 29216 -26562 29276 -26502
rect 29316 -26562 29350 -26502
rect 29350 -26562 29376 -26502
rect 29216 -26642 29276 -26582
rect 29316 -26642 29350 -26582
rect 29350 -26642 29376 -26582
rect 29216 -26822 29276 -26762
rect 29316 -26822 29350 -26762
rect 29350 -26822 29376 -26762
rect 29216 -26902 29276 -26842
rect 29316 -26902 29350 -26842
rect 29350 -26902 29376 -26842
rect 29216 -27182 29276 -27122
rect 29316 -27182 29350 -27122
rect 29350 -27182 29376 -27122
rect 29216 -27262 29276 -27202
rect 29316 -27262 29350 -27202
rect 29350 -27262 29376 -27202
rect 29216 -27402 29276 -27342
rect 29316 -27402 29350 -27342
rect 29350 -27402 29376 -27342
rect 29216 -27482 29276 -27422
rect 29316 -27482 29350 -27422
rect 29350 -27482 29376 -27422
rect 31156 -26562 31216 -26502
rect 31236 -26562 31336 -26502
rect 31356 -26562 31416 -26502
rect 31436 -26562 31496 -26502
rect 31516 -26562 31576 -26502
rect 31596 -26562 31656 -26502
rect 31676 -26562 31736 -26502
rect 31756 -26562 31816 -26502
rect 31836 -26562 31896 -26502
rect 31916 -26562 31976 -26502
rect 31996 -26562 32056 -26502
rect 32076 -26562 32136 -26502
rect 32156 -26562 32216 -26502
rect 32236 -26562 32296 -26502
rect 31156 -26662 31216 -26602
rect 31236 -26662 31336 -26602
rect 31356 -26662 31416 -26602
rect 31436 -26662 31496 -26602
rect 31516 -26662 31576 -26602
rect 31596 -26662 31656 -26602
rect 31676 -26662 31736 -26602
rect 31756 -26662 31816 -26602
rect 31836 -26662 31896 -26602
rect 31916 -26662 31976 -26602
rect 31996 -26662 32056 -26602
rect 32076 -26662 32136 -26602
rect 32156 -26662 32216 -26602
rect 32236 -26662 32296 -26602
rect 22816 -29122 22896 -29042
rect 22956 -29122 23036 -29042
rect 23096 -29122 23176 -29042
rect 30616 -29122 30696 -29042
rect 30756 -29122 30836 -29042
rect 30896 -29122 30976 -29042
rect 22816 -29262 22896 -29182
rect 22956 -29262 23036 -29182
rect 23096 -29262 23176 -29182
rect 22816 -29402 22896 -29322
rect 22956 -29402 23036 -29322
rect 23096 -29402 23176 -29322
rect 30616 -29262 30696 -29182
rect 30756 -29262 30836 -29182
rect 30896 -29262 30976 -29182
rect 30616 -29402 30696 -29322
rect 30756 -29402 30836 -29322
rect 30896 -29402 30976 -29322
rect 26716 -29702 26776 -29642
rect 26816 -29702 26876 -29642
rect 26916 -29702 26976 -29642
rect 27016 -29702 27076 -29642
rect 26716 -29802 26776 -29742
rect 26816 -29802 26876 -29742
rect 26916 -29802 26976 -29742
rect 27016 -29802 27076 -29742
rect 26716 -29902 26776 -29842
rect 26816 -29902 26876 -29842
rect 26916 -29902 26976 -29842
rect 27016 -29902 27076 -29842
rect 26716 -30002 26776 -29942
rect 26816 -30002 26876 -29942
rect 26916 -30002 26976 -29942
rect 27016 -30002 27076 -29942
rect 21756 -30502 21816 -30442
rect 21856 -30502 21916 -30442
rect 21956 -30502 22016 -30442
rect 22056 -30502 22116 -30442
rect 21756 -30582 21816 -30522
rect 21856 -30582 21916 -30522
rect 21956 -30582 22016 -30522
rect 22056 -30582 22116 -30522
rect 21756 -30682 21816 -30622
rect 21856 -30682 21916 -30622
rect 21956 -30682 22016 -30622
rect 22056 -30682 22116 -30622
rect 21756 -30782 21816 -30722
rect 21856 -30782 21916 -30722
rect 21956 -30782 22016 -30722
rect 22056 -30782 22116 -30722
rect 31676 -30502 31736 -30442
rect 31776 -30502 31836 -30442
rect 31876 -30502 31936 -30442
rect 31976 -30502 32036 -30442
rect 31676 -30582 31736 -30522
rect 31776 -30582 31836 -30522
rect 31876 -30582 31936 -30522
rect 31976 -30582 32036 -30522
rect 31676 -30682 31736 -30622
rect 31776 -30682 31836 -30622
rect 31876 -30682 31936 -30622
rect 31976 -30682 32036 -30622
rect 31676 -30782 31736 -30722
rect 31776 -30782 31836 -30722
rect 31876 -30782 31936 -30722
rect 31976 -30782 32036 -30722
<< metal2 >>
rect 24816 -21002 28836 -20982
rect 24816 -21062 24896 -21002
rect 24956 -21062 24996 -21002
rect 25056 -21062 26136 -21002
rect 26196 -21062 26236 -21002
rect 26296 -21062 26716 -21002
rect 24816 -21082 26716 -21062
rect 26796 -21082 26856 -21002
rect 26936 -21082 26996 -21002
rect 27076 -21062 27356 -21002
rect 27416 -21062 27456 -21002
rect 27516 -21062 28596 -21002
rect 28656 -21062 28696 -21002
rect 28756 -21062 28836 -21002
rect 27076 -21082 28836 -21062
rect 24816 -21142 24896 -21082
rect 24956 -21142 24996 -21082
rect 25056 -21142 26136 -21082
rect 26196 -21142 26236 -21082
rect 26296 -21122 27356 -21082
rect 26296 -21142 26716 -21122
rect 24816 -21202 26716 -21142
rect 26796 -21202 26856 -21122
rect 26936 -21202 26996 -21122
rect 27076 -21142 27356 -21122
rect 27416 -21142 27456 -21082
rect 27516 -21142 28596 -21082
rect 28656 -21142 28696 -21082
rect 28756 -21142 28836 -21082
rect 27076 -21202 28836 -21142
rect 24816 -21262 24896 -21202
rect 24956 -21262 24996 -21202
rect 25056 -21262 26136 -21202
rect 26196 -21262 26236 -21202
rect 26296 -21262 27356 -21202
rect 27416 -21262 27456 -21202
rect 27516 -21262 28596 -21202
rect 28656 -21262 28696 -21202
rect 28756 -21262 28836 -21202
rect 24816 -21282 26716 -21262
rect 24816 -21342 24896 -21282
rect 24956 -21342 24996 -21282
rect 25056 -21342 26136 -21282
rect 26196 -21342 26236 -21282
rect 26296 -21342 26716 -21282
rect 26796 -21342 26856 -21262
rect 26936 -21342 26996 -21262
rect 27076 -21282 28836 -21262
rect 27076 -21342 27356 -21282
rect 27416 -21342 27456 -21282
rect 27516 -21342 28596 -21282
rect 28656 -21342 28696 -21282
rect 28756 -21342 28836 -21282
rect 24816 -21362 28836 -21342
rect 20856 -21902 23636 -21882
rect 20856 -21962 20896 -21902
rect 20956 -21962 21496 -21902
rect 21556 -21962 21776 -21902
rect 21836 -21962 21896 -21902
rect 21976 -21962 22036 -21902
rect 22096 -21962 22136 -21902
rect 22196 -21962 22736 -21902
rect 22796 -21962 23376 -21902
rect 23436 -21962 23636 -21902
rect 30136 -21902 32916 -21882
rect 20856 -22082 23636 -21962
rect 20856 -22142 20896 -22082
rect 20956 -22142 21496 -22082
rect 21556 -22142 21776 -22082
rect 21836 -22142 21896 -22082
rect 21976 -22142 22036 -22082
rect 22096 -22142 22136 -22082
rect 22196 -22142 22736 -22082
rect 22796 -22142 23376 -22082
rect 23436 -22142 23636 -22082
rect 20856 -22162 23636 -22142
rect 23816 -21962 29956 -21942
rect 23816 -22042 24236 -21962
rect 24316 -22042 24376 -21962
rect 24456 -22042 24516 -21962
rect 24596 -22042 24636 -21962
rect 24716 -22042 24756 -21962
rect 24836 -22042 24876 -21962
rect 24956 -22042 24996 -21962
rect 25076 -22042 25116 -21962
rect 25196 -22042 25236 -21962
rect 25316 -22042 25356 -21962
rect 25436 -22042 25476 -21962
rect 25556 -22042 25596 -21962
rect 25676 -22042 25716 -21962
rect 25796 -22042 25836 -21962
rect 25916 -22042 25956 -21962
rect 26036 -22042 26076 -21962
rect 26156 -22042 26196 -21962
rect 26276 -22042 26316 -21962
rect 26396 -22042 26436 -21962
rect 26516 -22042 26556 -21962
rect 26636 -22042 26676 -21962
rect 26756 -22042 26796 -21962
rect 26876 -22042 26916 -21962
rect 26996 -22042 27036 -21962
rect 27116 -22042 27156 -21962
rect 27236 -22042 27276 -21962
rect 27356 -22042 27396 -21962
rect 27476 -22042 27516 -21962
rect 27596 -22042 27636 -21962
rect 27716 -22042 27756 -21962
rect 27836 -22042 27876 -21962
rect 27956 -22042 27996 -21962
rect 28076 -22042 28116 -21962
rect 28196 -22042 28236 -21962
rect 28316 -22042 28356 -21962
rect 28436 -22042 28476 -21962
rect 28556 -22042 28596 -21962
rect 28676 -22042 28716 -21962
rect 28796 -22042 28836 -21962
rect 28916 -22042 28956 -21962
rect 29036 -22042 29076 -21962
rect 29156 -22042 29196 -21962
rect 29276 -22042 29336 -21962
rect 29416 -22042 29476 -21962
rect 29556 -22042 29956 -21962
rect 23816 -22102 29956 -22042
rect 23816 -22182 24236 -22102
rect 24316 -22182 24376 -22102
rect 24456 -22182 24516 -22102
rect 24596 -22182 24636 -22102
rect 24716 -22182 24756 -22102
rect 24836 -22182 24876 -22102
rect 24956 -22182 24996 -22102
rect 25076 -22182 25116 -22102
rect 25196 -22182 25236 -22102
rect 25316 -22182 25356 -22102
rect 25436 -22182 25476 -22102
rect 25556 -22182 25596 -22102
rect 25676 -22182 25716 -22102
rect 25796 -22182 25836 -22102
rect 25916 -22182 25956 -22102
rect 26036 -22182 26076 -22102
rect 26156 -22182 26196 -22102
rect 26276 -22182 26316 -22102
rect 26396 -22182 26436 -22102
rect 26516 -22182 26556 -22102
rect 26636 -22182 26676 -22102
rect 26756 -22182 26796 -22102
rect 26876 -22182 26916 -22102
rect 26996 -22182 27036 -22102
rect 27116 -22182 27156 -22102
rect 27236 -22182 27276 -22102
rect 27356 -22182 27396 -22102
rect 27476 -22182 27516 -22102
rect 27596 -22182 27636 -22102
rect 27716 -22182 27756 -22102
rect 27836 -22182 27876 -22102
rect 27956 -22182 27996 -22102
rect 28076 -22182 28116 -22102
rect 28196 -22182 28236 -22102
rect 28316 -22182 28356 -22102
rect 28436 -22182 28476 -22102
rect 28556 -22182 28596 -22102
rect 28676 -22182 28716 -22102
rect 28796 -22182 28836 -22102
rect 28916 -22182 28956 -22102
rect 29036 -22182 29076 -22102
rect 29156 -22182 29196 -22102
rect 29276 -22182 29336 -22102
rect 29416 -22182 29476 -22102
rect 29556 -22182 29956 -22102
rect 30136 -21962 30336 -21902
rect 30396 -21962 30936 -21902
rect 30996 -21962 31576 -21902
rect 31636 -21962 31696 -21902
rect 31756 -21962 31816 -21902
rect 31896 -21962 31956 -21902
rect 32016 -21962 32176 -21902
rect 32236 -21962 32796 -21902
rect 32856 -21962 32916 -21902
rect 30136 -22082 32916 -21962
rect 30136 -22142 30336 -22082
rect 30396 -22142 30936 -22082
rect 30996 -22142 31576 -22082
rect 31636 -22142 31696 -22082
rect 31756 -22142 31816 -22082
rect 31896 -22142 31956 -22082
rect 32016 -22142 32176 -22082
rect 32236 -22142 32796 -22082
rect 32856 -22142 32916 -22082
rect 30136 -22162 32916 -22142
rect 23816 -22242 29956 -22182
rect 23816 -22322 24236 -22242
rect 24316 -22322 24376 -22242
rect 24456 -22322 24516 -22242
rect 24596 -22322 24636 -22242
rect 24716 -22322 24756 -22242
rect 24836 -22322 24876 -22242
rect 24956 -22322 24996 -22242
rect 25076 -22322 25116 -22242
rect 25196 -22322 25236 -22242
rect 25316 -22322 25356 -22242
rect 25436 -22322 25476 -22242
rect 25556 -22322 25596 -22242
rect 25676 -22322 25716 -22242
rect 25796 -22322 25836 -22242
rect 25916 -22322 25956 -22242
rect 26036 -22322 26076 -22242
rect 26156 -22322 26196 -22242
rect 26276 -22322 26316 -22242
rect 26396 -22322 26436 -22242
rect 26516 -22322 26556 -22242
rect 26636 -22322 26676 -22242
rect 26756 -22322 26796 -22242
rect 26876 -22322 26916 -22242
rect 26996 -22322 27036 -22242
rect 27116 -22322 27156 -22242
rect 27236 -22322 27276 -22242
rect 27356 -22322 27396 -22242
rect 27476 -22322 27516 -22242
rect 27596 -22322 27636 -22242
rect 27716 -22322 27756 -22242
rect 27836 -22322 27876 -22242
rect 27956 -22322 27996 -22242
rect 28076 -22322 28116 -22242
rect 28196 -22322 28236 -22242
rect 28316 -22322 28356 -22242
rect 28436 -22322 28476 -22242
rect 28556 -22322 28596 -22242
rect 28676 -22322 28716 -22242
rect 28796 -22322 28836 -22242
rect 28916 -22322 28956 -22242
rect 29036 -22322 29076 -22242
rect 29156 -22322 29196 -22242
rect 29276 -22322 29336 -22242
rect 29416 -22322 29476 -22242
rect 29556 -22322 29956 -22242
rect 23816 -22342 29956 -22322
rect 20956 -22442 32816 -22422
rect 20956 -22522 20976 -22442
rect 21056 -22522 21076 -22442
rect 21156 -22522 21176 -22442
rect 21256 -22522 21276 -22442
rect 21356 -22522 21376 -22442
rect 21456 -22522 21476 -22442
rect 21556 -22522 21576 -22442
rect 21656 -22522 21676 -22442
rect 21756 -22522 21776 -22442
rect 21856 -22522 21876 -22442
rect 21956 -22522 21976 -22442
rect 22056 -22522 22076 -22442
rect 22156 -22522 22176 -22442
rect 22256 -22522 22276 -22442
rect 22356 -22522 22376 -22442
rect 22456 -22522 22476 -22442
rect 22556 -22522 22576 -22442
rect 22656 -22522 22676 -22442
rect 22756 -22522 22776 -22442
rect 22856 -22522 22876 -22442
rect 22956 -22522 22976 -22442
rect 23056 -22522 23076 -22442
rect 23156 -22522 23176 -22442
rect 23256 -22522 23276 -22442
rect 23356 -22502 23516 -22442
rect 23576 -22502 23616 -22442
rect 23676 -22502 23756 -22442
rect 23836 -22502 23916 -22442
rect 23976 -22502 24016 -22442
rect 24076 -22502 25216 -22442
rect 23356 -22522 25216 -22502
rect 25296 -22522 25356 -22442
rect 25436 -22522 25496 -22442
rect 25576 -22522 26716 -22442
rect 26796 -22522 26856 -22442
rect 26936 -22522 26996 -22442
rect 27076 -22522 28216 -22442
rect 28296 -22522 28356 -22442
rect 28436 -22522 28496 -22442
rect 28576 -22502 29716 -22442
rect 29776 -22502 29816 -22442
rect 29876 -22502 29956 -22442
rect 30036 -22502 30116 -22442
rect 30176 -22502 30216 -22442
rect 30276 -22502 30416 -22442
rect 28576 -22522 30416 -22502
rect 30496 -22522 30516 -22442
rect 30596 -22522 30616 -22442
rect 30696 -22522 30716 -22442
rect 30796 -22522 30816 -22442
rect 30896 -22522 30916 -22442
rect 30996 -22522 31016 -22442
rect 31096 -22522 31116 -22442
rect 31196 -22522 31216 -22442
rect 31296 -22522 31316 -22442
rect 31396 -22522 31416 -22442
rect 31496 -22522 31516 -22442
rect 31596 -22522 31616 -22442
rect 31696 -22522 31716 -22442
rect 31796 -22522 31816 -22442
rect 31896 -22522 31916 -22442
rect 31996 -22522 32016 -22442
rect 32096 -22522 32116 -22442
rect 32196 -22522 32216 -22442
rect 32296 -22522 32316 -22442
rect 32396 -22522 32416 -22442
rect 32496 -22522 32516 -22442
rect 32596 -22522 32616 -22442
rect 32696 -22522 32716 -22442
rect 32796 -22522 32816 -22442
rect 20956 -22582 32816 -22522
rect 20956 -22662 20976 -22582
rect 21056 -22662 21076 -22582
rect 21156 -22662 21176 -22582
rect 21256 -22662 21276 -22582
rect 21356 -22662 21376 -22582
rect 21456 -22662 21476 -22582
rect 21556 -22662 21576 -22582
rect 21656 -22662 21676 -22582
rect 21756 -22662 21776 -22582
rect 21856 -22662 21876 -22582
rect 21956 -22662 21976 -22582
rect 22056 -22662 22076 -22582
rect 22156 -22662 22176 -22582
rect 22256 -22662 22276 -22582
rect 22356 -22662 22376 -22582
rect 22456 -22662 22476 -22582
rect 22556 -22662 22576 -22582
rect 22656 -22662 22676 -22582
rect 22756 -22662 22776 -22582
rect 22856 -22662 22876 -22582
rect 22956 -22662 22976 -22582
rect 23056 -22662 23076 -22582
rect 23156 -22662 23176 -22582
rect 23256 -22662 23276 -22582
rect 23356 -22662 23516 -22582
rect 23596 -22662 23636 -22582
rect 23696 -22662 23756 -22582
rect 23836 -22662 23896 -22582
rect 23956 -22662 23996 -22582
rect 24076 -22662 25216 -22582
rect 25296 -22662 25356 -22582
rect 25436 -22662 25496 -22582
rect 25576 -22662 26716 -22582
rect 26796 -22662 26856 -22582
rect 26936 -22662 26996 -22582
rect 27076 -22662 28216 -22582
rect 28296 -22662 28356 -22582
rect 28436 -22662 28496 -22582
rect 28576 -22662 29716 -22582
rect 29796 -22662 29836 -22582
rect 29896 -22662 29956 -22582
rect 30036 -22662 30096 -22582
rect 30156 -22662 30196 -22582
rect 30276 -22662 30416 -22582
rect 30496 -22662 30516 -22582
rect 30596 -22662 30616 -22582
rect 30696 -22662 30716 -22582
rect 30796 -22662 30816 -22582
rect 30896 -22662 30916 -22582
rect 30996 -22662 31016 -22582
rect 31096 -22662 31116 -22582
rect 31196 -22662 31216 -22582
rect 31296 -22662 31316 -22582
rect 31396 -22662 31416 -22582
rect 31496 -22662 31516 -22582
rect 31596 -22662 31616 -22582
rect 31696 -22662 31716 -22582
rect 31796 -22662 31816 -22582
rect 31896 -22662 31916 -22582
rect 31996 -22662 32016 -22582
rect 32096 -22662 32116 -22582
rect 32196 -22662 32216 -22582
rect 32296 -22662 32316 -22582
rect 32396 -22662 32416 -22582
rect 32496 -22662 32516 -22582
rect 32596 -22662 32616 -22582
rect 32696 -22662 32716 -22582
rect 32796 -22662 32816 -22582
rect 20956 -22722 32816 -22662
rect 20956 -22802 20976 -22722
rect 21056 -22802 21076 -22722
rect 21156 -22802 21176 -22722
rect 21256 -22802 21276 -22722
rect 21356 -22802 21376 -22722
rect 21456 -22802 21476 -22722
rect 21556 -22802 21576 -22722
rect 21656 -22802 21676 -22722
rect 21756 -22802 21776 -22722
rect 21856 -22802 21876 -22722
rect 21956 -22802 21976 -22722
rect 22056 -22802 22076 -22722
rect 22156 -22802 22176 -22722
rect 22256 -22802 22276 -22722
rect 22356 -22802 22376 -22722
rect 22456 -22802 22476 -22722
rect 22556 -22802 22576 -22722
rect 22656 -22802 22676 -22722
rect 22756 -22802 22776 -22722
rect 22856 -22802 22876 -22722
rect 22956 -22802 22976 -22722
rect 23056 -22802 23076 -22722
rect 23156 -22802 23176 -22722
rect 23256 -22802 23276 -22722
rect 23356 -22742 25216 -22722
rect 23356 -22802 23516 -22742
rect 23576 -22802 23616 -22742
rect 23676 -22802 23756 -22742
rect 23836 -22802 23916 -22742
rect 23976 -22802 24016 -22742
rect 24076 -22802 25216 -22742
rect 25296 -22802 25356 -22722
rect 25436 -22802 25496 -22722
rect 25576 -22802 26716 -22722
rect 26796 -22802 26856 -22722
rect 26936 -22802 26996 -22722
rect 27076 -22802 28216 -22722
rect 28296 -22802 28356 -22722
rect 28436 -22802 28496 -22722
rect 28576 -22742 30416 -22722
rect 28576 -22802 29716 -22742
rect 29776 -22802 29816 -22742
rect 29876 -22802 29956 -22742
rect 30036 -22802 30116 -22742
rect 30176 -22802 30216 -22742
rect 30276 -22802 30416 -22742
rect 30496 -22802 30516 -22722
rect 30596 -22802 30616 -22722
rect 30696 -22802 30716 -22722
rect 30796 -22802 30816 -22722
rect 30896 -22802 30916 -22722
rect 30996 -22802 31016 -22722
rect 31096 -22802 31116 -22722
rect 31196 -22802 31216 -22722
rect 31296 -22802 31316 -22722
rect 31396 -22802 31416 -22722
rect 31496 -22802 31516 -22722
rect 31596 -22802 31616 -22722
rect 31696 -22802 31716 -22722
rect 31796 -22802 31816 -22722
rect 31896 -22802 31916 -22722
rect 31996 -22802 32016 -22722
rect 32096 -22802 32116 -22722
rect 32196 -22802 32216 -22722
rect 32296 -22802 32316 -22722
rect 32396 -22802 32416 -22722
rect 32496 -22802 32516 -22722
rect 32596 -22802 32616 -22722
rect 32696 -22802 32716 -22722
rect 32796 -22802 32816 -22722
rect 20956 -22822 32816 -22802
rect 26696 -22922 27096 -22902
rect 20676 -22982 22416 -22962
rect 20676 -23042 21856 -22982
rect 21916 -23042 22316 -22982
rect 22376 -23042 22416 -22982
rect 20676 -23062 20836 -23042
rect 20676 -23122 20716 -23062
rect 20796 -23102 20836 -23062
rect 20896 -23062 21096 -23042
rect 20896 -23102 20956 -23062
rect 20796 -23122 20956 -23102
rect 21036 -23102 21096 -23062
rect 21156 -23062 22416 -23042
rect 21156 -23102 21196 -23062
rect 21036 -23122 21196 -23102
rect 21276 -23122 22416 -23062
rect 20676 -23162 22416 -23122
rect 20676 -23222 20716 -23162
rect 20796 -23222 20836 -23162
rect 20896 -23222 20956 -23162
rect 21036 -23222 21096 -23162
rect 21156 -23222 21196 -23162
rect 21276 -23222 21856 -23162
rect 21916 -23222 22316 -23162
rect 22376 -23222 22416 -23162
rect 20676 -23242 22416 -23222
rect 26696 -23002 26716 -22922
rect 26796 -23002 26856 -22922
rect 26936 -23002 26996 -22922
rect 27076 -23002 27096 -22922
rect 26696 -23042 27096 -23002
rect 26696 -23122 26716 -23042
rect 26796 -23122 26856 -23042
rect 26936 -23122 26996 -23042
rect 27076 -23122 27096 -23042
rect 26696 -23162 27096 -23122
rect 26696 -23242 26716 -23162
rect 26796 -23242 26856 -23162
rect 26936 -23242 26996 -23162
rect 27076 -23242 27096 -23162
rect 31436 -22982 33176 -22962
rect 31436 -23042 31456 -22982
rect 31516 -23042 31916 -22982
rect 31976 -23042 33176 -22982
rect 31436 -23062 32636 -23042
rect 31436 -23122 32516 -23062
rect 32596 -23102 32636 -23062
rect 32696 -23062 32896 -23042
rect 32696 -23102 32756 -23062
rect 32596 -23122 32756 -23102
rect 32836 -23102 32896 -23062
rect 32956 -23062 33176 -23042
rect 32956 -23102 32996 -23062
rect 32836 -23122 32996 -23102
rect 33076 -23122 33176 -23062
rect 31436 -23162 33176 -23122
rect 31436 -23222 31456 -23162
rect 31516 -23222 31916 -23162
rect 31976 -23222 32516 -23162
rect 32596 -23222 32636 -23162
rect 32696 -23222 32756 -23162
rect 32836 -23222 32896 -23162
rect 32956 -23222 32996 -23162
rect 33076 -23222 33176 -23162
rect 31436 -23242 33176 -23222
rect 26696 -23282 27096 -23242
rect 26696 -23362 26716 -23282
rect 26796 -23362 26856 -23282
rect 26936 -23362 26996 -23282
rect 27076 -23362 27096 -23282
rect 26696 -23402 27096 -23362
rect 23796 -23442 24596 -23422
rect 21736 -23462 22236 -23442
rect 21736 -23522 21916 -23462
rect 21976 -23522 22016 -23462
rect 22076 -23522 22116 -23462
rect 22176 -23522 22236 -23462
rect 21736 -23562 22236 -23522
rect 21736 -23622 21916 -23562
rect 21976 -23622 22016 -23562
rect 22076 -23622 22116 -23562
rect 22176 -23622 22236 -23562
rect 21736 -23642 22236 -23622
rect 23776 -23462 24236 -23442
rect 23776 -23522 23796 -23462
rect 23856 -23522 24116 -23462
rect 24176 -23522 24236 -23462
rect 24316 -23522 24356 -23442
rect 24456 -23522 24496 -23442
rect 24576 -23522 24596 -23442
rect 23776 -23542 24596 -23522
rect 23776 -23602 23796 -23542
rect 23856 -23602 24116 -23542
rect 24176 -23602 24596 -23542
rect 23776 -23622 24596 -23602
rect 23776 -23682 23796 -23622
rect 23856 -23682 24116 -23622
rect 24176 -23682 24236 -23622
rect 23776 -23702 24236 -23682
rect 24316 -23702 24356 -23622
rect 24456 -23702 24496 -23622
rect 24576 -23702 24596 -23622
rect 23796 -23722 24596 -23702
rect 25196 -23442 25976 -23422
rect 25196 -23522 25216 -23442
rect 25296 -23522 25336 -23442
rect 25456 -23522 25496 -23442
rect 25576 -23462 25996 -23442
rect 25576 -23522 25596 -23462
rect 25656 -23522 25916 -23462
rect 25976 -23522 25996 -23462
rect 25196 -23542 25996 -23522
rect 25196 -23602 25596 -23542
rect 25656 -23602 25916 -23542
rect 25976 -23602 25996 -23542
rect 25196 -23622 25996 -23602
rect 25196 -23702 25216 -23622
rect 25296 -23702 25336 -23622
rect 25456 -23702 25496 -23622
rect 25576 -23682 25596 -23622
rect 25656 -23682 25916 -23622
rect 25976 -23682 25996 -23622
rect 25576 -23702 25996 -23682
rect 26696 -23482 26716 -23402
rect 26796 -23482 26856 -23402
rect 26936 -23482 26996 -23402
rect 27076 -23482 27096 -23402
rect 27796 -23442 28596 -23422
rect 26696 -23522 27096 -23482
rect 26696 -23602 26716 -23522
rect 26796 -23602 26856 -23522
rect 26936 -23602 26996 -23522
rect 27076 -23602 27096 -23522
rect 26696 -23642 27096 -23602
rect 25196 -23722 25976 -23702
rect 26696 -23722 26716 -23642
rect 26796 -23722 26856 -23642
rect 26936 -23722 26996 -23642
rect 27076 -23722 27096 -23642
rect 27776 -23462 28216 -23442
rect 27776 -23522 27796 -23462
rect 27856 -23522 28116 -23462
rect 28176 -23522 28216 -23462
rect 28296 -23522 28336 -23442
rect 28456 -23522 28496 -23442
rect 28576 -23522 28596 -23442
rect 27776 -23542 28596 -23522
rect 27776 -23602 27796 -23542
rect 27856 -23602 28116 -23542
rect 28176 -23602 28596 -23542
rect 27776 -23622 28596 -23602
rect 27776 -23682 27796 -23622
rect 27856 -23682 28116 -23622
rect 28176 -23682 28216 -23622
rect 27776 -23702 28216 -23682
rect 28296 -23702 28336 -23622
rect 28456 -23702 28496 -23622
rect 28576 -23702 28596 -23622
rect 27796 -23722 28596 -23702
rect 29196 -23442 29976 -23422
rect 29196 -23522 29216 -23442
rect 29296 -23522 29336 -23442
rect 29436 -23522 29476 -23442
rect 29556 -23462 29996 -23442
rect 29556 -23522 29596 -23462
rect 29656 -23522 29916 -23462
rect 29976 -23522 29996 -23462
rect 29196 -23542 29996 -23522
rect 29196 -23602 29596 -23542
rect 29656 -23602 29916 -23542
rect 29976 -23602 29996 -23542
rect 29196 -23622 29996 -23602
rect 29196 -23702 29216 -23622
rect 29296 -23702 29336 -23622
rect 29436 -23702 29476 -23622
rect 29556 -23682 29596 -23622
rect 29656 -23682 29916 -23622
rect 29976 -23682 29996 -23622
rect 31556 -23462 32056 -23442
rect 31556 -23522 31636 -23462
rect 31696 -23522 31756 -23462
rect 31816 -23522 31856 -23462
rect 31916 -23522 32056 -23462
rect 31556 -23562 32056 -23522
rect 31556 -23622 31636 -23562
rect 31696 -23622 31756 -23562
rect 31816 -23622 31856 -23562
rect 31916 -23622 32056 -23562
rect 31556 -23642 32056 -23622
rect 29556 -23702 29996 -23682
rect 29196 -23722 29976 -23702
rect 26696 -23762 27096 -23722
rect 26696 -23842 26716 -23762
rect 26796 -23842 26856 -23762
rect 26936 -23842 26996 -23762
rect 27076 -23842 27096 -23762
rect 26696 -23882 27096 -23842
rect 26416 -23942 26596 -23922
rect 26416 -24082 26436 -23942
rect 26576 -24082 26596 -23942
rect 22796 -24122 23156 -24102
rect 22796 -24202 22816 -24122
rect 22896 -24202 22936 -24122
rect 23016 -24202 23056 -24122
rect 23136 -24202 23156 -24122
rect 22796 -24242 23156 -24202
rect 22796 -24302 22816 -24242
rect 22876 -24302 22936 -24242
rect 23016 -24302 23076 -24242
rect 23136 -24262 23156 -24242
rect 23856 -24142 24116 -24122
rect 23856 -24202 23876 -24142
rect 23936 -24202 24036 -24142
rect 24096 -24202 24116 -24142
rect 23856 -24262 24116 -24202
rect 24936 -24142 25916 -24122
rect 24996 -24202 25036 -24142
rect 25096 -24202 25676 -24142
rect 25736 -24202 25836 -24142
rect 25896 -24202 25916 -24142
rect 24936 -24222 25916 -24202
rect 26416 -24262 26596 -24082
rect 23136 -24282 26596 -24262
rect 23136 -24302 24696 -24282
rect 22796 -24342 24696 -24302
rect 24756 -24342 26596 -24282
rect 22796 -24422 22816 -24342
rect 22896 -24422 22936 -24342
rect 23016 -24422 23056 -24342
rect 23136 -24362 26596 -24342
rect 23136 -24422 24776 -24362
rect 24836 -24422 26596 -24362
rect 22796 -24442 26596 -24422
rect 26696 -23962 26716 -23882
rect 26796 -23962 26856 -23882
rect 26936 -23962 26996 -23882
rect 27076 -23962 27096 -23882
rect 26696 -24002 27096 -23962
rect 26696 -24082 26716 -24002
rect 26796 -24082 26856 -24002
rect 26936 -24082 26996 -24002
rect 27076 -24082 27096 -24002
rect 26696 -24122 27096 -24082
rect 26696 -24202 26716 -24122
rect 26796 -24202 26856 -24122
rect 26936 -24202 26996 -24122
rect 27076 -24202 27096 -24122
rect 26696 -24242 27096 -24202
rect 26696 -24322 26716 -24242
rect 26796 -24322 26856 -24242
rect 26936 -24322 26996 -24242
rect 27076 -24322 27096 -24242
rect 26696 -24362 27096 -24322
rect 26696 -24442 26716 -24362
rect 26796 -24442 26856 -24362
rect 26936 -24442 26996 -24362
rect 27076 -24442 27096 -24362
rect 27196 -23942 27376 -23922
rect 27196 -24082 27216 -23942
rect 27356 -24082 27376 -23942
rect 27196 -24262 27376 -24082
rect 27856 -24142 28856 -24122
rect 27856 -24202 27876 -24142
rect 27936 -24202 28036 -24142
rect 28096 -24202 28696 -24142
rect 28756 -24202 28796 -24142
rect 27856 -24222 28856 -24202
rect 29656 -24142 29916 -24122
rect 29656 -24202 29676 -24142
rect 29736 -24202 29836 -24142
rect 29896 -24202 29916 -24142
rect 29656 -24262 29916 -24202
rect 30636 -24262 30996 -24102
rect 27196 -24282 30996 -24262
rect 27196 -24342 29036 -24282
rect 29096 -24342 30996 -24282
rect 27196 -24362 30996 -24342
rect 27196 -24422 28956 -24362
rect 29016 -24422 30996 -24362
rect 27196 -24442 30996 -24422
rect 26696 -24482 27096 -24442
rect 22796 -24522 26596 -24502
rect 22796 -24582 25036 -24522
rect 25096 -24582 26596 -24522
rect 22796 -24602 26596 -24582
rect 22796 -24662 24956 -24602
rect 25016 -24662 26596 -24602
rect 22796 -24682 26596 -24662
rect 22796 -24842 23156 -24682
rect 23856 -24742 24116 -24682
rect 23856 -24802 23876 -24742
rect 23936 -24802 24036 -24742
rect 24096 -24802 24116 -24742
rect 23856 -24822 24116 -24802
rect 24676 -24742 25916 -24722
rect 24676 -24802 24696 -24742
rect 24756 -24802 24796 -24742
rect 24856 -24802 25676 -24742
rect 25736 -24802 25836 -24742
rect 25896 -24802 25916 -24742
rect 24676 -24822 25916 -24802
rect 26416 -24862 26596 -24682
rect 23796 -24942 25596 -24922
rect 23776 -24962 25216 -24942
rect 21216 -24982 22916 -24962
rect 21216 -25042 21416 -24982
rect 21476 -25042 21776 -24982
rect 21836 -25042 21896 -24982
rect 21956 -25042 22036 -24982
rect 22096 -25042 22636 -24982
rect 22696 -25042 22916 -24982
rect 21216 -25162 22916 -25042
rect 21216 -25222 21416 -25162
rect 21476 -25222 21776 -25162
rect 21836 -25222 21896 -25162
rect 21956 -25222 22036 -25162
rect 22096 -25222 22636 -25162
rect 22696 -25222 22916 -25162
rect 23776 -25022 23796 -24962
rect 23856 -25022 24116 -24962
rect 24176 -25022 25216 -24962
rect 25296 -25022 25336 -24942
rect 25456 -25022 25496 -24942
rect 25576 -25022 25596 -24942
rect 26416 -25002 26436 -24862
rect 26576 -25002 26596 -24862
rect 26416 -25022 26596 -25002
rect 26696 -24562 26716 -24482
rect 26796 -24562 26856 -24482
rect 26936 -24562 26996 -24482
rect 27076 -24562 27096 -24482
rect 26696 -24602 27096 -24562
rect 26696 -24682 26716 -24602
rect 26796 -24682 26856 -24602
rect 26936 -24682 26996 -24602
rect 27076 -24682 27096 -24602
rect 26696 -24722 27096 -24682
rect 26696 -24802 26716 -24722
rect 26796 -24802 26856 -24722
rect 26936 -24802 26996 -24722
rect 27076 -24802 27096 -24722
rect 26696 -24842 27096 -24802
rect 26696 -24922 26716 -24842
rect 26796 -24922 26856 -24842
rect 26936 -24922 26996 -24842
rect 27076 -24922 27096 -24842
rect 26696 -24962 27096 -24922
rect 23776 -25042 25596 -25022
rect 23776 -25102 23796 -25042
rect 23856 -25102 24116 -25042
rect 24176 -25102 25596 -25042
rect 23776 -25122 25596 -25102
rect 23776 -25182 23796 -25122
rect 23856 -25182 24116 -25122
rect 24176 -25182 25216 -25122
rect 23776 -25202 25216 -25182
rect 25296 -25202 25336 -25122
rect 25456 -25202 25496 -25122
rect 25576 -25202 25596 -25122
rect 23796 -25222 25596 -25202
rect 26696 -25042 26716 -24962
rect 26796 -25042 26856 -24962
rect 26936 -25042 26996 -24962
rect 27076 -25042 27096 -24962
rect 27196 -24522 30996 -24502
rect 27196 -24582 28696 -24522
rect 28756 -24582 30656 -24522
rect 27196 -24602 30656 -24582
rect 30736 -24602 30776 -24522
rect 30856 -24602 30896 -24522
rect 30976 -24602 30996 -24522
rect 27196 -24662 28776 -24602
rect 28836 -24642 30996 -24602
rect 28836 -24662 30656 -24642
rect 27196 -24682 30656 -24662
rect 27196 -24862 27376 -24682
rect 27856 -24742 29116 -24722
rect 27856 -24802 27876 -24742
rect 27936 -24802 28036 -24742
rect 28096 -24802 28936 -24742
rect 28996 -24802 29036 -24742
rect 29096 -24802 29116 -24742
rect 27856 -24822 29116 -24802
rect 29656 -24742 29916 -24682
rect 29656 -24802 29676 -24742
rect 29736 -24802 29836 -24742
rect 29896 -24802 29916 -24742
rect 29656 -24822 29916 -24802
rect 30636 -24702 30656 -24682
rect 30736 -24702 30776 -24642
rect 30856 -24702 30896 -24642
rect 30976 -24702 30996 -24642
rect 30636 -24742 30996 -24702
rect 30636 -24822 30656 -24742
rect 30736 -24822 30776 -24742
rect 30856 -24822 30896 -24742
rect 30976 -24822 30996 -24742
rect 30636 -24842 30996 -24822
rect 27196 -25002 27216 -24862
rect 27356 -25002 27376 -24862
rect 27196 -25022 27376 -25002
rect 28196 -24942 29976 -24922
rect 28196 -25022 28216 -24942
rect 28296 -25022 28336 -24942
rect 28456 -25022 28496 -24942
rect 28576 -24962 29996 -24942
rect 28576 -25022 29596 -24962
rect 29656 -25022 29916 -24962
rect 29976 -25022 29996 -24962
rect 26696 -25082 27096 -25042
rect 26696 -25162 26716 -25082
rect 26796 -25162 26856 -25082
rect 26936 -25162 26996 -25082
rect 27076 -25162 27096 -25082
rect 26696 -25202 27096 -25162
rect 21216 -25242 22916 -25222
rect 26696 -25282 26716 -25202
rect 26796 -25282 26856 -25202
rect 26936 -25282 26996 -25202
rect 27076 -25282 27096 -25202
rect 28196 -25042 29996 -25022
rect 28196 -25102 29596 -25042
rect 29656 -25102 29916 -25042
rect 29976 -25102 29996 -25042
rect 28196 -25122 29996 -25102
rect 28196 -25202 28216 -25122
rect 28296 -25202 28336 -25122
rect 28456 -25202 28496 -25122
rect 28576 -25182 29596 -25122
rect 29656 -25182 29916 -25122
rect 29976 -25182 29996 -25122
rect 28576 -25202 29996 -25182
rect 30876 -24982 32576 -24962
rect 30876 -25042 31076 -24982
rect 31136 -25042 31696 -24982
rect 31756 -25042 31836 -24982
rect 31896 -25042 31956 -24982
rect 32016 -25042 32296 -24982
rect 32356 -25042 32576 -24982
rect 30876 -25162 32576 -25042
rect 28196 -25222 29976 -25202
rect 30876 -25222 31076 -25162
rect 31136 -25222 31696 -25162
rect 31756 -25222 31836 -25162
rect 31896 -25222 31956 -25162
rect 32016 -25222 32296 -25162
rect 32356 -25222 32576 -25162
rect 30876 -25242 32576 -25222
rect 26696 -25322 27096 -25282
rect 26696 -25402 26716 -25322
rect 26796 -25402 26856 -25322
rect 26936 -25402 26996 -25322
rect 27076 -25402 27096 -25322
rect 26696 -25442 27096 -25402
rect 26696 -25522 26716 -25442
rect 26796 -25522 26856 -25442
rect 26936 -25522 26996 -25442
rect 27076 -25522 27096 -25442
rect 24196 -25542 25976 -25522
rect 24196 -25622 24236 -25542
rect 24316 -25622 24356 -25542
rect 24476 -25622 24516 -25542
rect 24596 -25562 25996 -25542
rect 24596 -25622 25596 -25562
rect 25656 -25622 25916 -25562
rect 25976 -25622 25996 -25562
rect 24196 -25642 25996 -25622
rect 24196 -25702 25596 -25642
rect 25656 -25702 25916 -25642
rect 25976 -25702 25996 -25642
rect 24196 -25722 25996 -25702
rect 24196 -25802 24236 -25722
rect 24316 -25802 24356 -25722
rect 24476 -25802 24516 -25722
rect 24596 -25782 25596 -25722
rect 25656 -25782 25916 -25722
rect 25976 -25782 25996 -25722
rect 24596 -25802 25996 -25782
rect 26696 -25562 27096 -25522
rect 27796 -25542 29596 -25522
rect 26696 -25642 26716 -25562
rect 26796 -25642 26856 -25562
rect 26936 -25642 26996 -25562
rect 27076 -25642 27096 -25562
rect 26696 -25682 27096 -25642
rect 26696 -25762 26716 -25682
rect 26796 -25762 26856 -25682
rect 26936 -25762 26996 -25682
rect 27076 -25762 27096 -25682
rect 26696 -25802 27096 -25762
rect 27776 -25562 29196 -25542
rect 27776 -25622 27796 -25562
rect 27856 -25622 28116 -25562
rect 28176 -25622 29196 -25562
rect 29276 -25622 29316 -25542
rect 29436 -25622 29476 -25542
rect 29556 -25622 29596 -25542
rect 27776 -25642 29596 -25622
rect 27776 -25702 27796 -25642
rect 27856 -25702 28116 -25642
rect 28176 -25702 29596 -25642
rect 27776 -25722 29596 -25702
rect 27776 -25782 27796 -25722
rect 27856 -25782 28116 -25722
rect 28176 -25782 29196 -25722
rect 27776 -25802 29196 -25782
rect 29276 -25802 29316 -25722
rect 29436 -25802 29476 -25722
rect 29556 -25802 29596 -25722
rect 24196 -25822 25976 -25802
rect 26696 -25882 26716 -25802
rect 26796 -25882 26856 -25802
rect 26936 -25882 26996 -25802
rect 27076 -25882 27096 -25802
rect 27796 -25822 29596 -25802
rect 26696 -25922 27096 -25882
rect 26696 -26002 26716 -25922
rect 26796 -26002 26856 -25922
rect 26936 -26002 26996 -25922
rect 27076 -26002 27096 -25922
rect 26696 -26482 27096 -26002
rect 21396 -26502 24696 -26482
rect 21396 -26562 21496 -26502
rect 21556 -26562 21576 -26502
rect 21636 -26562 21656 -26502
rect 21716 -26562 21736 -26502
rect 21796 -26562 21816 -26502
rect 21876 -26562 21896 -26502
rect 21956 -26562 21976 -26502
rect 22036 -26562 22056 -26502
rect 22116 -26562 22136 -26502
rect 22196 -26562 22216 -26502
rect 22276 -26562 22296 -26502
rect 22356 -26562 22376 -26502
rect 22436 -26562 22456 -26502
rect 22556 -26562 22576 -26502
rect 22636 -26562 24376 -26502
rect 24436 -26562 24476 -26502
rect 24536 -26562 24696 -26502
rect 21396 -26582 24696 -26562
rect 21396 -26602 24376 -26582
rect 21396 -26662 21496 -26602
rect 21556 -26662 21576 -26602
rect 21636 -26662 21656 -26602
rect 21716 -26662 21736 -26602
rect 21796 -26662 21816 -26602
rect 21876 -26662 21896 -26602
rect 21956 -26662 21976 -26602
rect 22036 -26662 22056 -26602
rect 22116 -26662 22136 -26602
rect 22196 -26662 22216 -26602
rect 22276 -26662 22296 -26602
rect 22356 -26662 22376 -26602
rect 22436 -26662 22456 -26602
rect 22556 -26662 22576 -26602
rect 22636 -26642 24376 -26602
rect 24436 -26642 24476 -26582
rect 24536 -26642 24696 -26582
rect 22636 -26662 24696 -26642
rect 21396 -26762 24696 -26662
rect 21396 -26822 24376 -26762
rect 24436 -26822 24476 -26762
rect 24536 -26822 24696 -26762
rect 21396 -26842 24696 -26822
rect 21396 -26902 24376 -26842
rect 24436 -26902 24476 -26842
rect 24536 -26902 24696 -26842
rect 21396 -26922 24696 -26902
rect 24790 -26522 28930 -26482
rect 24790 -26582 24956 -26522
rect 25016 -26582 25036 -26522
rect 25096 -26582 26176 -26522
rect 26236 -26582 26256 -26522
rect 26316 -26582 27416 -26522
rect 27476 -26582 27496 -26522
rect 27556 -26582 28636 -26522
rect 28696 -26582 28716 -26522
rect 28776 -26582 28930 -26522
rect 24790 -26602 28930 -26582
rect 24790 -26662 24956 -26602
rect 25016 -26662 25036 -26602
rect 25096 -26662 26176 -26602
rect 26236 -26662 26256 -26602
rect 26316 -26662 27416 -26602
rect 27476 -26662 27496 -26602
rect 27556 -26662 28636 -26602
rect 28696 -26662 28716 -26602
rect 28776 -26662 28930 -26602
rect 24790 -26682 28930 -26662
rect 24790 -26742 24956 -26682
rect 25016 -26742 25036 -26682
rect 25096 -26742 26176 -26682
rect 26236 -26742 26256 -26682
rect 26316 -26742 27416 -26682
rect 27476 -26742 27496 -26682
rect 27556 -26742 28636 -26682
rect 28696 -26742 28716 -26682
rect 28776 -26742 28930 -26682
rect 24790 -26762 28930 -26742
rect 24790 -26822 24956 -26762
rect 25016 -26822 25036 -26762
rect 25096 -26822 26176 -26762
rect 26236 -26822 26256 -26762
rect 26316 -26822 27416 -26762
rect 27476 -26822 27496 -26762
rect 27556 -26822 28636 -26762
rect 28696 -26822 28716 -26762
rect 28776 -26822 28930 -26762
rect 24790 -26842 28930 -26822
rect 24790 -26902 24956 -26842
rect 25016 -26902 25036 -26842
rect 25096 -26902 26176 -26842
rect 26236 -26902 26256 -26842
rect 26316 -26902 27416 -26842
rect 27476 -26902 27496 -26842
rect 27556 -26902 28636 -26842
rect 28696 -26902 28716 -26842
rect 28776 -26902 28930 -26842
rect 24790 -26922 28930 -26902
rect 29056 -26502 32356 -26482
rect 29056 -26562 29216 -26502
rect 29276 -26562 29316 -26502
rect 29376 -26562 31156 -26502
rect 31216 -26562 31236 -26502
rect 31336 -26562 31356 -26502
rect 31416 -26562 31436 -26502
rect 31496 -26562 31516 -26502
rect 31576 -26562 31596 -26502
rect 31656 -26562 31676 -26502
rect 31736 -26562 31756 -26502
rect 31816 -26562 31836 -26502
rect 31896 -26562 31916 -26502
rect 31976 -26562 31996 -26502
rect 32056 -26562 32076 -26502
rect 32136 -26562 32156 -26502
rect 32216 -26562 32236 -26502
rect 32296 -26562 32356 -26502
rect 29056 -26582 32356 -26562
rect 29056 -26642 29216 -26582
rect 29276 -26642 29316 -26582
rect 29376 -26602 32356 -26582
rect 29376 -26642 31156 -26602
rect 29056 -26662 31156 -26642
rect 31216 -26662 31236 -26602
rect 31336 -26662 31356 -26602
rect 31416 -26662 31436 -26602
rect 31496 -26662 31516 -26602
rect 31576 -26662 31596 -26602
rect 31656 -26662 31676 -26602
rect 31736 -26662 31756 -26602
rect 31816 -26662 31836 -26602
rect 31896 -26662 31916 -26602
rect 31976 -26662 31996 -26602
rect 32056 -26662 32076 -26602
rect 32136 -26662 32156 -26602
rect 32216 -26662 32236 -26602
rect 32296 -26662 32356 -26602
rect 29056 -26762 32356 -26662
rect 29056 -26822 29216 -26762
rect 29276 -26822 29316 -26762
rect 29376 -26822 32356 -26762
rect 29056 -26842 32356 -26822
rect 29056 -26902 29216 -26842
rect 29276 -26902 29316 -26842
rect 29376 -26902 32356 -26842
rect 29056 -26922 32356 -26902
rect 24356 -27102 24696 -26922
rect 29056 -27102 29396 -26922
rect 24356 -27122 29396 -27102
rect 24356 -27182 24376 -27122
rect 24436 -27182 24476 -27122
rect 24536 -27182 25556 -27122
rect 25616 -27182 25656 -27122
rect 25716 -27182 26796 -27122
rect 26856 -27182 26896 -27122
rect 26956 -27182 28016 -27122
rect 28076 -27182 28116 -27122
rect 28176 -27182 29216 -27122
rect 29276 -27182 29316 -27122
rect 29376 -27182 29396 -27122
rect 24356 -27202 29396 -27182
rect 24356 -27262 24376 -27202
rect 24436 -27262 24476 -27202
rect 24536 -27262 25556 -27202
rect 25616 -27262 25656 -27202
rect 25716 -27262 26796 -27202
rect 26856 -27262 26896 -27202
rect 26956 -27262 28016 -27202
rect 28076 -27262 28116 -27202
rect 28176 -27262 29216 -27202
rect 29276 -27262 29316 -27202
rect 29376 -27262 29396 -27202
rect 24356 -27342 29396 -27262
rect 24356 -27402 24376 -27342
rect 24436 -27402 24476 -27342
rect 24536 -27402 25556 -27342
rect 25616 -27402 25656 -27342
rect 25716 -27402 26796 -27342
rect 26856 -27402 26896 -27342
rect 26956 -27402 28016 -27342
rect 28076 -27402 28116 -27342
rect 28176 -27402 29216 -27342
rect 29276 -27402 29316 -27342
rect 29376 -27402 29396 -27342
rect 24356 -27422 29396 -27402
rect 24356 -27482 24376 -27422
rect 24436 -27482 24476 -27422
rect 24536 -27482 25556 -27422
rect 25616 -27482 25656 -27422
rect 25716 -27482 26796 -27422
rect 26856 -27482 26896 -27422
rect 26956 -27482 28016 -27422
rect 28076 -27482 28116 -27422
rect 28176 -27482 29216 -27422
rect 29276 -27482 29316 -27422
rect 29376 -27482 29396 -27422
rect 24356 -27502 29396 -27482
rect 22796 -29042 23196 -29022
rect 22796 -29122 22816 -29042
rect 22896 -29122 22956 -29042
rect 23036 -29122 23096 -29042
rect 23176 -29122 23196 -29042
rect 22796 -29182 23196 -29122
rect 22796 -29262 22816 -29182
rect 22896 -29262 22956 -29182
rect 23036 -29262 23096 -29182
rect 23176 -29262 23196 -29182
rect 22796 -29322 23196 -29262
rect 22796 -29402 22816 -29322
rect 22896 -29402 22956 -29322
rect 23036 -29402 23096 -29322
rect 23176 -29402 23196 -29322
rect 22796 -29422 23196 -29402
rect 26696 -29642 27096 -27502
rect 30596 -29042 30996 -29022
rect 30596 -29122 30616 -29042
rect 30696 -29122 30756 -29042
rect 30836 -29122 30896 -29042
rect 30976 -29122 30996 -29042
rect 30596 -29182 30996 -29122
rect 30596 -29262 30616 -29182
rect 30696 -29262 30756 -29182
rect 30836 -29262 30896 -29182
rect 30976 -29262 30996 -29182
rect 30596 -29322 30996 -29262
rect 30596 -29402 30616 -29322
rect 30696 -29402 30756 -29322
rect 30836 -29402 30896 -29322
rect 30976 -29402 30996 -29322
rect 30596 -29422 30996 -29402
rect 26696 -29702 26716 -29642
rect 26776 -29702 26816 -29642
rect 26876 -29702 26916 -29642
rect 26976 -29702 27016 -29642
rect 27076 -29702 27096 -29642
rect 26696 -29742 27096 -29702
rect 26696 -29802 26716 -29742
rect 26776 -29802 26816 -29742
rect 26876 -29802 26916 -29742
rect 26976 -29802 27016 -29742
rect 27076 -29802 27096 -29742
rect 26696 -29842 27096 -29802
rect 26696 -29902 26716 -29842
rect 26776 -29902 26816 -29842
rect 26876 -29902 26916 -29842
rect 26976 -29902 27016 -29842
rect 27076 -29902 27096 -29842
rect 26696 -29942 27096 -29902
rect 26696 -30002 26716 -29942
rect 26776 -30002 26816 -29942
rect 26876 -30002 26916 -29942
rect 26976 -30002 27016 -29942
rect 27076 -30002 27096 -29942
rect 21736 -30442 22136 -30422
rect 21736 -30502 21756 -30442
rect 21816 -30502 21856 -30442
rect 21916 -30502 21956 -30442
rect 22016 -30502 22056 -30442
rect 22116 -30502 22136 -30442
rect 21736 -30522 22136 -30502
rect 21736 -30582 21756 -30522
rect 21816 -30582 21856 -30522
rect 21916 -30582 21956 -30522
rect 22016 -30582 22056 -30522
rect 22116 -30582 22136 -30522
rect 21736 -30622 22136 -30582
rect 21736 -30682 21756 -30622
rect 21816 -30682 21856 -30622
rect 21916 -30682 21956 -30622
rect 22016 -30682 22056 -30622
rect 22116 -30682 22136 -30622
rect 21736 -30722 22136 -30682
rect 21736 -30782 21756 -30722
rect 21816 -30782 21856 -30722
rect 21916 -30782 21956 -30722
rect 22016 -30782 22056 -30722
rect 22116 -30782 22136 -30722
rect 21736 -30802 22136 -30782
rect 31656 -30442 32056 -30422
rect 31656 -30502 31676 -30442
rect 31736 -30502 31776 -30442
rect 31836 -30502 31876 -30442
rect 31936 -30502 31976 -30442
rect 32036 -30502 32056 -30442
rect 31656 -30522 32056 -30502
rect 31656 -30582 31676 -30522
rect 31736 -30582 31776 -30522
rect 31836 -30582 31876 -30522
rect 31936 -30582 31976 -30522
rect 32036 -30582 32056 -30522
rect 31656 -30622 32056 -30582
rect 31656 -30682 31676 -30622
rect 31736 -30682 31776 -30622
rect 31836 -30682 31876 -30622
rect 31936 -30682 31976 -30622
rect 32036 -30682 32056 -30622
rect 31656 -30722 32056 -30682
rect 31656 -30782 31676 -30722
rect 31736 -30782 31776 -30722
rect 31836 -30782 31876 -30722
rect 31936 -30782 31976 -30722
rect 32036 -30782 32056 -30722
rect 31656 -30802 32056 -30782
<< via2 >>
rect 26716 -21082 26796 -21002
rect 26856 -21082 26936 -21002
rect 26996 -21082 27076 -21002
rect 26716 -21202 26796 -21122
rect 26856 -21202 26936 -21122
rect 26996 -21202 27076 -21122
rect 26716 -21342 26796 -21262
rect 26856 -21342 26936 -21262
rect 26996 -21342 27076 -21262
rect 21776 -21962 21836 -21902
rect 21896 -21962 21976 -21902
rect 22036 -21962 22096 -21902
rect 21776 -22142 21836 -22082
rect 21896 -22142 21976 -22082
rect 22036 -22142 22096 -22082
rect 24236 -22042 24316 -21962
rect 24376 -22042 24456 -21962
rect 24516 -22042 24596 -21962
rect 29196 -22042 29276 -21962
rect 29336 -22042 29416 -21962
rect 29476 -22042 29556 -21962
rect 24236 -22182 24316 -22102
rect 24376 -22182 24456 -22102
rect 24516 -22182 24596 -22102
rect 29196 -22182 29276 -22102
rect 29336 -22182 29416 -22102
rect 29476 -22182 29556 -22102
rect 31696 -21962 31756 -21902
rect 31816 -21962 31896 -21902
rect 31956 -21962 32016 -21902
rect 31696 -22142 31756 -22082
rect 31816 -22142 31896 -22082
rect 31956 -22142 32016 -22082
rect 24236 -22322 24316 -22242
rect 24376 -22322 24456 -22242
rect 24516 -22322 24596 -22242
rect 29196 -22322 29276 -22242
rect 29336 -22322 29416 -22242
rect 29476 -22322 29556 -22242
rect 23516 -22502 23576 -22442
rect 23616 -22502 23676 -22442
rect 23756 -22502 23836 -22442
rect 23916 -22502 23976 -22442
rect 24016 -22502 24076 -22442
rect 25216 -22522 25296 -22442
rect 25356 -22522 25436 -22442
rect 25496 -22522 25576 -22442
rect 26716 -22522 26796 -22442
rect 26856 -22522 26936 -22442
rect 26996 -22522 27076 -22442
rect 28216 -22522 28296 -22442
rect 28356 -22522 28436 -22442
rect 28496 -22522 28576 -22442
rect 29716 -22502 29776 -22442
rect 29816 -22502 29876 -22442
rect 29956 -22502 30036 -22442
rect 30116 -22502 30176 -22442
rect 30216 -22502 30276 -22442
rect 23516 -22662 23596 -22582
rect 23636 -22662 23696 -22582
rect 23756 -22662 23836 -22582
rect 23896 -22662 23956 -22582
rect 23996 -22662 24076 -22582
rect 25216 -22662 25296 -22582
rect 25356 -22662 25436 -22582
rect 25496 -22662 25576 -22582
rect 26716 -22662 26796 -22582
rect 26856 -22662 26936 -22582
rect 26996 -22662 27076 -22582
rect 28216 -22662 28296 -22582
rect 28356 -22662 28436 -22582
rect 28496 -22662 28576 -22582
rect 29716 -22662 29796 -22582
rect 29836 -22662 29896 -22582
rect 29956 -22662 30036 -22582
rect 30096 -22662 30156 -22582
rect 30196 -22662 30276 -22582
rect 23516 -22802 23576 -22742
rect 23616 -22802 23676 -22742
rect 23756 -22802 23836 -22742
rect 23916 -22802 23976 -22742
rect 24016 -22802 24076 -22742
rect 25216 -22802 25296 -22722
rect 25356 -22802 25436 -22722
rect 25496 -22802 25576 -22722
rect 26716 -22802 26796 -22722
rect 26856 -22802 26936 -22722
rect 26996 -22802 27076 -22722
rect 28216 -22802 28296 -22722
rect 28356 -22802 28436 -22722
rect 28496 -22802 28576 -22722
rect 29716 -22802 29776 -22742
rect 29816 -22802 29876 -22742
rect 29956 -22802 30036 -22742
rect 30116 -22802 30176 -22742
rect 30216 -22802 30276 -22742
rect 20716 -23122 20796 -23062
rect 20836 -23102 20896 -23042
rect 20956 -23122 21036 -23062
rect 21096 -23102 21156 -23042
rect 21196 -23122 21276 -23062
rect 20716 -23222 20796 -23162
rect 20836 -23222 20896 -23162
rect 20956 -23222 21036 -23162
rect 21096 -23222 21156 -23162
rect 21196 -23222 21276 -23162
rect 32516 -23122 32596 -23062
rect 32636 -23102 32696 -23042
rect 32756 -23122 32836 -23062
rect 32896 -23102 32956 -23042
rect 32996 -23122 33076 -23062
rect 32516 -23222 32596 -23162
rect 32636 -23222 32696 -23162
rect 32756 -23222 32836 -23162
rect 32896 -23222 32956 -23162
rect 32996 -23222 33076 -23162
rect 21916 -23522 21976 -23462
rect 22016 -23522 22076 -23462
rect 21916 -23622 21976 -23562
rect 22016 -23622 22076 -23562
rect 24236 -23522 24316 -23442
rect 24356 -23522 24456 -23442
rect 24496 -23522 24576 -23442
rect 24236 -23702 24316 -23622
rect 24356 -23702 24456 -23622
rect 24496 -23702 24576 -23622
rect 25216 -23522 25296 -23442
rect 25336 -23522 25456 -23442
rect 25496 -23522 25576 -23442
rect 25216 -23702 25296 -23622
rect 25336 -23702 25456 -23622
rect 25496 -23702 25576 -23622
rect 28216 -23522 28296 -23442
rect 28336 -23522 28456 -23442
rect 28496 -23522 28576 -23442
rect 28216 -23702 28296 -23622
rect 28336 -23702 28456 -23622
rect 28496 -23702 28576 -23622
rect 29216 -23522 29296 -23442
rect 29336 -23522 29436 -23442
rect 29476 -23522 29556 -23442
rect 29216 -23702 29296 -23622
rect 29336 -23702 29436 -23622
rect 29476 -23702 29556 -23622
rect 31756 -23522 31816 -23462
rect 31856 -23522 31916 -23462
rect 31756 -23622 31816 -23562
rect 31856 -23622 31916 -23562
rect 26436 -24082 26576 -23942
rect 22816 -24202 22896 -24122
rect 22936 -24202 23016 -24122
rect 23056 -24202 23136 -24122
rect 22816 -24302 22876 -24242
rect 22936 -24302 23016 -24242
rect 23076 -24302 23136 -24242
rect 24936 -24202 24996 -24142
rect 25036 -24202 25096 -24142
rect 24696 -24342 24756 -24282
rect 22816 -24422 22896 -24342
rect 22936 -24422 23016 -24342
rect 23056 -24422 23136 -24342
rect 24776 -24422 24836 -24362
rect 27216 -24082 27356 -23942
rect 28696 -24202 28756 -24142
rect 28796 -24202 28856 -24142
rect 29036 -24342 29096 -24282
rect 28956 -24422 29016 -24362
rect 25036 -24582 25096 -24522
rect 24956 -24662 25016 -24602
rect 24696 -24802 24756 -24742
rect 24796 -24802 24856 -24742
rect 21776 -25042 21836 -24982
rect 21896 -25042 21956 -24982
rect 21776 -25222 21836 -25162
rect 21896 -25222 21956 -25162
rect 25216 -25022 25296 -24942
rect 25336 -25022 25456 -24942
rect 25496 -25022 25576 -24942
rect 26436 -25002 26576 -24862
rect 25216 -25202 25296 -25122
rect 25336 -25202 25456 -25122
rect 25496 -25202 25576 -25122
rect 28696 -24582 28756 -24522
rect 30656 -24602 30736 -24522
rect 30776 -24602 30856 -24522
rect 30896 -24602 30976 -24522
rect 28776 -24662 28836 -24602
rect 28936 -24802 28996 -24742
rect 29036 -24802 29096 -24742
rect 30656 -24702 30736 -24642
rect 30776 -24702 30856 -24642
rect 30896 -24702 30976 -24642
rect 30656 -24822 30736 -24742
rect 30776 -24822 30856 -24742
rect 30896 -24822 30976 -24742
rect 27216 -25002 27356 -24862
rect 28216 -25022 28296 -24942
rect 28336 -25022 28456 -24942
rect 28496 -25022 28576 -24942
rect 28216 -25202 28296 -25122
rect 28336 -25202 28456 -25122
rect 28496 -25202 28576 -25122
rect 31836 -25042 31896 -24982
rect 31956 -25042 32016 -24982
rect 31836 -25222 31896 -25162
rect 31956 -25222 32016 -25162
rect 24236 -25622 24316 -25542
rect 24356 -25622 24476 -25542
rect 24516 -25622 24596 -25542
rect 24236 -25802 24316 -25722
rect 24356 -25802 24476 -25722
rect 24516 -25802 24596 -25722
rect 29196 -25622 29276 -25542
rect 29316 -25622 29436 -25542
rect 29476 -25622 29556 -25542
rect 29196 -25802 29276 -25722
rect 29316 -25802 29436 -25722
rect 29476 -25802 29556 -25722
rect 22816 -29122 22896 -29042
rect 22956 -29122 23036 -29042
rect 23096 -29122 23176 -29042
rect 22816 -29262 22896 -29182
rect 22956 -29262 23036 -29182
rect 23096 -29262 23176 -29182
rect 22816 -29402 22896 -29322
rect 22956 -29402 23036 -29322
rect 23096 -29402 23176 -29322
rect 30616 -29122 30696 -29042
rect 30756 -29122 30836 -29042
rect 30896 -29122 30976 -29042
rect 30616 -29262 30696 -29182
rect 30756 -29262 30836 -29182
rect 30896 -29262 30976 -29182
rect 30616 -29402 30696 -29322
rect 30756 -29402 30836 -29322
rect 30896 -29402 30976 -29322
rect 21756 -30502 21816 -30442
rect 21856 -30502 21916 -30442
rect 21956 -30502 22016 -30442
rect 22056 -30502 22116 -30442
rect 21756 -30782 21816 -30722
rect 21856 -30782 21916 -30722
rect 21956 -30782 22016 -30722
rect 22056 -30782 22116 -30722
rect 31676 -30502 31736 -30442
rect 31776 -30502 31836 -30442
rect 31876 -30502 31936 -30442
rect 31976 -30502 32036 -30442
rect 31676 -30782 31736 -30722
rect 31776 -30782 31836 -30722
rect 31876 -30782 31936 -30722
rect 31976 -30782 32036 -30722
<< metal3 >>
rect 200 -10440 14400 3760
rect 39200 1718 53400 3560
rect 39200 -3306 40866 1718
rect 40930 -3306 46478 1718
rect 46542 -3306 53400 1718
rect 39200 -3602 53400 -3306
rect 39200 -8626 40866 -3602
rect 40930 -8626 46478 -3602
rect 46542 -8626 53400 -3602
rect 39200 -10440 53400 -8626
rect 9496 -18930 14868 -18902
rect 9496 -23954 14784 -18930
rect 14848 -23954 14868 -18930
rect 9496 -23982 14868 -23954
rect 15108 -18930 20480 -18902
rect 15108 -23954 20396 -18930
rect 20460 -23954 20480 -18930
rect 33296 -18930 38668 -18902
rect 26696 -21002 27096 -20982
rect 26696 -21082 26716 -21002
rect 26796 -21082 26856 -21002
rect 26936 -21082 26996 -21002
rect 27076 -21082 27096 -21002
rect 26696 -21122 27096 -21082
rect 26696 -21202 26716 -21122
rect 26796 -21202 26856 -21122
rect 26936 -21202 26996 -21122
rect 27076 -21202 27096 -21122
rect 26696 -21262 27096 -21202
rect 26696 -21342 26716 -21262
rect 26796 -21342 26856 -21262
rect 26936 -21342 26996 -21262
rect 27076 -21342 27096 -21262
rect 21736 -21902 22136 -21882
rect 21736 -21962 21776 -21902
rect 21836 -21962 21896 -21902
rect 21976 -21962 22036 -21902
rect 22096 -21962 22136 -21902
rect 21736 -22082 22136 -21962
rect 21736 -22142 21776 -22082
rect 21836 -22142 21896 -22082
rect 21976 -22142 22036 -22082
rect 22096 -22142 22136 -22082
rect 20696 -23042 21296 -23022
rect 20696 -23122 20716 -23042
rect 20796 -23122 20816 -23042
rect 20896 -23122 20956 -23042
rect 21036 -23122 21096 -23042
rect 21176 -23122 21196 -23042
rect 21276 -23122 21296 -23042
rect 20696 -23162 21296 -23122
rect 20696 -23242 20716 -23162
rect 20796 -23242 20816 -23162
rect 20896 -23242 20956 -23162
rect 21036 -23242 21096 -23162
rect 21176 -23242 21196 -23162
rect 21276 -23242 21296 -23162
rect 15108 -23982 20480 -23954
rect 21736 -23462 22136 -22142
rect 24216 -21962 24616 -21942
rect 24216 -22042 24236 -21962
rect 24316 -22042 24376 -21962
rect 24456 -22042 24516 -21962
rect 24596 -22042 24616 -21962
rect 24216 -22102 24616 -22042
rect 24216 -22182 24236 -22102
rect 24316 -22182 24376 -22102
rect 24456 -22182 24516 -22102
rect 24596 -22182 24616 -22102
rect 24216 -22242 24616 -22182
rect 24216 -22322 24236 -22242
rect 24316 -22322 24376 -22242
rect 24456 -22322 24516 -22242
rect 24596 -22322 24616 -22242
rect 23496 -22442 24096 -22422
rect 23496 -22522 23516 -22442
rect 23596 -22522 23616 -22442
rect 23696 -22522 23756 -22442
rect 23836 -22522 23896 -22442
rect 23976 -22522 23996 -22442
rect 24076 -22522 24096 -22442
rect 23496 -22582 24096 -22522
rect 23496 -22662 23516 -22582
rect 23596 -22662 23616 -22582
rect 23696 -22662 23756 -22582
rect 23836 -22662 23896 -22582
rect 23976 -22662 23996 -22582
rect 24076 -22662 24096 -22582
rect 23496 -22722 24096 -22662
rect 23496 -22802 23516 -22722
rect 23596 -22802 23616 -22722
rect 23696 -22802 23756 -22722
rect 23836 -22802 23896 -22722
rect 23976 -22802 23996 -22722
rect 24076 -22802 24096 -22722
rect 23496 -22822 24096 -22802
rect 21736 -23522 21916 -23462
rect 21976 -23522 22016 -23462
rect 22076 -23522 22136 -23462
rect 21736 -23562 22136 -23522
rect 21736 -23622 21916 -23562
rect 21976 -23622 22016 -23562
rect 22076 -23622 22136 -23562
rect 9496 -24250 14868 -24222
rect 9496 -29274 14784 -24250
rect 14848 -29274 14868 -24250
rect 9496 -29302 14868 -29274
rect 15108 -24250 20480 -24222
rect 15108 -29274 20396 -24250
rect 20460 -29274 20480 -24250
rect 15108 -29302 20480 -29274
rect 21736 -24982 22136 -23622
rect 24216 -23442 24616 -22322
rect 24216 -23522 24236 -23442
rect 24316 -23522 24356 -23442
rect 24456 -23522 24496 -23442
rect 24576 -23522 24616 -23442
rect 24216 -23622 24616 -23522
rect 24216 -23702 24236 -23622
rect 24316 -23702 24356 -23622
rect 24456 -23702 24496 -23622
rect 24576 -23702 24616 -23622
rect 21736 -25042 21776 -24982
rect 21836 -25042 21896 -24982
rect 21956 -25042 22136 -24982
rect 21736 -25162 22136 -25042
rect 21736 -25222 21776 -25162
rect 21836 -25222 21896 -25162
rect 21956 -25222 22136 -25162
rect 21736 -30422 22136 -25222
rect 22796 -24122 23156 -24102
rect 22796 -24202 22816 -24122
rect 22896 -24202 22936 -24122
rect 23016 -24202 23056 -24122
rect 23136 -24202 23156 -24122
rect 22796 -24242 23156 -24202
rect 22796 -24302 22816 -24242
rect 22876 -24302 22936 -24242
rect 23016 -24302 23076 -24242
rect 23136 -24262 23156 -24242
rect 23136 -24302 23196 -24262
rect 22796 -24342 23196 -24302
rect 22796 -24422 22816 -24342
rect 22896 -24422 22936 -24342
rect 23016 -24422 23056 -24342
rect 23136 -24422 23196 -24342
rect 22796 -29042 23196 -24422
rect 24216 -25542 24616 -23702
rect 25196 -22442 25596 -22422
rect 25196 -22522 25216 -22442
rect 25296 -22522 25356 -22442
rect 25436 -22522 25496 -22442
rect 25576 -22522 25596 -22442
rect 25196 -22582 25596 -22522
rect 25196 -22662 25216 -22582
rect 25296 -22662 25356 -22582
rect 25436 -22662 25496 -22582
rect 25576 -22662 25596 -22582
rect 25196 -22722 25596 -22662
rect 25196 -22802 25216 -22722
rect 25296 -22802 25356 -22722
rect 25436 -22802 25496 -22722
rect 25576 -22802 25596 -22722
rect 25196 -23442 25596 -22802
rect 26696 -22442 27096 -21342
rect 31656 -21902 32056 -21882
rect 29176 -21962 29576 -21942
rect 29176 -22042 29196 -21962
rect 29276 -22042 29336 -21962
rect 29416 -22042 29476 -21962
rect 29556 -22042 29576 -21962
rect 29176 -22102 29576 -22042
rect 29176 -22182 29196 -22102
rect 29276 -22182 29336 -22102
rect 29416 -22182 29476 -22102
rect 29556 -22182 29576 -22102
rect 29176 -22242 29576 -22182
rect 29176 -22322 29196 -22242
rect 29276 -22322 29336 -22242
rect 29416 -22322 29476 -22242
rect 29556 -22322 29576 -22242
rect 26696 -22522 26716 -22442
rect 26796 -22522 26856 -22442
rect 26936 -22522 26996 -22442
rect 27076 -22522 27096 -22442
rect 26696 -22582 27096 -22522
rect 26696 -22662 26716 -22582
rect 26796 -22662 26856 -22582
rect 26936 -22662 26996 -22582
rect 27076 -22662 27096 -22582
rect 26696 -22722 27096 -22662
rect 26696 -22802 26716 -22722
rect 26796 -22802 26856 -22722
rect 26936 -22802 26996 -22722
rect 27076 -22802 27096 -22722
rect 26696 -22822 27096 -22802
rect 28196 -22442 28596 -22422
rect 28196 -22522 28216 -22442
rect 28296 -22522 28356 -22442
rect 28436 -22522 28496 -22442
rect 28576 -22522 28596 -22442
rect 28196 -22582 28596 -22522
rect 28196 -22662 28216 -22582
rect 28296 -22662 28356 -22582
rect 28436 -22662 28496 -22582
rect 28576 -22662 28596 -22582
rect 28196 -22722 28596 -22662
rect 28196 -22802 28216 -22722
rect 28296 -22802 28356 -22722
rect 28436 -22802 28496 -22722
rect 28576 -22802 28596 -22722
rect 25196 -23522 25216 -23442
rect 25296 -23522 25336 -23442
rect 25456 -23522 25496 -23442
rect 25576 -23522 25596 -23442
rect 25196 -23622 25596 -23522
rect 25196 -23702 25216 -23622
rect 25296 -23702 25336 -23622
rect 25456 -23702 25496 -23622
rect 25576 -23702 25596 -23622
rect 24916 -24142 25116 -24122
rect 24916 -24202 24936 -24142
rect 24996 -24202 25036 -24142
rect 25096 -24202 25116 -24142
rect 24916 -24222 25116 -24202
rect 24676 -24282 24856 -24262
rect 24676 -24342 24696 -24282
rect 24756 -24342 24856 -24282
rect 24676 -24362 24856 -24342
rect 24676 -24422 24776 -24362
rect 24836 -24422 24856 -24362
rect 24676 -24722 24856 -24422
rect 24936 -24522 25116 -24222
rect 24936 -24582 25036 -24522
rect 25096 -24582 25116 -24522
rect 24936 -24602 25116 -24582
rect 24936 -24662 24956 -24602
rect 25016 -24662 25116 -24602
rect 24936 -24682 25116 -24662
rect 24676 -24742 24876 -24722
rect 24676 -24802 24696 -24742
rect 24756 -24802 24796 -24742
rect 24856 -24802 24876 -24742
rect 24676 -24822 24876 -24802
rect 24216 -25622 24236 -25542
rect 24316 -25622 24356 -25542
rect 24476 -25622 24516 -25542
rect 24596 -25622 24616 -25542
rect 24216 -25722 24616 -25622
rect 24216 -25802 24236 -25722
rect 24316 -25802 24356 -25722
rect 24476 -25802 24516 -25722
rect 24596 -25802 24616 -25722
rect 24216 -26122 24616 -25802
rect 25196 -24942 25596 -23702
rect 28196 -23442 28596 -22802
rect 28196 -23522 28216 -23442
rect 28296 -23522 28336 -23442
rect 28456 -23522 28496 -23442
rect 28576 -23522 28596 -23442
rect 28196 -23622 28596 -23522
rect 28196 -23702 28216 -23622
rect 28296 -23702 28336 -23622
rect 28456 -23702 28496 -23622
rect 28576 -23702 28596 -23622
rect 26416 -23942 27376 -23922
rect 26416 -24082 26436 -23942
rect 26576 -24082 27216 -23942
rect 27356 -24082 27376 -23942
rect 26416 -24102 27376 -24082
rect 25196 -25022 25216 -24942
rect 25296 -25022 25336 -24942
rect 25456 -25022 25496 -24942
rect 25576 -25022 25596 -24942
rect 26416 -24862 27376 -24842
rect 26416 -25002 26436 -24862
rect 26576 -25002 27216 -24862
rect 27356 -25002 27376 -24862
rect 26416 -25022 27376 -25002
rect 28196 -24942 28596 -23702
rect 29176 -23442 29576 -22322
rect 31656 -21962 31696 -21902
rect 31756 -21962 31816 -21902
rect 31896 -21962 31956 -21902
rect 32016 -21962 32056 -21902
rect 31656 -22082 32056 -21962
rect 31656 -22142 31696 -22082
rect 31756 -22142 31816 -22082
rect 31896 -22142 31956 -22082
rect 32016 -22142 32056 -22082
rect 29696 -22442 30296 -22422
rect 29696 -22522 29716 -22442
rect 29796 -22522 29816 -22442
rect 29896 -22522 29956 -22442
rect 30036 -22522 30096 -22442
rect 30176 -22522 30196 -22442
rect 30276 -22522 30296 -22442
rect 29696 -22582 30296 -22522
rect 29696 -22662 29716 -22582
rect 29796 -22662 29816 -22582
rect 29896 -22662 29956 -22582
rect 30036 -22662 30096 -22582
rect 30176 -22662 30196 -22582
rect 30276 -22662 30296 -22582
rect 29696 -22722 30296 -22662
rect 29696 -22802 29716 -22722
rect 29796 -22802 29816 -22722
rect 29896 -22802 29956 -22722
rect 30036 -22802 30096 -22722
rect 30176 -22802 30196 -22722
rect 30276 -22802 30296 -22722
rect 29696 -22822 30296 -22802
rect 29176 -23522 29216 -23442
rect 29296 -23522 29336 -23442
rect 29436 -23522 29476 -23442
rect 29556 -23522 29576 -23442
rect 29176 -23622 29576 -23522
rect 29176 -23702 29216 -23622
rect 29296 -23702 29336 -23622
rect 29436 -23702 29476 -23622
rect 29556 -23702 29576 -23622
rect 28676 -24142 28876 -24122
rect 28676 -24202 28696 -24142
rect 28756 -24202 28796 -24142
rect 28856 -24202 28876 -24142
rect 28676 -24222 28876 -24202
rect 28676 -24522 28856 -24222
rect 28676 -24582 28696 -24522
rect 28756 -24582 28856 -24522
rect 28676 -24602 28856 -24582
rect 28676 -24662 28776 -24602
rect 28836 -24662 28856 -24602
rect 28676 -24682 28856 -24662
rect 28936 -24282 29116 -24262
rect 28936 -24342 29036 -24282
rect 29096 -24342 29116 -24282
rect 28936 -24362 29116 -24342
rect 28936 -24422 28956 -24362
rect 29016 -24422 29116 -24362
rect 28936 -24722 29116 -24422
rect 28916 -24742 29116 -24722
rect 28916 -24802 28936 -24742
rect 28996 -24802 29036 -24742
rect 29096 -24802 29116 -24742
rect 28916 -24822 29116 -24802
rect 28196 -25022 28216 -24942
rect 28296 -25022 28336 -24942
rect 28456 -25022 28496 -24942
rect 28576 -25022 28596 -24942
rect 25196 -25122 25596 -25022
rect 25196 -25202 25216 -25122
rect 25296 -25202 25336 -25122
rect 25456 -25202 25496 -25122
rect 25576 -25202 25596 -25122
rect 25196 -26122 25596 -25202
rect 28196 -25122 28596 -25022
rect 28196 -25202 28216 -25122
rect 28296 -25202 28336 -25122
rect 28456 -25202 28496 -25122
rect 28576 -25202 28596 -25122
rect 28196 -26122 28596 -25202
rect 29176 -25542 29576 -23702
rect 31656 -23462 32056 -22142
rect 32496 -23042 33096 -23022
rect 32496 -23122 32516 -23042
rect 32596 -23122 32616 -23042
rect 32696 -23122 32756 -23042
rect 32836 -23122 32896 -23042
rect 32976 -23122 32996 -23042
rect 33076 -23122 33096 -23042
rect 32496 -23162 33096 -23122
rect 32496 -23242 32516 -23162
rect 32596 -23242 32616 -23162
rect 32696 -23242 32756 -23162
rect 32836 -23242 32896 -23162
rect 32976 -23242 32996 -23162
rect 33076 -23242 33096 -23162
rect 31656 -23522 31756 -23462
rect 31816 -23522 31856 -23462
rect 31916 -23522 32056 -23462
rect 31656 -23562 32056 -23522
rect 31656 -23622 31756 -23562
rect 31816 -23622 31856 -23562
rect 31916 -23622 32056 -23562
rect 30636 -24262 30996 -24102
rect 29176 -25622 29196 -25542
rect 29276 -25622 29316 -25542
rect 29436 -25622 29476 -25542
rect 29556 -25622 29576 -25542
rect 29176 -25722 29576 -25622
rect 29176 -25802 29196 -25722
rect 29276 -25802 29316 -25722
rect 29436 -25802 29476 -25722
rect 29556 -25802 29576 -25722
rect 29176 -26122 29576 -25802
rect 30596 -24522 30996 -24262
rect 30596 -24602 30656 -24522
rect 30736 -24602 30776 -24522
rect 30856 -24602 30896 -24522
rect 30976 -24602 30996 -24522
rect 30596 -24642 30996 -24602
rect 30596 -24702 30656 -24642
rect 30736 -24702 30776 -24642
rect 30856 -24702 30896 -24642
rect 30976 -24702 30996 -24642
rect 30596 -24742 30996 -24702
rect 30596 -24822 30656 -24742
rect 30736 -24822 30776 -24742
rect 30856 -24822 30896 -24742
rect 30976 -24822 30996 -24742
rect 22796 -29122 22816 -29042
rect 22896 -29122 22956 -29042
rect 23036 -29122 23096 -29042
rect 23176 -29122 23196 -29042
rect 22796 -29182 23196 -29122
rect 22796 -29262 22816 -29182
rect 22896 -29262 22956 -29182
rect 23036 -29262 23096 -29182
rect 23176 -29262 23196 -29182
rect 22796 -29322 23196 -29262
rect 22796 -29402 22816 -29322
rect 22896 -29402 22956 -29322
rect 23036 -29402 23096 -29322
rect 23176 -29402 23196 -29322
rect 22796 -29422 23196 -29402
rect 30596 -29042 30996 -24822
rect 30596 -29122 30616 -29042
rect 30696 -29122 30756 -29042
rect 30836 -29122 30896 -29042
rect 30976 -29122 30996 -29042
rect 30596 -29182 30996 -29122
rect 30596 -29262 30616 -29182
rect 30696 -29262 30756 -29182
rect 30836 -29262 30896 -29182
rect 30976 -29262 30996 -29182
rect 30596 -29322 30996 -29262
rect 30596 -29402 30616 -29322
rect 30696 -29402 30756 -29322
rect 30836 -29402 30896 -29322
rect 30976 -29402 30996 -29322
rect 30596 -29422 30996 -29402
rect 31656 -24982 32056 -23622
rect 33296 -23954 33316 -18930
rect 33380 -23954 38668 -18930
rect 33296 -23982 38668 -23954
rect 38908 -18930 44280 -18902
rect 38908 -23954 38928 -18930
rect 38992 -23954 44280 -18930
rect 38908 -23982 44280 -23954
rect 31656 -25042 31836 -24982
rect 31896 -25042 31956 -24982
rect 32016 -25042 32056 -24982
rect 31656 -25162 32056 -25042
rect 31656 -25222 31836 -25162
rect 31896 -25222 31956 -25162
rect 32016 -25222 32056 -25162
rect 31656 -30422 32056 -25222
rect 33296 -24250 38668 -24222
rect 33296 -29274 33316 -24250
rect 33380 -29274 38668 -24250
rect 33296 -29302 38668 -29274
rect 38908 -24250 44280 -24222
rect 38908 -29274 38928 -24250
rect 38992 -29274 44280 -24250
rect 38908 -29302 44280 -29274
rect 21736 -30442 32056 -30422
rect 21736 -30502 21756 -30442
rect 21816 -30502 21856 -30442
rect 21916 -30502 21956 -30442
rect 22016 -30502 22056 -30442
rect 22116 -30502 31676 -30442
rect 31736 -30502 31776 -30442
rect 31836 -30502 31876 -30442
rect 31936 -30502 31976 -30442
rect 32036 -30502 32056 -30442
rect 21736 -30722 32056 -30502
rect 21736 -30782 21756 -30722
rect 21816 -30782 21856 -30722
rect 21916 -30782 21956 -30722
rect 22016 -30782 22056 -30722
rect 22116 -30782 31676 -30722
rect 31736 -30782 31776 -30722
rect 31836 -30782 31876 -30722
rect 31936 -30782 31976 -30722
rect 32036 -30782 32056 -30722
rect 21736 -30802 32056 -30782
<< via3 >>
rect 40866 -3306 40930 1718
rect 46478 -3306 46542 1718
rect 40866 -8626 40930 -3602
rect 46478 -8626 46542 -3602
rect 14784 -23954 14848 -18930
rect 20396 -23954 20460 -18930
rect 20716 -23062 20796 -23042
rect 20716 -23122 20796 -23062
rect 20816 -23102 20836 -23042
rect 20836 -23102 20896 -23042
rect 20816 -23122 20896 -23102
rect 20956 -23062 21036 -23042
rect 20956 -23122 21036 -23062
rect 21096 -23102 21156 -23042
rect 21156 -23102 21176 -23042
rect 21096 -23122 21176 -23102
rect 21196 -23062 21276 -23042
rect 21196 -23122 21276 -23062
rect 20716 -23222 20796 -23162
rect 20716 -23242 20796 -23222
rect 20816 -23222 20836 -23162
rect 20836 -23222 20896 -23162
rect 20816 -23242 20896 -23222
rect 20956 -23222 21036 -23162
rect 20956 -23242 21036 -23222
rect 21096 -23222 21156 -23162
rect 21156 -23222 21176 -23162
rect 21096 -23242 21176 -23222
rect 21196 -23222 21276 -23162
rect 21196 -23242 21276 -23222
rect 23516 -22502 23576 -22442
rect 23576 -22502 23596 -22442
rect 23516 -22522 23596 -22502
rect 23616 -22502 23676 -22442
rect 23676 -22502 23696 -22442
rect 23616 -22522 23696 -22502
rect 23756 -22502 23836 -22442
rect 23756 -22522 23836 -22502
rect 23896 -22502 23916 -22442
rect 23916 -22502 23976 -22442
rect 23896 -22522 23976 -22502
rect 23996 -22502 24016 -22442
rect 24016 -22502 24076 -22442
rect 23996 -22522 24076 -22502
rect 23516 -22662 23596 -22582
rect 23616 -22662 23636 -22582
rect 23636 -22662 23696 -22582
rect 23756 -22662 23836 -22582
rect 23896 -22662 23956 -22582
rect 23956 -22662 23976 -22582
rect 23996 -22662 24076 -22582
rect 23516 -22742 23596 -22722
rect 23516 -22802 23576 -22742
rect 23576 -22802 23596 -22742
rect 23616 -22742 23696 -22722
rect 23616 -22802 23676 -22742
rect 23676 -22802 23696 -22742
rect 23756 -22742 23836 -22722
rect 23756 -22802 23836 -22742
rect 23896 -22742 23976 -22722
rect 23896 -22802 23916 -22742
rect 23916 -22802 23976 -22742
rect 23996 -22742 24076 -22722
rect 23996 -22802 24016 -22742
rect 24016 -22802 24076 -22742
rect 14784 -29274 14848 -24250
rect 20396 -29274 20460 -24250
rect 29716 -22502 29776 -22442
rect 29776 -22502 29796 -22442
rect 29716 -22522 29796 -22502
rect 29816 -22502 29876 -22442
rect 29876 -22502 29896 -22442
rect 29816 -22522 29896 -22502
rect 29956 -22502 30036 -22442
rect 29956 -22522 30036 -22502
rect 30096 -22502 30116 -22442
rect 30116 -22502 30176 -22442
rect 30096 -22522 30176 -22502
rect 30196 -22502 30216 -22442
rect 30216 -22502 30276 -22442
rect 30196 -22522 30276 -22502
rect 29716 -22662 29796 -22582
rect 29816 -22662 29836 -22582
rect 29836 -22662 29896 -22582
rect 29956 -22662 30036 -22582
rect 30096 -22662 30156 -22582
rect 30156 -22662 30176 -22582
rect 30196 -22662 30276 -22582
rect 29716 -22742 29796 -22722
rect 29716 -22802 29776 -22742
rect 29776 -22802 29796 -22742
rect 29816 -22742 29896 -22722
rect 29816 -22802 29876 -22742
rect 29876 -22802 29896 -22742
rect 29956 -22742 30036 -22722
rect 29956 -22802 30036 -22742
rect 30096 -22742 30176 -22722
rect 30096 -22802 30116 -22742
rect 30116 -22802 30176 -22742
rect 30196 -22742 30276 -22722
rect 30196 -22802 30216 -22742
rect 30216 -22802 30276 -22742
rect 32516 -23062 32596 -23042
rect 32516 -23122 32596 -23062
rect 32616 -23102 32636 -23042
rect 32636 -23102 32696 -23042
rect 32616 -23122 32696 -23102
rect 32756 -23062 32836 -23042
rect 32756 -23122 32836 -23062
rect 32896 -23102 32956 -23042
rect 32956 -23102 32976 -23042
rect 32896 -23122 32976 -23102
rect 32996 -23062 33076 -23042
rect 32996 -23122 33076 -23062
rect 32516 -23222 32596 -23162
rect 32516 -23242 32596 -23222
rect 32616 -23222 32636 -23162
rect 32636 -23222 32696 -23162
rect 32616 -23242 32696 -23222
rect 32756 -23222 32836 -23162
rect 32756 -23242 32836 -23222
rect 32896 -23222 32956 -23162
rect 32956 -23222 32976 -23162
rect 32896 -23242 32976 -23222
rect 32996 -23222 33076 -23162
rect 32996 -23242 33076 -23222
rect 33316 -23954 33380 -18930
rect 38928 -23954 38992 -18930
rect 33316 -29274 33380 -24250
rect 38928 -29274 38992 -24250
<< mimcap >>
rect 41178 1666 46178 1706
rect 41178 -3254 41218 1666
rect 46138 -3254 46178 1666
rect 41178 -3294 46178 -3254
rect 46790 1666 51790 1706
rect 46790 -3254 46830 1666
rect 51750 -3254 51790 1666
rect 46790 -3294 51790 -3254
rect 41178 -3654 46178 -3614
rect 41178 -8574 41218 -3654
rect 46138 -8574 46178 -3654
rect 41178 -8614 46178 -8574
rect 46790 -3654 51790 -3614
rect 46790 -8574 46830 -3654
rect 51750 -8574 51790 -3654
rect 46790 -8614 51790 -8574
rect 9536 -18982 14536 -18942
rect 9536 -23902 9576 -18982
rect 14496 -23902 14536 -18982
rect 9536 -23942 14536 -23902
rect 15148 -18982 20148 -18942
rect 15148 -23902 15188 -18982
rect 20108 -23902 20148 -18982
rect 15148 -23942 20148 -23902
rect 33628 -18982 38628 -18942
rect 33628 -23902 33668 -18982
rect 38588 -23902 38628 -18982
rect 33628 -23942 38628 -23902
rect 39240 -18982 44240 -18942
rect 39240 -23902 39280 -18982
rect 44200 -23902 44240 -18982
rect 39240 -23942 44240 -23902
rect 9536 -24302 14536 -24262
rect 9536 -29222 9576 -24302
rect 14496 -29222 14536 -24302
rect 9536 -29262 14536 -29222
rect 15148 -24302 20148 -24262
rect 15148 -29222 15188 -24302
rect 20108 -29222 20148 -24302
rect 15148 -29262 20148 -29222
rect 33628 -24302 38628 -24262
rect 33628 -29222 33668 -24302
rect 38588 -29222 38628 -24302
rect 33628 -29262 38628 -29222
rect 39240 -24302 44240 -24262
rect 39240 -29222 39280 -24302
rect 44200 -29222 44240 -24302
rect 39240 -29262 44240 -29222
<< mimcapcontact >>
rect 41218 -3254 46138 1666
rect 46830 -3254 51750 1666
rect 41218 -8574 46138 -3654
rect 46830 -8574 51750 -3654
rect 9576 -23902 14496 -18982
rect 15188 -23902 20108 -18982
rect 33668 -23902 38588 -18982
rect 39280 -23902 44200 -18982
rect 9576 -29222 14496 -24302
rect 15188 -29222 20108 -24302
rect 33668 -29222 38588 -24302
rect 39280 -29222 44200 -24302
<< metal4 >>
rect 40846 1718 40950 1866
rect 40846 -3306 40866 1718
rect 40930 -3306 40950 1718
rect 43626 1667 43730 1866
rect 46458 1718 46562 1866
rect 41217 1666 46139 1667
rect 41217 -3254 41218 1666
rect 46138 -3254 46139 1666
rect 41217 -3255 46139 -3254
rect 40846 -3602 40950 -3306
rect 40846 -8626 40866 -3602
rect 40930 -8626 40950 -3602
rect 43626 -3653 43730 -3255
rect 46458 -3306 46478 1718
rect 46542 -3306 46562 1718
rect 49238 1667 49342 1866
rect 46829 1666 51751 1667
rect 46829 -3254 46830 1666
rect 51750 -3254 51751 1666
rect 46829 -3255 51751 -3254
rect 46458 -3602 46562 -3306
rect 41217 -3654 46139 -3653
rect 41217 -8574 41218 -3654
rect 46138 -8574 46139 -3654
rect 41217 -8575 46139 -8574
rect 40846 -8774 40950 -8626
rect 43626 -8774 43730 -8575
rect 46458 -8626 46478 -3602
rect 46542 -8626 46562 -3602
rect 49238 -3653 49342 -3255
rect 46829 -3654 51751 -3653
rect 46829 -8574 46830 -3654
rect 51750 -8574 51751 -3654
rect 46829 -8575 51751 -8574
rect 46458 -8774 46562 -8626
rect 49238 -8774 49342 -8575
rect 6000 -32000 8000 -10000
rect 14696 -18622 39096 -18022
rect 11984 -18981 12088 -18782
rect 14696 -18822 14936 -18622
rect 20296 -18782 20536 -18622
rect 14764 -18930 14868 -18822
rect 9575 -18982 14497 -18981
rect 9575 -23902 9576 -18982
rect 14496 -23902 14497 -18982
rect 9575 -23903 14497 -23902
rect 11984 -24301 12088 -23903
rect 14764 -23954 14784 -18930
rect 14848 -23954 14868 -18930
rect 17596 -18981 17700 -18782
rect 20376 -18930 20480 -18782
rect 15187 -18982 20109 -18981
rect 15187 -23902 15188 -18982
rect 20108 -23902 20109 -18982
rect 15187 -23903 20109 -23902
rect 14764 -24250 14868 -23954
rect 9575 -24302 14497 -24301
rect 9575 -29222 9576 -24302
rect 14496 -29222 14497 -24302
rect 9575 -29223 14497 -29222
rect 11984 -29422 12088 -29223
rect 14764 -29274 14784 -24250
rect 14848 -29274 14868 -24250
rect 17596 -24301 17700 -23903
rect 20376 -23954 20396 -18930
rect 20460 -23954 20480 -18930
rect 23496 -22442 24096 -18622
rect 23496 -22522 23516 -22442
rect 23596 -22522 23616 -22442
rect 23696 -22522 23756 -22442
rect 23836 -22522 23896 -22442
rect 23976 -22522 23996 -22442
rect 24076 -22522 24096 -22442
rect 23496 -22582 24096 -22522
rect 23496 -22662 23516 -22582
rect 23596 -22662 23616 -22582
rect 23696 -22662 23756 -22582
rect 23836 -22662 23896 -22582
rect 23976 -22662 23996 -22582
rect 24076 -22662 24096 -22582
rect 23496 -22722 24096 -22662
rect 23496 -22802 23516 -22722
rect 23596 -22802 23616 -22722
rect 23696 -22802 23756 -22722
rect 23836 -22802 23896 -22722
rect 23976 -22802 23996 -22722
rect 24076 -22802 24096 -22722
rect 23496 -22822 24096 -22802
rect 29696 -22442 30296 -18622
rect 33216 -18782 33456 -18622
rect 38856 -18782 39096 -18622
rect 29696 -22522 29716 -22442
rect 29796 -22522 29816 -22442
rect 29896 -22522 29956 -22442
rect 30036 -22522 30096 -22442
rect 30176 -22522 30196 -22442
rect 30276 -22522 30296 -22442
rect 29696 -22582 30296 -22522
rect 29696 -22662 29716 -22582
rect 29796 -22662 29816 -22582
rect 29896 -22662 29956 -22582
rect 30036 -22662 30096 -22582
rect 30176 -22662 30196 -22582
rect 30276 -22662 30296 -22582
rect 29696 -22722 30296 -22662
rect 29696 -22802 29716 -22722
rect 29796 -22802 29816 -22722
rect 29896 -22802 29956 -22722
rect 30036 -22802 30096 -22722
rect 30176 -22802 30196 -22722
rect 30276 -22802 30296 -22722
rect 29696 -22822 30296 -22802
rect 33296 -18930 33400 -18782
rect 20376 -24250 20480 -23954
rect 15187 -24302 20109 -24301
rect 15187 -29222 15188 -24302
rect 20108 -29222 20109 -24302
rect 15187 -29223 20109 -29222
rect 14764 -29422 14868 -29274
rect 17596 -29422 17700 -29223
rect 20376 -29274 20396 -24250
rect 20460 -29274 20480 -24250
rect 20376 -29422 20480 -29274
rect 20696 -23042 21296 -23022
rect 20696 -23122 20716 -23042
rect 20796 -23122 20816 -23042
rect 20896 -23122 20956 -23042
rect 21036 -23122 21096 -23042
rect 21176 -23122 21196 -23042
rect 21276 -23122 21296 -23042
rect 20696 -23162 21296 -23122
rect 20696 -23242 20716 -23162
rect 20796 -23242 20816 -23162
rect 20896 -23242 20956 -23162
rect 21036 -23242 21096 -23162
rect 21176 -23242 21196 -23162
rect 21276 -23242 21296 -23162
rect 11896 -29622 12176 -29422
rect 17516 -29622 17776 -29422
rect 20696 -29622 21296 -23242
rect 32496 -23042 33096 -23022
rect 32496 -23122 32516 -23042
rect 32596 -23122 32616 -23042
rect 32696 -23122 32756 -23042
rect 32836 -23122 32896 -23042
rect 32976 -23122 32996 -23042
rect 33076 -23122 33096 -23042
rect 32496 -23162 33096 -23122
rect 32496 -23242 32516 -23162
rect 32596 -23242 32616 -23162
rect 32696 -23242 32756 -23162
rect 32836 -23242 32896 -23162
rect 32976 -23242 32996 -23162
rect 33076 -23242 33096 -23162
rect 32496 -29622 33096 -23242
rect 33296 -23954 33316 -18930
rect 33380 -23954 33400 -18930
rect 36076 -18981 36180 -18782
rect 38908 -18930 39012 -18782
rect 33667 -18982 38589 -18981
rect 33667 -23902 33668 -18982
rect 38588 -23902 38589 -18982
rect 33667 -23903 38589 -23902
rect 33296 -24250 33400 -23954
rect 33296 -29274 33316 -24250
rect 33380 -29274 33400 -24250
rect 36076 -24301 36180 -23903
rect 38908 -23954 38928 -18930
rect 38992 -23954 39012 -18930
rect 41688 -18981 41792 -18782
rect 39279 -18982 44201 -18981
rect 39279 -23902 39280 -18982
rect 44200 -23902 44201 -18982
rect 39279 -23903 44201 -23902
rect 38908 -24250 39012 -23954
rect 33667 -24302 38589 -24301
rect 33667 -29222 33668 -24302
rect 38588 -29222 38589 -24302
rect 33667 -29223 38589 -29222
rect 33296 -29422 33400 -29274
rect 36076 -29402 36180 -29223
rect 38908 -29274 38928 -24250
rect 38992 -29274 39012 -24250
rect 41688 -24301 41792 -23903
rect 39279 -24302 44201 -24301
rect 39279 -29222 39280 -24302
rect 44200 -29222 44201 -24302
rect 39279 -29223 44201 -29222
rect 35996 -29622 36256 -29402
rect 38908 -29422 39012 -29274
rect 41688 -29402 41792 -29223
rect 41616 -29622 41896 -29402
rect 11896 -30222 41896 -29622
rect 46000 -32000 48000 -10000
rect 6000 -34000 22000 -32000
rect 26000 -46000 28000 -32000
rect 32000 -34000 48000 -32000
<< metal5 >>
rect 4000 6000 50000 10000
rect 4000 -16000 50000 -12000
rect 4000 -38000 50000 -34000
use 1st-stage  1st-stage_1 error-amplifier2/layout
timestamp 1770370310
transform 1 0 13496 0 1 -19022
box -4000 -11780 30784 1000
use serpentine259k  serpentine259k_0 serpentine259k/topology2
timestamp 1770177229
transform 1 0 57500 0 1 26500
box -1500 -72500 10000 -5500
use serpentine259k  serpentine259k_1
timestamp 1770177229
transform 1 0 -12500 0 1 26500
box -1500 -72500 10000 -5500
use sky130_fd_pr__cap_mim_m3_1_RK594X  sky130_fd_pr__cap_mim_m3_1_RK594X_1 error-amplifier2/layout
timestamp 1770370310
transform -1 0 46338 0 -1 -3454
box -5492 -5320 5492 5320
use sky130_fd_pr__cap_mim_m3_1_RK594X  XC2
timestamp 1770370310
transform 1 0 7262 0 1 -3426
box -5492 -5320 5492 5320
use sky130_fd_pr__pfet_g5v0d10v5_YYQDC9  XM1
timestamp 1770370310
transform 1 0 27285 0 1 1328
box -5285 -1328 5285 1328
use sky130_fd_pr__nfet_g5v0d10v5_MLLFC6  XM3
timestamp 1770370310
transform 1 0 26711 0 1 -7582
box -10311 -2258 10311 2258
<< labels >>
flabel metal1 21836 -30702 22036 -30502 0 FreeSans 800 0 0 0 OUT
port 14 nsew
flabel metal1 26796 -29922 26996 -29722 0 FreeSans 256 0 0 0 IBIAS
port 9 nsew
flabel metal1 30696 -29322 30896 -29122 0 FreeSans 256 0 0 0 VN
port 4 nsew
flabel metal1 22896 -29322 23096 -29122 0 FreeSans 256 0 0 0 VP
port 3 nsew
flabel metal1 27896 -28722 28096 -28522 0 FreeSans 256 0 0 0 VSS
port 11 nsew
flabel metal1 26416 -19202 26616 -19002 0 FreeSans 800 0 0 0 VDD
port 17 nsew
<< end >>
