magic
tech sky130A
magscale 1 2
timestamp 1769170054
<< nwell >>
rect -1461 -767 1461 767
<< mvpmos >>
rect -1203 -470 -953 470
rect -895 -470 -645 470
rect -587 -470 -337 470
rect -279 -470 -29 470
rect 29 -470 279 470
rect 337 -470 587 470
rect 645 -470 895 470
rect 953 -470 1203 470
<< mvpdiff >>
rect -1261 458 -1203 470
rect -1261 -458 -1249 458
rect -1215 -458 -1203 458
rect -1261 -470 -1203 -458
rect -953 458 -895 470
rect -953 -458 -941 458
rect -907 -458 -895 458
rect -953 -470 -895 -458
rect -645 458 -587 470
rect -645 -458 -633 458
rect -599 -458 -587 458
rect -645 -470 -587 -458
rect -337 458 -279 470
rect -337 -458 -325 458
rect -291 -458 -279 458
rect -337 -470 -279 -458
rect -29 458 29 470
rect -29 -458 -17 458
rect 17 -458 29 458
rect -29 -470 29 -458
rect 279 458 337 470
rect 279 -458 291 458
rect 325 -458 337 458
rect 279 -470 337 -458
rect 587 458 645 470
rect 587 -458 599 458
rect 633 -458 645 458
rect 587 -470 645 -458
rect 895 458 953 470
rect 895 -458 907 458
rect 941 -458 953 458
rect 895 -470 953 -458
rect 1203 458 1261 470
rect 1203 -458 1215 458
rect 1249 -458 1261 458
rect 1203 -470 1261 -458
<< mvpdiffc >>
rect -1249 -458 -1215 458
rect -941 -458 -907 458
rect -633 -458 -599 458
rect -325 -458 -291 458
rect -17 -458 17 458
rect 291 -458 325 458
rect 599 -458 633 458
rect 907 -458 941 458
rect 1215 -458 1249 458
<< mvnsubdiff >>
rect -1395 689 1395 701
rect -1395 655 -1287 689
rect 1287 655 1395 689
rect -1395 643 1395 655
rect -1395 593 -1337 643
rect -1395 -593 -1383 593
rect -1349 -593 -1337 593
rect 1337 593 1395 643
rect -1395 -643 -1337 -593
rect 1337 -593 1349 593
rect 1383 -593 1395 593
rect 1337 -643 1395 -593
rect -1395 -655 1395 -643
rect -1395 -689 -1287 -655
rect 1287 -689 1395 -655
rect -1395 -701 1395 -689
<< mvnsubdiffcont >>
rect -1287 655 1287 689
rect -1383 -593 -1349 593
rect 1349 -593 1383 593
rect -1287 -689 1287 -655
<< poly >>
rect -1203 551 -953 567
rect -1203 517 -1187 551
rect -969 517 -953 551
rect -1203 470 -953 517
rect -895 551 -645 567
rect -895 517 -879 551
rect -661 517 -645 551
rect -895 470 -645 517
rect -587 551 -337 567
rect -587 517 -571 551
rect -353 517 -337 551
rect -587 470 -337 517
rect -279 551 -29 567
rect -279 517 -263 551
rect -45 517 -29 551
rect -279 470 -29 517
rect 29 551 279 567
rect 29 517 45 551
rect 263 517 279 551
rect 29 470 279 517
rect 337 551 587 567
rect 337 517 353 551
rect 571 517 587 551
rect 337 470 587 517
rect 645 551 895 567
rect 645 517 661 551
rect 879 517 895 551
rect 645 470 895 517
rect 953 551 1203 567
rect 953 517 969 551
rect 1187 517 1203 551
rect 953 470 1203 517
rect -1203 -517 -953 -470
rect -1203 -551 -1187 -517
rect -969 -551 -953 -517
rect -1203 -567 -953 -551
rect -895 -517 -645 -470
rect -895 -551 -879 -517
rect -661 -551 -645 -517
rect -895 -567 -645 -551
rect -587 -517 -337 -470
rect -587 -551 -571 -517
rect -353 -551 -337 -517
rect -587 -567 -337 -551
rect -279 -517 -29 -470
rect -279 -551 -263 -517
rect -45 -551 -29 -517
rect -279 -567 -29 -551
rect 29 -517 279 -470
rect 29 -551 45 -517
rect 263 -551 279 -517
rect 29 -567 279 -551
rect 337 -517 587 -470
rect 337 -551 353 -517
rect 571 -551 587 -517
rect 337 -567 587 -551
rect 645 -517 895 -470
rect 645 -551 661 -517
rect 879 -551 895 -517
rect 645 -567 895 -551
rect 953 -517 1203 -470
rect 953 -551 969 -517
rect 1187 -551 1203 -517
rect 953 -567 1203 -551
<< polycont >>
rect -1187 517 -969 551
rect -879 517 -661 551
rect -571 517 -353 551
rect -263 517 -45 551
rect 45 517 263 551
rect 353 517 571 551
rect 661 517 879 551
rect 969 517 1187 551
rect -1187 -551 -969 -517
rect -879 -551 -661 -517
rect -571 -551 -353 -517
rect -263 -551 -45 -517
rect 45 -551 263 -517
rect 353 -551 571 -517
rect 661 -551 879 -517
rect 969 -551 1187 -517
<< locali >>
rect -1383 655 -1287 689
rect 1287 655 1383 689
rect -1383 593 -1349 655
rect 1349 593 1383 655
rect -1203 517 -1187 551
rect -969 517 -953 551
rect -895 517 -879 551
rect -661 517 -645 551
rect -587 517 -571 551
rect -353 517 -337 551
rect -279 517 -263 551
rect -45 517 -29 551
rect 29 517 45 551
rect 263 517 279 551
rect 337 517 353 551
rect 571 517 587 551
rect 645 517 661 551
rect 879 517 895 551
rect 953 517 969 551
rect 1187 517 1203 551
rect -1249 458 -1215 474
rect -1249 -474 -1215 -458
rect -941 458 -907 474
rect -941 -474 -907 -458
rect -633 458 -599 474
rect -633 -474 -599 -458
rect -325 458 -291 474
rect -325 -474 -291 -458
rect -17 458 17 474
rect -17 -474 17 -458
rect 291 458 325 474
rect 291 -474 325 -458
rect 599 458 633 474
rect 599 -474 633 -458
rect 907 458 941 474
rect 907 -474 941 -458
rect 1215 458 1249 474
rect 1215 -474 1249 -458
rect -1203 -551 -1187 -517
rect -969 -551 -953 -517
rect -895 -551 -879 -517
rect -661 -551 -645 -517
rect -587 -551 -571 -517
rect -353 -551 -337 -517
rect -279 -551 -263 -517
rect -45 -551 -29 -517
rect 29 -551 45 -517
rect 263 -551 279 -517
rect 337 -551 353 -517
rect 571 -551 587 -517
rect 645 -551 661 -517
rect 879 -551 895 -517
rect 953 -551 969 -517
rect 1187 -551 1203 -517
rect -1383 -655 -1349 -593
rect 1349 -655 1383 -593
rect -1383 -689 -1287 -655
rect 1287 -689 1383 -655
<< viali >>
rect -1187 517 -969 551
rect -879 517 -661 551
rect -571 517 -353 551
rect -263 517 -45 551
rect 45 517 263 551
rect 353 517 571 551
rect 661 517 879 551
rect 969 517 1187 551
rect -1249 -458 -1215 458
rect -941 -458 -907 458
rect -633 -458 -599 458
rect -325 -458 -291 458
rect -17 -458 17 458
rect 291 -458 325 458
rect 599 -458 633 458
rect 907 -458 941 458
rect 1215 -458 1249 458
rect -1187 -551 -969 -517
rect -879 -551 -661 -517
rect -571 -551 -353 -517
rect -263 -551 -45 -517
rect 45 -551 263 -517
rect 353 -551 571 -517
rect 661 -551 879 -517
rect 969 -551 1187 -517
<< metal1 >>
rect -1199 551 -957 557
rect -1199 517 -1187 551
rect -969 517 -957 551
rect -1199 511 -957 517
rect -891 551 -649 557
rect -891 517 -879 551
rect -661 517 -649 551
rect -891 511 -649 517
rect -583 551 -341 557
rect -583 517 -571 551
rect -353 517 -341 551
rect -583 511 -341 517
rect -275 551 -33 557
rect -275 517 -263 551
rect -45 517 -33 551
rect -275 511 -33 517
rect 33 551 275 557
rect 33 517 45 551
rect 263 517 275 551
rect 33 511 275 517
rect 341 551 583 557
rect 341 517 353 551
rect 571 517 583 551
rect 341 511 583 517
rect 649 551 891 557
rect 649 517 661 551
rect 879 517 891 551
rect 649 511 891 517
rect 957 551 1199 557
rect 957 517 969 551
rect 1187 517 1199 551
rect 957 511 1199 517
rect -1255 458 -1209 470
rect -1255 -458 -1249 458
rect -1215 -458 -1209 458
rect -1255 -470 -1209 -458
rect -947 458 -901 470
rect -947 -458 -941 458
rect -907 -458 -901 458
rect -947 -470 -901 -458
rect -639 458 -593 470
rect -639 -458 -633 458
rect -599 -458 -593 458
rect -639 -470 -593 -458
rect -331 458 -285 470
rect -331 -458 -325 458
rect -291 -458 -285 458
rect -331 -470 -285 -458
rect -23 458 23 470
rect -23 -458 -17 458
rect 17 -458 23 458
rect -23 -470 23 -458
rect 285 458 331 470
rect 285 -458 291 458
rect 325 -458 331 458
rect 285 -470 331 -458
rect 593 458 639 470
rect 593 -458 599 458
rect 633 -458 639 458
rect 593 -470 639 -458
rect 901 458 947 470
rect 901 -458 907 458
rect 941 -458 947 458
rect 901 -470 947 -458
rect 1209 458 1255 470
rect 1209 -458 1215 458
rect 1249 -458 1255 458
rect 1209 -470 1255 -458
rect -1199 -517 -957 -511
rect -1199 -551 -1187 -517
rect -969 -551 -957 -517
rect -1199 -557 -957 -551
rect -891 -517 -649 -511
rect -891 -551 -879 -517
rect -661 -551 -649 -517
rect -891 -557 -649 -551
rect -583 -517 -341 -511
rect -583 -551 -571 -517
rect -353 -551 -341 -517
rect -583 -557 -341 -551
rect -275 -517 -33 -511
rect -275 -551 -263 -517
rect -45 -551 -33 -517
rect -275 -557 -33 -551
rect 33 -517 275 -511
rect 33 -551 45 -517
rect 263 -551 275 -517
rect 33 -557 275 -551
rect 341 -517 583 -511
rect 341 -551 353 -517
rect 571 -551 583 -517
rect 341 -557 583 -551
rect 649 -517 891 -511
rect 649 -551 661 -517
rect 879 -551 891 -517
rect 649 -557 891 -551
rect 957 -517 1199 -511
rect 957 -551 969 -517
rect 1187 -551 1199 -517
rect 957 -557 1199 -551
<< properties >>
string FIXED_BBOX -1366 -672 1366 672
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.7 l 1.25 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
