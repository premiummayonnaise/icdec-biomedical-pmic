magic
tech sky130A
magscale 1 2
timestamp 1769412267
<< error_p >>
rect -1112 791 -1044 797
rect -804 791 -736 797
rect -496 791 -428 797
rect -188 791 -120 797
rect 120 791 188 797
rect 428 791 496 797
rect 736 791 804 797
rect 1044 791 1112 797
rect -1112 757 -1100 791
rect -804 757 -792 791
rect -496 757 -484 791
rect -188 757 -176 791
rect 120 757 132 791
rect 428 757 440 791
rect 736 757 748 791
rect 1044 757 1056 791
rect -1112 751 -1044 757
rect -804 751 -736 757
rect -496 751 -428 757
rect -188 751 -120 757
rect 120 751 188 757
rect 428 751 496 757
rect 736 751 804 757
rect 1044 751 1112 757
<< mvnmos >>
rect -1203 -781 -953 719
rect -895 -781 -645 719
rect -587 -781 -337 719
rect -279 -781 -29 719
rect 29 -781 279 719
rect 337 -781 587 719
rect 645 -781 895 719
rect 953 -781 1203 719
<< mvndiff >>
rect -1261 707 -1203 719
rect -1261 -769 -1249 707
rect -1215 -769 -1203 707
rect -1261 -781 -1203 -769
rect -953 707 -895 719
rect -953 -769 -941 707
rect -907 -769 -895 707
rect -953 -781 -895 -769
rect -645 707 -587 719
rect -645 -769 -633 707
rect -599 -769 -587 707
rect -645 -781 -587 -769
rect -337 707 -279 719
rect -337 -769 -325 707
rect -291 -769 -279 707
rect -337 -781 -279 -769
rect -29 707 29 719
rect -29 -769 -17 707
rect 17 -769 29 707
rect -29 -781 29 -769
rect 279 707 337 719
rect 279 -769 291 707
rect 325 -769 337 707
rect 279 -781 337 -769
rect 587 707 645 719
rect 587 -769 599 707
rect 633 -769 645 707
rect 587 -781 645 -769
rect 895 707 953 719
rect 895 -769 907 707
rect 941 -769 953 707
rect 895 -781 953 -769
rect 1203 707 1261 719
rect 1203 -769 1215 707
rect 1249 -769 1261 707
rect 1203 -781 1261 -769
<< mvndiffc >>
rect -1249 -769 -1215 707
rect -941 -769 -907 707
rect -633 -769 -599 707
rect -325 -769 -291 707
rect -17 -769 17 707
rect 291 -769 325 707
rect 599 -769 633 707
rect 907 -769 941 707
rect 1215 -769 1249 707
<< poly >>
rect -1116 791 -1040 807
rect -1116 774 -1100 791
rect -1203 757 -1100 774
rect -1056 774 -1040 791
rect -808 791 -732 807
rect -808 774 -792 791
rect -1056 757 -953 774
rect -1203 719 -953 757
rect -895 757 -792 774
rect -748 774 -732 791
rect -500 791 -424 807
rect -500 774 -484 791
rect -748 757 -645 774
rect -895 719 -645 757
rect -587 757 -484 774
rect -440 774 -424 791
rect -192 791 -116 807
rect -192 774 -176 791
rect -440 757 -337 774
rect -587 719 -337 757
rect -279 757 -176 774
rect -132 774 -116 791
rect 116 791 192 807
rect 116 774 132 791
rect -132 757 -29 774
rect -279 719 -29 757
rect 29 757 132 774
rect 176 774 192 791
rect 424 791 500 807
rect 424 774 440 791
rect 176 757 279 774
rect 29 719 279 757
rect 337 757 440 774
rect 484 774 500 791
rect 732 791 808 807
rect 732 774 748 791
rect 484 757 587 774
rect 337 719 587 757
rect 645 757 748 774
rect 792 774 808 791
rect 1040 791 1116 807
rect 1040 774 1056 791
rect 792 757 895 774
rect 645 719 895 757
rect 953 757 1056 774
rect 1100 774 1116 791
rect 1100 757 1203 774
rect 953 719 1203 757
rect -1203 -807 -953 -781
rect -895 -807 -645 -781
rect -587 -807 -337 -781
rect -279 -807 -29 -781
rect 29 -807 279 -781
rect 337 -807 587 -781
rect 645 -807 895 -781
rect 953 -807 1203 -781
<< polycont >>
rect -1100 757 -1056 791
rect -792 757 -748 791
rect -484 757 -440 791
rect -176 757 -132 791
rect 132 757 176 791
rect 440 757 484 791
rect 748 757 792 791
rect 1056 757 1100 791
<< locali >>
rect -1116 757 -1100 791
rect -1056 757 -1040 791
rect -808 757 -792 791
rect -748 757 -732 791
rect -500 757 -484 791
rect -440 757 -424 791
rect -192 757 -176 791
rect -132 757 -116 791
rect 116 757 132 791
rect 176 757 192 791
rect 424 757 440 791
rect 484 757 500 791
rect 732 757 748 791
rect 792 757 808 791
rect 1040 757 1056 791
rect 1100 757 1116 791
rect -1249 707 -1215 723
rect -1249 -785 -1215 -769
rect -941 707 -907 723
rect -941 -785 -907 -769
rect -633 707 -599 723
rect -633 -785 -599 -769
rect -325 707 -291 723
rect -325 -785 -291 -769
rect -17 707 17 723
rect -17 -785 17 -769
rect 291 707 325 723
rect 291 -785 325 -769
rect 599 707 633 723
rect 599 -785 633 -769
rect 907 707 941 723
rect 907 -785 941 -769
rect 1215 707 1249 723
rect 1215 -785 1249 -769
<< viali >>
rect -1100 757 -1056 791
rect -792 757 -748 791
rect -484 757 -440 791
rect -176 757 -132 791
rect 132 757 176 791
rect 440 757 484 791
rect 748 757 792 791
rect 1056 757 1100 791
rect -1249 -769 -1215 707
rect -941 -769 -907 707
rect -633 -769 -599 707
rect -325 -769 -291 707
rect -17 -769 17 707
rect 291 -769 325 707
rect 599 -769 633 707
rect 907 -769 941 707
rect 1215 -769 1249 707
<< metal1 >>
rect -1112 791 -1044 797
rect -1112 757 -1100 791
rect -1056 757 -1044 791
rect -1112 751 -1044 757
rect -804 791 -736 797
rect -804 757 -792 791
rect -748 757 -736 791
rect -804 751 -736 757
rect -496 791 -428 797
rect -496 757 -484 791
rect -440 757 -428 791
rect -496 751 -428 757
rect -188 791 -120 797
rect -188 757 -176 791
rect -132 757 -120 791
rect -188 751 -120 757
rect 120 791 188 797
rect 120 757 132 791
rect 176 757 188 791
rect 120 751 188 757
rect 428 791 496 797
rect 428 757 440 791
rect 484 757 496 791
rect 428 751 496 757
rect 736 791 804 797
rect 736 757 748 791
rect 792 757 804 791
rect 736 751 804 757
rect 1044 791 1112 797
rect 1044 757 1056 791
rect 1100 757 1112 791
rect 1044 751 1112 757
rect -1255 707 -1209 719
rect -1255 -769 -1249 707
rect -1215 -769 -1209 707
rect -1255 -781 -1209 -769
rect -947 707 -901 719
rect -947 -769 -941 707
rect -907 -769 -901 707
rect -947 -781 -901 -769
rect -639 707 -593 719
rect -639 -769 -633 707
rect -599 -769 -593 707
rect -639 -781 -593 -769
rect -331 707 -285 719
rect -331 -769 -325 707
rect -291 -769 -285 707
rect -331 -781 -285 -769
rect -23 707 23 719
rect -23 -769 -17 707
rect 17 -769 23 707
rect -23 -781 23 -769
rect 285 707 331 719
rect 285 -769 291 707
rect 325 -769 331 707
rect 285 -781 331 -769
rect 593 707 639 719
rect 593 -769 599 707
rect 633 -769 639 707
rect 593 -781 639 -769
rect 901 707 947 719
rect 901 -769 907 707
rect 941 -769 947 707
rect 901 -781 947 -769
rect 1209 707 1255 719
rect 1209 -769 1215 707
rect 1249 -769 1255 707
rect 1209 -781 1255 -769
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 8 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
