magic
tech sky130A
magscale 1 2
timestamp 1769436194
<< pwell >>
rect -3448 -1932 3448 1932
<< psubdiff >>
rect -3412 1862 -3316 1896
rect 3316 1862 3412 1896
rect -3412 1800 -3378 1862
rect 3378 1800 3412 1862
rect -3412 -1862 -3378 -1800
rect 3378 -1862 3412 -1800
rect -3412 -1896 -3316 -1862
rect 3316 -1896 3412 -1862
<< psubdiffcont >>
rect -3316 1862 3316 1896
rect -3412 -1800 -3378 1800
rect 3378 -1800 3412 1800
rect -3316 -1896 3316 -1862
<< xpolycontact >>
rect -3282 1334 -2712 1766
rect -3282 -1766 -2712 -1334
rect -2616 1334 -2046 1766
rect -2616 -1766 -2046 -1334
rect -1950 1334 -1380 1766
rect -1950 -1766 -1380 -1334
rect -1284 1334 -714 1766
rect -1284 -1766 -714 -1334
rect -618 1334 -48 1766
rect -618 -1766 -48 -1334
rect 48 1334 618 1766
rect 48 -1766 618 -1334
rect 714 1334 1284 1766
rect 714 -1766 1284 -1334
rect 1380 1334 1950 1766
rect 1380 -1766 1950 -1334
rect 2046 1334 2616 1766
rect 2046 -1766 2616 -1334
rect 2712 1334 3282 1766
rect 2712 -1766 3282 -1334
<< ppolyres >>
rect -3282 -1334 -2712 1334
rect -2616 -1334 -2046 1334
rect -1950 -1334 -1380 1334
rect -1284 -1334 -714 1334
rect -618 -1334 -48 1334
rect 48 -1334 618 1334
rect 714 -1334 1284 1334
rect 1380 -1334 1950 1334
rect 2046 -1334 2616 1334
rect 2712 -1334 3282 1334
<< locali >>
rect -3412 1862 -3316 1896
rect 3316 1862 3412 1896
rect -3412 1800 -3378 1862
rect 3378 1800 3412 1862
rect -3412 -1862 -3378 -1800
rect 3378 -1862 3412 -1800
rect -3412 -1896 -3316 -1862
rect 3316 -1896 3412 -1862
<< viali >>
rect -3266 1351 -2728 1748
rect -2600 1351 -2062 1748
rect -1934 1351 -1396 1748
rect -1268 1351 -730 1748
rect -602 1351 -64 1748
rect 64 1351 602 1748
rect 730 1351 1268 1748
rect 1396 1351 1934 1748
rect 2062 1351 2600 1748
rect 2728 1351 3266 1748
rect -3266 -1748 -2728 -1351
rect -2600 -1748 -2062 -1351
rect -1934 -1748 -1396 -1351
rect -1268 -1748 -730 -1351
rect -602 -1748 -64 -1351
rect 64 -1748 602 -1351
rect 730 -1748 1268 -1351
rect 1396 -1748 1934 -1351
rect 2062 -1748 2600 -1351
rect 2728 -1748 3266 -1351
<< metal1 >>
rect -3278 1748 -2716 1754
rect -3278 1351 -3266 1748
rect -2728 1351 -2716 1748
rect -3278 1345 -2716 1351
rect -2612 1748 -2050 1754
rect -2612 1351 -2600 1748
rect -2062 1351 -2050 1748
rect -2612 1345 -2050 1351
rect -1946 1748 -1384 1754
rect -1946 1351 -1934 1748
rect -1396 1351 -1384 1748
rect -1946 1345 -1384 1351
rect -1280 1748 -718 1754
rect -1280 1351 -1268 1748
rect -730 1351 -718 1748
rect -1280 1345 -718 1351
rect -614 1748 -52 1754
rect -614 1351 -602 1748
rect -64 1351 -52 1748
rect -614 1345 -52 1351
rect 52 1748 614 1754
rect 52 1351 64 1748
rect 602 1351 614 1748
rect 52 1345 614 1351
rect 718 1748 1280 1754
rect 718 1351 730 1748
rect 1268 1351 1280 1748
rect 718 1345 1280 1351
rect 1384 1748 1946 1754
rect 1384 1351 1396 1748
rect 1934 1351 1946 1748
rect 1384 1345 1946 1351
rect 2050 1748 2612 1754
rect 2050 1351 2062 1748
rect 2600 1351 2612 1748
rect 2050 1345 2612 1351
rect 2716 1748 3278 1754
rect 2716 1351 2728 1748
rect 3266 1351 3278 1748
rect 2716 1345 3278 1351
rect -3278 -1351 -2716 -1345
rect -3278 -1748 -3266 -1351
rect -2728 -1748 -2716 -1351
rect -3278 -1754 -2716 -1748
rect -2612 -1351 -2050 -1345
rect -2612 -1748 -2600 -1351
rect -2062 -1748 -2050 -1351
rect -2612 -1754 -2050 -1748
rect -1946 -1351 -1384 -1345
rect -1946 -1748 -1934 -1351
rect -1396 -1748 -1384 -1351
rect -1946 -1754 -1384 -1748
rect -1280 -1351 -718 -1345
rect -1280 -1748 -1268 -1351
rect -730 -1748 -718 -1351
rect -1280 -1754 -718 -1748
rect -614 -1351 -52 -1345
rect -614 -1748 -602 -1351
rect -64 -1748 -52 -1351
rect -614 -1754 -52 -1748
rect 52 -1351 614 -1345
rect 52 -1748 64 -1351
rect 602 -1748 614 -1351
rect 52 -1754 614 -1748
rect 718 -1351 1280 -1345
rect 718 -1748 730 -1351
rect 1268 -1748 1280 -1351
rect 718 -1754 1280 -1748
rect 1384 -1351 1946 -1345
rect 1384 -1748 1396 -1351
rect 1934 -1748 1946 -1351
rect 1384 -1754 1946 -1748
rect 2050 -1351 2612 -1345
rect 2050 -1748 2062 -1351
rect 2600 -1748 2612 -1351
rect 2050 -1754 2612 -1748
rect 2716 -1351 3278 -1345
rect 2716 -1748 2728 -1351
rect 3266 -1748 3278 -1351
rect 2716 -1754 3278 -1748
<< properties >>
string FIXED_BBOX -3395 -1879 3395 1879
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string parameters w 2.850 l 13.5 m 1 nx 10 wmin 2.850 lmin 0.50 class resistor rho 319.8 val 1.651k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 2.850 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
