magic
tech sky130A
magscale 1 2
timestamp 1770123317
<< pwell >>
rect -825 -527 825 527
<< mvnmos >>
rect -595 -331 -445 269
rect -387 -331 -237 269
rect -179 -331 -29 269
rect 29 -331 179 269
rect 237 -331 387 269
rect 445 -331 595 269
<< mvndiff >>
rect -653 257 -595 269
rect -653 -319 -641 257
rect -607 -319 -595 257
rect -653 -331 -595 -319
rect -445 257 -387 269
rect -445 -319 -433 257
rect -399 -319 -387 257
rect -445 -331 -387 -319
rect -237 257 -179 269
rect -237 -319 -225 257
rect -191 -319 -179 257
rect -237 -331 -179 -319
rect -29 257 29 269
rect -29 -319 -17 257
rect 17 -319 29 257
rect -29 -331 29 -319
rect 179 257 237 269
rect 179 -319 191 257
rect 225 -319 237 257
rect 179 -331 237 -319
rect 387 257 445 269
rect 387 -319 399 257
rect 433 -319 445 257
rect 387 -331 445 -319
rect 595 257 653 269
rect 595 -319 607 257
rect 641 -319 653 257
rect 595 -331 653 -319
<< mvndiffc >>
rect -641 -319 -607 257
rect -433 -319 -399 257
rect -225 -319 -191 257
rect -17 -319 17 257
rect 191 -319 225 257
rect 399 -319 433 257
rect 607 -319 641 257
<< mvpsubdiff >>
rect -789 433 789 491
rect -789 383 -731 433
rect -789 -383 -777 383
rect -743 -383 -731 383
rect 731 383 789 433
rect -789 -433 -731 -383
rect 731 -383 743 383
rect 777 -383 789 383
rect 731 -433 789 -383
rect -789 -445 789 -433
rect -789 -479 -681 -445
rect 681 -479 789 -445
rect -789 -491 789 -479
<< mvpsubdiffcont >>
rect -777 -383 -743 383
rect 743 -383 777 383
rect -681 -479 681 -445
<< poly >>
rect -595 341 -445 357
rect -595 307 -579 341
rect -461 307 -445 341
rect -595 269 -445 307
rect -387 341 -237 357
rect -387 307 -371 341
rect -253 307 -237 341
rect -387 269 -237 307
rect -179 341 -29 357
rect -179 307 -163 341
rect -45 307 -29 341
rect -179 269 -29 307
rect 29 341 179 357
rect 29 307 45 341
rect 163 307 179 341
rect 29 269 179 307
rect 237 341 387 357
rect 237 307 253 341
rect 371 307 387 341
rect 237 269 387 307
rect 445 341 595 357
rect 445 307 461 341
rect 579 307 595 341
rect 445 269 595 307
rect -595 -357 -445 -331
rect -387 -357 -237 -331
rect -179 -357 -29 -331
rect 29 -357 179 -331
rect 237 -357 387 -331
rect 445 -357 595 -331
<< polycont >>
rect -579 307 -461 341
rect -371 307 -253 341
rect -163 307 -45 341
rect 45 307 163 341
rect 253 307 371 341
rect 461 307 579 341
<< locali >>
rect -777 445 777 479
rect -777 383 -743 445
rect 743 383 777 445
rect -595 307 -579 341
rect -461 307 -445 341
rect -387 307 -371 341
rect -253 307 -237 341
rect -179 307 -163 341
rect -45 307 -29 341
rect 29 307 45 341
rect 163 307 179 341
rect 237 307 253 341
rect 371 307 387 341
rect 445 307 461 341
rect 579 307 595 341
rect -641 257 -607 273
rect -641 -335 -607 -319
rect -433 257 -399 273
rect -433 -335 -399 -319
rect -225 257 -191 273
rect -225 -335 -191 -319
rect -17 257 17 273
rect -17 -335 17 -319
rect 191 257 225 273
rect 191 -335 225 -319
rect 399 257 433 273
rect 399 -335 433 -319
rect 607 257 641 273
rect 607 -335 641 -319
rect -777 -445 -743 -383
rect 743 -445 777 -383
rect -777 -479 -681 -445
rect 681 -479 777 -445
<< viali >>
rect -579 307 -461 341
rect -371 307 -253 341
rect -163 307 -45 341
rect 45 307 163 341
rect 253 307 371 341
rect 461 307 579 341
rect -641 -319 -607 257
rect -433 -319 -399 257
rect -225 -319 -191 257
rect -17 -319 17 257
rect 191 -319 225 257
rect 399 -319 433 257
rect 607 -319 641 257
<< metal1 >>
rect -591 341 -449 347
rect -591 307 -579 341
rect -461 307 -449 341
rect -591 301 -449 307
rect -383 341 -241 347
rect -383 307 -371 341
rect -253 307 -241 341
rect -383 301 -241 307
rect -175 341 -33 347
rect -175 307 -163 341
rect -45 307 -33 341
rect -175 301 -33 307
rect 33 341 175 347
rect 33 307 45 341
rect 163 307 175 341
rect 33 301 175 307
rect 241 341 383 347
rect 241 307 253 341
rect 371 307 383 341
rect 241 301 383 307
rect 449 341 591 347
rect 449 307 461 341
rect 579 307 591 341
rect 449 301 591 307
rect -647 257 -601 269
rect -647 -319 -641 257
rect -607 -319 -601 257
rect -647 -331 -601 -319
rect -439 257 -393 269
rect -439 -319 -433 257
rect -399 -319 -393 257
rect -439 -331 -393 -319
rect -231 257 -185 269
rect -231 -319 -225 257
rect -191 -319 -185 257
rect -231 -331 -185 -319
rect -23 257 23 269
rect -23 -319 -17 257
rect 17 -319 23 257
rect -23 -331 23 -319
rect 185 257 231 269
rect 185 -319 191 257
rect 225 -319 231 257
rect 185 -331 231 -319
rect 393 257 439 269
rect 393 -319 399 257
rect 433 -319 439 257
rect 393 -331 439 -319
rect 601 257 647 269
rect 601 -319 607 257
rect 641 -319 647 257
rect 601 -331 647 -319
<< labels >>
rlabel mvpsubdiffcont 0 -462 0 -462 0 B
port 1 nsew
rlabel mvndiffc -624 -31 -624 -31 0 D0
port 2 nsew
rlabel polycont -520 324 -520 324 0 G0
port 3 nsew
rlabel mvndiffc -416 -31 -416 -31 0 S1
port 4 nsew
rlabel polycont -312 324 -312 324 0 G1
port 5 nsew
rlabel mvndiffc -208 -31 -208 -31 0 D2
port 6 nsew
rlabel polycont -104 324 -104 324 0 G2
port 7 nsew
rlabel mvndiffc 0 -31 0 -31 0 S3
port 8 nsew
rlabel polycont 104 324 104 324 0 G3
port 9 nsew
rlabel mvndiffc 208 -31 208 -31 0 D4
port 10 nsew
rlabel polycont 312 324 312 324 0 G4
port 11 nsew
rlabel mvndiffc 416 -31 416 -31 0 S5
port 12 nsew
rlabel polycont 520 324 520 324 0 G5
port 13 nsew
<< properties >>
string FIXED_BBOX -760 -462 760 462
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 0.75 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
