=============================================================
* tb_ac_pex_mc_final.spice  (PEX-backed, adapted to x1st-stage wrapper)
* =============================================================

.GLOBAL GND

* --- Models / Corner ---
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice mc

* --- Include extracted PEX netlist ---
* Must contain: .subckt x1st-stage VP VN IBIAS VSS OUT VDD
.include "1st-stage_pex.spice"

* =============================================================
* WRAPPER (KEEP YOUR SCHEM SYMBOL PIN ORDER)
* Schematic:  .subckt 1st-stage VDD OUT VN VP IBIAS VSS
* PEX cell:   .subckt x1st-stage VP VN IBIAS VSS OUT VDD
* =============================================================
.subckt 1st-stage VDD OUT VN VP IBIAS VSS
XPEX VP VN IBIAS VSS OUT VDD x1st-stage
.ends 1st-stage


* =============================================================
* TOP-LEVEL TESTBENCH (KEEP EXACT SETUP KAMU)
* =============================================================

* Differential inputs
V2 VN   VSS  AC -1m  DC 1.25
V3 VP   VSS  AC  1m  DC 1.25

* Supplies
V5 VDD  VSS  5
V7 VSS  GND  0

* Bias
I4 VDD  IBIAS 200u

* Output load
C2 OUT  VSS  1p

* Common-mode / CMRR path
V1 VCM  VSS  AC 1m  DC 1.25
C1 OUT2 VSS  5p

* PSRR path: inject AC on VDDr supply feeding x3
V4 VDDr VSS  DC 5  AC 1
C3 OUT3 VSS  10p
R1 OUT3 VN   1k

* DUT instances (WRAPPER subckt)
* Wrapper pin order matches your original schematic:
* .subckt 1st-stage VDD OUT VN VP IBIAS VSS
x1 VDDr OUT3 VN VP IBIAS VSS 1st-stage
x2 VDD  OUT2 VCM VCM IBIAS VSS 1st-stage
x3 VDD  OUT  VN  VP  IBIAS VSS 1st-stage


.control
  set noaskquit
  set temp = 27
  set filetype=ascii
  set appendwrite

  let mc_runs = 300
  let run = 0

  * init vectors (300 entries) — brute force
  compose a0_gain_vec values \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0

  compose pm_val_vec values \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0

  compose cmrr_val_vec values \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0

  compose psrr_val_vec values \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 \
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0

  dowhile run < mc_runs
    reset
    set temp = 27
    setseed (run+1)

    op

    * --- Gain/PM (differential) ---
    alter v1 acmag = 0
    alter v4 acmag = 0

    alter v2 acmag = 1m
    alter v3 acmag = 1m
    alter v2 acphase = 180
    alter v3 acphase = 0

    ac dec 100 1 100meg

    let g_inst = db( v(out) / (v(vp)-v(vn)) )
    let a0_gain_vec[run] = g_inst[0]

    let p_inst = (180/pi) * cph( v(out) / (v(vp)-v(vn)) )
    meas ac p_unity find p_inst when g_inst = 0
    let pm_val_vec[run] = 180 + p_unity

    * --- CMRR (common-mode) ---
    alter v2 acmag = 0
    alter v3 acmag = 0
    alter v1 acmag = 1m
    alter v4 acmag = 0

    ac dec 100 1 100meg
    let a_cm = db( v(out2) / v(vcm) )
    let cmrr_val_vec[run] = a0_gain_vec[run] - a_cm[0]

    * --- PSRR (supply injection) ---
    alter v1 acmag = 0
    alter v2 acmag = 0
    alter v3 acmag = 0
    alter v4 acmag = 1

    ac dec 100 1 100meg
    let psrr_inst = -db( v(out3) )
    let psrr_val_vec[run] = psrr_inst[0]

    echo "MC RUN " run " DONE | A0=" a0_gain_vec[run] " PM=" pm_val_vec[run] " CMRR=" cmrr_val_vec[run] " PSRR=" psrr_val_vec[run]
    let run = run + 1
  end

  echo "---------------- FINAL STATISTICAL REPORT (PEX) ----------------"
  print mean(a0_gain_vec) mean(pm_val_vec) mean(cmrr_val_vec) mean(psrr_val_vec)

  * =============================================================
  * RE-FIXED CSV OUTPUT BLOCK (INDEX EVALUATION)
  * =============================================================
  shell rm -f mc_results.csv
  shell echo "run,A0_dB,PM_deg,CMRR_dB,PSRR_dB" > mc_results.csv

  let i = 0
  dowhile i < mc_runs
    * Pull values into temp scalars so echo can find them easily
    let tmp_a0   = a0_gain_vec[i]
    let tmp_pm   = pm_val_vec[i]
    let tmp_cmrr = cmrr_val_vec[i]
    let tmp_psrr = psrr_val_vec[i]

    * Now echo the scalars
    echo "$&i, $&tmp_a0, $&tmp_pm, $&tmp_cmrr, $&tmp_psrr" >> mc_results.csv

    let i = i + 1
  end

  echo "CSV WRITTEN: mc_results.csv"
.endc
