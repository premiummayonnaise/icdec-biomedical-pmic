magic
tech sky130A
magscale 1 2
timestamp 1768990256
<< mvnmos >>
rect -5047 -781 -4797 719
rect -4619 -781 -4369 719
rect -4191 -781 -3941 719
rect -3763 -781 -3513 719
rect -3335 -781 -3085 719
rect -2907 -781 -2657 719
rect -2479 -781 -2229 719
rect -2051 -781 -1801 719
rect -1623 -781 -1373 719
rect -1195 -781 -945 719
rect -767 -781 -517 719
rect -339 -781 -89 719
rect 89 -781 339 719
rect 517 -781 767 719
rect 945 -781 1195 719
rect 1373 -781 1623 719
rect 1801 -781 2051 719
rect 2229 -781 2479 719
rect 2657 -781 2907 719
rect 3085 -781 3335 719
rect 3513 -781 3763 719
rect 3941 -781 4191 719
rect 4369 -781 4619 719
rect 4797 -781 5047 719
<< mvndiff >>
rect -5105 707 -5047 719
rect -5105 -769 -5093 707
rect -5059 -769 -5047 707
rect -5105 -781 -5047 -769
rect -4797 707 -4739 719
rect -4797 -769 -4785 707
rect -4751 -769 -4739 707
rect -4797 -781 -4739 -769
rect -4677 707 -4619 719
rect -4677 -769 -4665 707
rect -4631 -769 -4619 707
rect -4677 -781 -4619 -769
rect -4369 707 -4311 719
rect -4369 -769 -4357 707
rect -4323 -769 -4311 707
rect -4369 -781 -4311 -769
rect -4249 707 -4191 719
rect -4249 -769 -4237 707
rect -4203 -769 -4191 707
rect -4249 -781 -4191 -769
rect -3941 707 -3883 719
rect -3941 -769 -3929 707
rect -3895 -769 -3883 707
rect -3941 -781 -3883 -769
rect -3821 707 -3763 719
rect -3821 -769 -3809 707
rect -3775 -769 -3763 707
rect -3821 -781 -3763 -769
rect -3513 707 -3455 719
rect -3513 -769 -3501 707
rect -3467 -769 -3455 707
rect -3513 -781 -3455 -769
rect -3393 707 -3335 719
rect -3393 -769 -3381 707
rect -3347 -769 -3335 707
rect -3393 -781 -3335 -769
rect -3085 707 -3027 719
rect -3085 -769 -3073 707
rect -3039 -769 -3027 707
rect -3085 -781 -3027 -769
rect -2965 707 -2907 719
rect -2965 -769 -2953 707
rect -2919 -769 -2907 707
rect -2965 -781 -2907 -769
rect -2657 707 -2599 719
rect -2657 -769 -2645 707
rect -2611 -769 -2599 707
rect -2657 -781 -2599 -769
rect -2537 707 -2479 719
rect -2537 -769 -2525 707
rect -2491 -769 -2479 707
rect -2537 -781 -2479 -769
rect -2229 707 -2171 719
rect -2229 -769 -2217 707
rect -2183 -769 -2171 707
rect -2229 -781 -2171 -769
rect -2109 707 -2051 719
rect -2109 -769 -2097 707
rect -2063 -769 -2051 707
rect -2109 -781 -2051 -769
rect -1801 707 -1743 719
rect -1801 -769 -1789 707
rect -1755 -769 -1743 707
rect -1801 -781 -1743 -769
rect -1681 707 -1623 719
rect -1681 -769 -1669 707
rect -1635 -769 -1623 707
rect -1681 -781 -1623 -769
rect -1373 707 -1315 719
rect -1373 -769 -1361 707
rect -1327 -769 -1315 707
rect -1373 -781 -1315 -769
rect -1253 707 -1195 719
rect -1253 -769 -1241 707
rect -1207 -769 -1195 707
rect -1253 -781 -1195 -769
rect -945 707 -887 719
rect -945 -769 -933 707
rect -899 -769 -887 707
rect -945 -781 -887 -769
rect -825 707 -767 719
rect -825 -769 -813 707
rect -779 -769 -767 707
rect -825 -781 -767 -769
rect -517 707 -459 719
rect -517 -769 -505 707
rect -471 -769 -459 707
rect -517 -781 -459 -769
rect -397 707 -339 719
rect -397 -769 -385 707
rect -351 -769 -339 707
rect -397 -781 -339 -769
rect -89 707 -31 719
rect -89 -769 -77 707
rect -43 -769 -31 707
rect -89 -781 -31 -769
rect 31 707 89 719
rect 31 -769 43 707
rect 77 -769 89 707
rect 31 -781 89 -769
rect 339 707 397 719
rect 339 -769 351 707
rect 385 -769 397 707
rect 339 -781 397 -769
rect 459 707 517 719
rect 459 -769 471 707
rect 505 -769 517 707
rect 459 -781 517 -769
rect 767 707 825 719
rect 767 -769 779 707
rect 813 -769 825 707
rect 767 -781 825 -769
rect 887 707 945 719
rect 887 -769 899 707
rect 933 -769 945 707
rect 887 -781 945 -769
rect 1195 707 1253 719
rect 1195 -769 1207 707
rect 1241 -769 1253 707
rect 1195 -781 1253 -769
rect 1315 707 1373 719
rect 1315 -769 1327 707
rect 1361 -769 1373 707
rect 1315 -781 1373 -769
rect 1623 707 1681 719
rect 1623 -769 1635 707
rect 1669 -769 1681 707
rect 1623 -781 1681 -769
rect 1743 707 1801 719
rect 1743 -769 1755 707
rect 1789 -769 1801 707
rect 1743 -781 1801 -769
rect 2051 707 2109 719
rect 2051 -769 2063 707
rect 2097 -769 2109 707
rect 2051 -781 2109 -769
rect 2171 707 2229 719
rect 2171 -769 2183 707
rect 2217 -769 2229 707
rect 2171 -781 2229 -769
rect 2479 707 2537 719
rect 2479 -769 2491 707
rect 2525 -769 2537 707
rect 2479 -781 2537 -769
rect 2599 707 2657 719
rect 2599 -769 2611 707
rect 2645 -769 2657 707
rect 2599 -781 2657 -769
rect 2907 707 2965 719
rect 2907 -769 2919 707
rect 2953 -769 2965 707
rect 2907 -781 2965 -769
rect 3027 707 3085 719
rect 3027 -769 3039 707
rect 3073 -769 3085 707
rect 3027 -781 3085 -769
rect 3335 707 3393 719
rect 3335 -769 3347 707
rect 3381 -769 3393 707
rect 3335 -781 3393 -769
rect 3455 707 3513 719
rect 3455 -769 3467 707
rect 3501 -769 3513 707
rect 3455 -781 3513 -769
rect 3763 707 3821 719
rect 3763 -769 3775 707
rect 3809 -769 3821 707
rect 3763 -781 3821 -769
rect 3883 707 3941 719
rect 3883 -769 3895 707
rect 3929 -769 3941 707
rect 3883 -781 3941 -769
rect 4191 707 4249 719
rect 4191 -769 4203 707
rect 4237 -769 4249 707
rect 4191 -781 4249 -769
rect 4311 707 4369 719
rect 4311 -769 4323 707
rect 4357 -769 4369 707
rect 4311 -781 4369 -769
rect 4619 707 4677 719
rect 4619 -769 4631 707
rect 4665 -769 4677 707
rect 4619 -781 4677 -769
rect 4739 707 4797 719
rect 4739 -769 4751 707
rect 4785 -769 4797 707
rect 4739 -781 4797 -769
rect 5047 707 5105 719
rect 5047 -769 5059 707
rect 5093 -769 5105 707
rect 5047 -781 5105 -769
<< mvndiffc >>
rect -5093 -769 -5059 707
rect -4785 -769 -4751 707
rect -4665 -769 -4631 707
rect -4357 -769 -4323 707
rect -4237 -769 -4203 707
rect -3929 -769 -3895 707
rect -3809 -769 -3775 707
rect -3501 -769 -3467 707
rect -3381 -769 -3347 707
rect -3073 -769 -3039 707
rect -2953 -769 -2919 707
rect -2645 -769 -2611 707
rect -2525 -769 -2491 707
rect -2217 -769 -2183 707
rect -2097 -769 -2063 707
rect -1789 -769 -1755 707
rect -1669 -769 -1635 707
rect -1361 -769 -1327 707
rect -1241 -769 -1207 707
rect -933 -769 -899 707
rect -813 -769 -779 707
rect -505 -769 -471 707
rect -385 -769 -351 707
rect -77 -769 -43 707
rect 43 -769 77 707
rect 351 -769 385 707
rect 471 -769 505 707
rect 779 -769 813 707
rect 899 -769 933 707
rect 1207 -769 1241 707
rect 1327 -769 1361 707
rect 1635 -769 1669 707
rect 1755 -769 1789 707
rect 2063 -769 2097 707
rect 2183 -769 2217 707
rect 2491 -769 2525 707
rect 2611 -769 2645 707
rect 2919 -769 2953 707
rect 3039 -769 3073 707
rect 3347 -769 3381 707
rect 3467 -769 3501 707
rect 3775 -769 3809 707
rect 3895 -769 3929 707
rect 4203 -769 4237 707
rect 4323 -769 4357 707
rect 4631 -769 4665 707
rect 4751 -769 4785 707
rect 5059 -769 5093 707
<< poly >>
rect -5047 791 -4797 807
rect -5047 757 -5031 791
rect -4813 757 -4797 791
rect -5047 719 -4797 757
rect -4619 791 -4369 807
rect -4619 757 -4603 791
rect -4385 757 -4369 791
rect -4619 719 -4369 757
rect -4191 791 -3941 807
rect -4191 757 -4175 791
rect -3957 757 -3941 791
rect -4191 719 -3941 757
rect -3763 791 -3513 807
rect -3763 757 -3747 791
rect -3529 757 -3513 791
rect -3763 719 -3513 757
rect -3335 791 -3085 807
rect -3335 757 -3319 791
rect -3101 757 -3085 791
rect -3335 719 -3085 757
rect -2907 791 -2657 807
rect -2907 757 -2891 791
rect -2673 757 -2657 791
rect -2907 719 -2657 757
rect -2479 791 -2229 807
rect -2479 757 -2463 791
rect -2245 757 -2229 791
rect -2479 719 -2229 757
rect -2051 791 -1801 807
rect -2051 757 -2035 791
rect -1817 757 -1801 791
rect -2051 719 -1801 757
rect -1623 791 -1373 807
rect -1623 757 -1607 791
rect -1389 757 -1373 791
rect -1623 719 -1373 757
rect -1195 791 -945 807
rect -1195 757 -1179 791
rect -961 757 -945 791
rect -1195 719 -945 757
rect -767 791 -517 807
rect -767 757 -751 791
rect -533 757 -517 791
rect -767 719 -517 757
rect -339 791 -89 807
rect -339 757 -323 791
rect -105 757 -89 791
rect -339 719 -89 757
rect 89 791 339 807
rect 89 757 105 791
rect 323 757 339 791
rect 89 719 339 757
rect 517 791 767 807
rect 517 757 533 791
rect 751 757 767 791
rect 517 719 767 757
rect 945 791 1195 807
rect 945 757 961 791
rect 1179 757 1195 791
rect 945 719 1195 757
rect 1373 791 1623 807
rect 1373 757 1389 791
rect 1607 757 1623 791
rect 1373 719 1623 757
rect 1801 791 2051 807
rect 1801 757 1817 791
rect 2035 757 2051 791
rect 1801 719 2051 757
rect 2229 791 2479 807
rect 2229 757 2245 791
rect 2463 757 2479 791
rect 2229 719 2479 757
rect 2657 791 2907 807
rect 2657 757 2673 791
rect 2891 757 2907 791
rect 2657 719 2907 757
rect 3085 791 3335 807
rect 3085 757 3101 791
rect 3319 757 3335 791
rect 3085 719 3335 757
rect 3513 791 3763 807
rect 3513 757 3529 791
rect 3747 757 3763 791
rect 3513 719 3763 757
rect 3941 791 4191 807
rect 3941 757 3957 791
rect 4175 757 4191 791
rect 3941 719 4191 757
rect 4369 791 4619 807
rect 4369 757 4385 791
rect 4603 757 4619 791
rect 4369 719 4619 757
rect 4797 791 5047 807
rect 4797 757 4813 791
rect 5031 757 5047 791
rect 4797 719 5047 757
rect -5047 -807 -4797 -781
rect -4619 -807 -4369 -781
rect -4191 -807 -3941 -781
rect -3763 -807 -3513 -781
rect -3335 -807 -3085 -781
rect -2907 -807 -2657 -781
rect -2479 -807 -2229 -781
rect -2051 -807 -1801 -781
rect -1623 -807 -1373 -781
rect -1195 -807 -945 -781
rect -767 -807 -517 -781
rect -339 -807 -89 -781
rect 89 -807 339 -781
rect 517 -807 767 -781
rect 945 -807 1195 -781
rect 1373 -807 1623 -781
rect 1801 -807 2051 -781
rect 2229 -807 2479 -781
rect 2657 -807 2907 -781
rect 3085 -807 3335 -781
rect 3513 -807 3763 -781
rect 3941 -807 4191 -781
rect 4369 -807 4619 -781
rect 4797 -807 5047 -781
<< polycont >>
rect -5031 757 -4813 791
rect -4603 757 -4385 791
rect -4175 757 -3957 791
rect -3747 757 -3529 791
rect -3319 757 -3101 791
rect -2891 757 -2673 791
rect -2463 757 -2245 791
rect -2035 757 -1817 791
rect -1607 757 -1389 791
rect -1179 757 -961 791
rect -751 757 -533 791
rect -323 757 -105 791
rect 105 757 323 791
rect 533 757 751 791
rect 961 757 1179 791
rect 1389 757 1607 791
rect 1817 757 2035 791
rect 2245 757 2463 791
rect 2673 757 2891 791
rect 3101 757 3319 791
rect 3529 757 3747 791
rect 3957 757 4175 791
rect 4385 757 4603 791
rect 4813 757 5031 791
<< locali >>
rect -5047 757 -5031 791
rect -4813 757 -4797 791
rect -4619 757 -4603 791
rect -4385 757 -4369 791
rect -4191 757 -4175 791
rect -3957 757 -3941 791
rect -3763 757 -3747 791
rect -3529 757 -3513 791
rect -3335 757 -3319 791
rect -3101 757 -3085 791
rect -2907 757 -2891 791
rect -2673 757 -2657 791
rect -2479 757 -2463 791
rect -2245 757 -2229 791
rect -2051 757 -2035 791
rect -1817 757 -1801 791
rect -1623 757 -1607 791
rect -1389 757 -1373 791
rect -1195 757 -1179 791
rect -961 757 -945 791
rect -767 757 -751 791
rect -533 757 -517 791
rect -339 757 -323 791
rect -105 757 -89 791
rect 89 757 105 791
rect 323 757 339 791
rect 517 757 533 791
rect 751 757 767 791
rect 945 757 961 791
rect 1179 757 1195 791
rect 1373 757 1389 791
rect 1607 757 1623 791
rect 1801 757 1817 791
rect 2035 757 2051 791
rect 2229 757 2245 791
rect 2463 757 2479 791
rect 2657 757 2673 791
rect 2891 757 2907 791
rect 3085 757 3101 791
rect 3319 757 3335 791
rect 3513 757 3529 791
rect 3747 757 3763 791
rect 3941 757 3957 791
rect 4175 757 4191 791
rect 4369 757 4385 791
rect 4603 757 4619 791
rect 4797 757 4813 791
rect 5031 757 5047 791
rect -5093 707 -5059 723
rect -5093 -785 -5059 -769
rect -4785 707 -4751 723
rect -4785 -785 -4751 -769
rect -4665 707 -4631 723
rect -4665 -785 -4631 -769
rect -4357 707 -4323 723
rect -4357 -785 -4323 -769
rect -4237 707 -4203 723
rect -4237 -785 -4203 -769
rect -3929 707 -3895 723
rect -3929 -785 -3895 -769
rect -3809 707 -3775 723
rect -3809 -785 -3775 -769
rect -3501 707 -3467 723
rect -3501 -785 -3467 -769
rect -3381 707 -3347 723
rect -3381 -785 -3347 -769
rect -3073 707 -3039 723
rect -3073 -785 -3039 -769
rect -2953 707 -2919 723
rect -2953 -785 -2919 -769
rect -2645 707 -2611 723
rect -2645 -785 -2611 -769
rect -2525 707 -2491 723
rect -2525 -785 -2491 -769
rect -2217 707 -2183 723
rect -2217 -785 -2183 -769
rect -2097 707 -2063 723
rect -2097 -785 -2063 -769
rect -1789 707 -1755 723
rect -1789 -785 -1755 -769
rect -1669 707 -1635 723
rect -1669 -785 -1635 -769
rect -1361 707 -1327 723
rect -1361 -785 -1327 -769
rect -1241 707 -1207 723
rect -1241 -785 -1207 -769
rect -933 707 -899 723
rect -933 -785 -899 -769
rect -813 707 -779 723
rect -813 -785 -779 -769
rect -505 707 -471 723
rect -505 -785 -471 -769
rect -385 707 -351 723
rect -385 -785 -351 -769
rect -77 707 -43 723
rect -77 -785 -43 -769
rect 43 707 77 723
rect 43 -785 77 -769
rect 351 707 385 723
rect 351 -785 385 -769
rect 471 707 505 723
rect 471 -785 505 -769
rect 779 707 813 723
rect 779 -785 813 -769
rect 899 707 933 723
rect 899 -785 933 -769
rect 1207 707 1241 723
rect 1207 -785 1241 -769
rect 1327 707 1361 723
rect 1327 -785 1361 -769
rect 1635 707 1669 723
rect 1635 -785 1669 -769
rect 1755 707 1789 723
rect 1755 -785 1789 -769
rect 2063 707 2097 723
rect 2063 -785 2097 -769
rect 2183 707 2217 723
rect 2183 -785 2217 -769
rect 2491 707 2525 723
rect 2491 -785 2525 -769
rect 2611 707 2645 723
rect 2611 -785 2645 -769
rect 2919 707 2953 723
rect 2919 -785 2953 -769
rect 3039 707 3073 723
rect 3039 -785 3073 -769
rect 3347 707 3381 723
rect 3347 -785 3381 -769
rect 3467 707 3501 723
rect 3467 -785 3501 -769
rect 3775 707 3809 723
rect 3775 -785 3809 -769
rect 3895 707 3929 723
rect 3895 -785 3929 -769
rect 4203 707 4237 723
rect 4203 -785 4237 -769
rect 4323 707 4357 723
rect 4323 -785 4357 -769
rect 4631 707 4665 723
rect 4631 -785 4665 -769
rect 4751 707 4785 723
rect 4751 -785 4785 -769
rect 5059 707 5093 723
rect 5059 -785 5093 -769
<< viali >>
rect -5031 757 -4813 791
rect -4603 757 -4385 791
rect -4175 757 -3957 791
rect -3747 757 -3529 791
rect -3319 757 -3101 791
rect -2891 757 -2673 791
rect -2463 757 -2245 791
rect -2035 757 -1817 791
rect -1607 757 -1389 791
rect -1179 757 -961 791
rect -751 757 -533 791
rect -323 757 -105 791
rect 105 757 323 791
rect 533 757 751 791
rect 961 757 1179 791
rect 1389 757 1607 791
rect 1817 757 2035 791
rect 2245 757 2463 791
rect 2673 757 2891 791
rect 3101 757 3319 791
rect 3529 757 3747 791
rect 3957 757 4175 791
rect 4385 757 4603 791
rect 4813 757 5031 791
rect -5093 -769 -5059 707
rect -4785 -769 -4751 707
rect -4665 -769 -4631 707
rect -4357 -769 -4323 707
rect -4237 -769 -4203 707
rect -3929 -769 -3895 707
rect -3809 -769 -3775 707
rect -3501 -769 -3467 707
rect -3381 -769 -3347 707
rect -3073 -769 -3039 707
rect -2953 -769 -2919 707
rect -2645 -769 -2611 707
rect -2525 -769 -2491 707
rect -2217 -769 -2183 707
rect -2097 -769 -2063 707
rect -1789 -769 -1755 707
rect -1669 -769 -1635 707
rect -1361 -769 -1327 707
rect -1241 -769 -1207 707
rect -933 -769 -899 707
rect -813 -769 -779 707
rect -505 -769 -471 707
rect -385 -769 -351 707
rect -77 -769 -43 707
rect 43 -769 77 707
rect 351 -769 385 707
rect 471 -769 505 707
rect 779 -769 813 707
rect 899 -769 933 707
rect 1207 -769 1241 707
rect 1327 -769 1361 707
rect 1635 -769 1669 707
rect 1755 -769 1789 707
rect 2063 -769 2097 707
rect 2183 -769 2217 707
rect 2491 -769 2525 707
rect 2611 -769 2645 707
rect 2919 -769 2953 707
rect 3039 -769 3073 707
rect 3347 -769 3381 707
rect 3467 -769 3501 707
rect 3775 -769 3809 707
rect 3895 -769 3929 707
rect 4203 -769 4237 707
rect 4323 -769 4357 707
rect 4631 -769 4665 707
rect 4751 -769 4785 707
rect 5059 -769 5093 707
<< metal1 >>
rect -5043 791 -4801 797
rect -5043 757 -5031 791
rect -4813 757 -4801 791
rect -5043 751 -4801 757
rect -4615 791 -4373 797
rect -4615 757 -4603 791
rect -4385 757 -4373 791
rect -4615 751 -4373 757
rect -4187 791 -3945 797
rect -4187 757 -4175 791
rect -3957 757 -3945 791
rect -4187 751 -3945 757
rect -3759 791 -3517 797
rect -3759 757 -3747 791
rect -3529 757 -3517 791
rect -3759 751 -3517 757
rect -3331 791 -3089 797
rect -3331 757 -3319 791
rect -3101 757 -3089 791
rect -3331 751 -3089 757
rect -2903 791 -2661 797
rect -2903 757 -2891 791
rect -2673 757 -2661 791
rect -2903 751 -2661 757
rect -2475 791 -2233 797
rect -2475 757 -2463 791
rect -2245 757 -2233 791
rect -2475 751 -2233 757
rect -2047 791 -1805 797
rect -2047 757 -2035 791
rect -1817 757 -1805 791
rect -2047 751 -1805 757
rect -1619 791 -1377 797
rect -1619 757 -1607 791
rect -1389 757 -1377 791
rect -1619 751 -1377 757
rect -1191 791 -949 797
rect -1191 757 -1179 791
rect -961 757 -949 791
rect -1191 751 -949 757
rect -763 791 -521 797
rect -763 757 -751 791
rect -533 757 -521 791
rect -763 751 -521 757
rect -335 791 -93 797
rect -335 757 -323 791
rect -105 757 -93 791
rect -335 751 -93 757
rect 93 791 335 797
rect 93 757 105 791
rect 323 757 335 791
rect 93 751 335 757
rect 521 791 763 797
rect 521 757 533 791
rect 751 757 763 791
rect 521 751 763 757
rect 949 791 1191 797
rect 949 757 961 791
rect 1179 757 1191 791
rect 949 751 1191 757
rect 1377 791 1619 797
rect 1377 757 1389 791
rect 1607 757 1619 791
rect 1377 751 1619 757
rect 1805 791 2047 797
rect 1805 757 1817 791
rect 2035 757 2047 791
rect 1805 751 2047 757
rect 2233 791 2475 797
rect 2233 757 2245 791
rect 2463 757 2475 791
rect 2233 751 2475 757
rect 2661 791 2903 797
rect 2661 757 2673 791
rect 2891 757 2903 791
rect 2661 751 2903 757
rect 3089 791 3331 797
rect 3089 757 3101 791
rect 3319 757 3331 791
rect 3089 751 3331 757
rect 3517 791 3759 797
rect 3517 757 3529 791
rect 3747 757 3759 791
rect 3517 751 3759 757
rect 3945 791 4187 797
rect 3945 757 3957 791
rect 4175 757 4187 791
rect 3945 751 4187 757
rect 4373 791 4615 797
rect 4373 757 4385 791
rect 4603 757 4615 791
rect 4373 751 4615 757
rect 4801 791 5043 797
rect 4801 757 4813 791
rect 5031 757 5043 791
rect 4801 751 5043 757
rect -5099 707 -5053 719
rect -5099 -769 -5093 707
rect -5059 -769 -5053 707
rect -5099 -781 -5053 -769
rect -4791 707 -4745 719
rect -4791 -769 -4785 707
rect -4751 -769 -4745 707
rect -4791 -781 -4745 -769
rect -4671 707 -4625 719
rect -4671 -769 -4665 707
rect -4631 -769 -4625 707
rect -4671 -781 -4625 -769
rect -4363 707 -4317 719
rect -4363 -769 -4357 707
rect -4323 -769 -4317 707
rect -4363 -781 -4317 -769
rect -4243 707 -4197 719
rect -4243 -769 -4237 707
rect -4203 -769 -4197 707
rect -4243 -781 -4197 -769
rect -3935 707 -3889 719
rect -3935 -769 -3929 707
rect -3895 -769 -3889 707
rect -3935 -781 -3889 -769
rect -3815 707 -3769 719
rect -3815 -769 -3809 707
rect -3775 -769 -3769 707
rect -3815 -781 -3769 -769
rect -3507 707 -3461 719
rect -3507 -769 -3501 707
rect -3467 -769 -3461 707
rect -3507 -781 -3461 -769
rect -3387 707 -3341 719
rect -3387 -769 -3381 707
rect -3347 -769 -3341 707
rect -3387 -781 -3341 -769
rect -3079 707 -3033 719
rect -3079 -769 -3073 707
rect -3039 -769 -3033 707
rect -3079 -781 -3033 -769
rect -2959 707 -2913 719
rect -2959 -769 -2953 707
rect -2919 -769 -2913 707
rect -2959 -781 -2913 -769
rect -2651 707 -2605 719
rect -2651 -769 -2645 707
rect -2611 -769 -2605 707
rect -2651 -781 -2605 -769
rect -2531 707 -2485 719
rect -2531 -769 -2525 707
rect -2491 -769 -2485 707
rect -2531 -781 -2485 -769
rect -2223 707 -2177 719
rect -2223 -769 -2217 707
rect -2183 -769 -2177 707
rect -2223 -781 -2177 -769
rect -2103 707 -2057 719
rect -2103 -769 -2097 707
rect -2063 -769 -2057 707
rect -2103 -781 -2057 -769
rect -1795 707 -1749 719
rect -1795 -769 -1789 707
rect -1755 -769 -1749 707
rect -1795 -781 -1749 -769
rect -1675 707 -1629 719
rect -1675 -769 -1669 707
rect -1635 -769 -1629 707
rect -1675 -781 -1629 -769
rect -1367 707 -1321 719
rect -1367 -769 -1361 707
rect -1327 -769 -1321 707
rect -1367 -781 -1321 -769
rect -1247 707 -1201 719
rect -1247 -769 -1241 707
rect -1207 -769 -1201 707
rect -1247 -781 -1201 -769
rect -939 707 -893 719
rect -939 -769 -933 707
rect -899 -769 -893 707
rect -939 -781 -893 -769
rect -819 707 -773 719
rect -819 -769 -813 707
rect -779 -769 -773 707
rect -819 -781 -773 -769
rect -511 707 -465 719
rect -511 -769 -505 707
rect -471 -769 -465 707
rect -511 -781 -465 -769
rect -391 707 -345 719
rect -391 -769 -385 707
rect -351 -769 -345 707
rect -391 -781 -345 -769
rect -83 707 -37 719
rect -83 -769 -77 707
rect -43 -769 -37 707
rect -83 -781 -37 -769
rect 37 707 83 719
rect 37 -769 43 707
rect 77 -769 83 707
rect 37 -781 83 -769
rect 345 707 391 719
rect 345 -769 351 707
rect 385 -769 391 707
rect 345 -781 391 -769
rect 465 707 511 719
rect 465 -769 471 707
rect 505 -769 511 707
rect 465 -781 511 -769
rect 773 707 819 719
rect 773 -769 779 707
rect 813 -769 819 707
rect 773 -781 819 -769
rect 893 707 939 719
rect 893 -769 899 707
rect 933 -769 939 707
rect 893 -781 939 -769
rect 1201 707 1247 719
rect 1201 -769 1207 707
rect 1241 -769 1247 707
rect 1201 -781 1247 -769
rect 1321 707 1367 719
rect 1321 -769 1327 707
rect 1361 -769 1367 707
rect 1321 -781 1367 -769
rect 1629 707 1675 719
rect 1629 -769 1635 707
rect 1669 -769 1675 707
rect 1629 -781 1675 -769
rect 1749 707 1795 719
rect 1749 -769 1755 707
rect 1789 -769 1795 707
rect 1749 -781 1795 -769
rect 2057 707 2103 719
rect 2057 -769 2063 707
rect 2097 -769 2103 707
rect 2057 -781 2103 -769
rect 2177 707 2223 719
rect 2177 -769 2183 707
rect 2217 -769 2223 707
rect 2177 -781 2223 -769
rect 2485 707 2531 719
rect 2485 -769 2491 707
rect 2525 -769 2531 707
rect 2485 -781 2531 -769
rect 2605 707 2651 719
rect 2605 -769 2611 707
rect 2645 -769 2651 707
rect 2605 -781 2651 -769
rect 2913 707 2959 719
rect 2913 -769 2919 707
rect 2953 -769 2959 707
rect 2913 -781 2959 -769
rect 3033 707 3079 719
rect 3033 -769 3039 707
rect 3073 -769 3079 707
rect 3033 -781 3079 -769
rect 3341 707 3387 719
rect 3341 -769 3347 707
rect 3381 -769 3387 707
rect 3341 -781 3387 -769
rect 3461 707 3507 719
rect 3461 -769 3467 707
rect 3501 -769 3507 707
rect 3461 -781 3507 -769
rect 3769 707 3815 719
rect 3769 -769 3775 707
rect 3809 -769 3815 707
rect 3769 -781 3815 -769
rect 3889 707 3935 719
rect 3889 -769 3895 707
rect 3929 -769 3935 707
rect 3889 -781 3935 -769
rect 4197 707 4243 719
rect 4197 -769 4203 707
rect 4237 -769 4243 707
rect 4197 -781 4243 -769
rect 4317 707 4363 719
rect 4317 -769 4323 707
rect 4357 -769 4363 707
rect 4317 -781 4363 -769
rect 4625 707 4671 719
rect 4625 -769 4631 707
rect 4665 -769 4671 707
rect 4625 -781 4671 -769
rect 4745 707 4791 719
rect 4745 -769 4751 707
rect 4785 -769 4791 707
rect 4745 -781 4791 -769
rect 5053 707 5099 719
rect 5053 -769 5059 707
rect 5093 -769 5099 707
rect 5053 -781 5099 -769
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 24 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
