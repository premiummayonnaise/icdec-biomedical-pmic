magic
tech sky130A
timestamp 1769135993
<< nmos >>
rect -440 -68 -365 37
rect -279 -68 -204 37
rect -118 -68 -43 37
rect 43 -68 118 37
rect 204 -68 279 37
rect 365 -68 440 37
<< ndiff >>
rect -469 31 -440 37
rect -469 -62 -463 31
rect -446 -62 -440 31
rect -469 -68 -440 -62
rect -365 31 -336 37
rect -365 -62 -359 31
rect -342 -62 -336 31
rect -365 -68 -336 -62
rect -308 31 -279 37
rect -308 -62 -302 31
rect -285 -62 -279 31
rect -308 -68 -279 -62
rect -204 31 -175 37
rect -204 -62 -198 31
rect -181 -62 -175 31
rect -204 -68 -175 -62
rect -147 31 -118 37
rect -147 -62 -141 31
rect -124 -62 -118 31
rect -147 -68 -118 -62
rect -43 31 -14 37
rect -43 -62 -37 31
rect -20 -62 -14 31
rect -43 -68 -14 -62
rect 14 31 43 37
rect 14 -62 20 31
rect 37 -62 43 31
rect 14 -68 43 -62
rect 118 31 147 37
rect 118 -62 124 31
rect 141 -62 147 31
rect 118 -68 147 -62
rect 175 31 204 37
rect 175 -62 181 31
rect 198 -62 204 31
rect 175 -68 204 -62
rect 279 31 308 37
rect 279 -62 285 31
rect 302 -62 308 31
rect 279 -68 308 -62
rect 336 31 365 37
rect 336 -62 342 31
rect 359 -62 365 31
rect 336 -68 365 -62
rect 440 31 469 37
rect 440 -62 446 31
rect 463 -62 469 31
rect 440 -68 469 -62
<< ndiffc >>
rect -463 -62 -446 31
rect -359 -62 -342 31
rect -302 -62 -285 31
rect -198 -62 -181 31
rect -141 -62 -124 31
rect -37 -62 -20 31
rect 20 -62 37 31
rect 124 -62 141 31
rect 181 -62 198 31
rect 285 -62 302 31
rect 342 -62 359 31
rect 446 -62 463 31
<< poly >>
rect -440 73 -365 81
rect -440 56 -432 73
rect -373 56 -365 73
rect -440 37 -365 56
rect -279 73 -204 81
rect -279 56 -271 73
rect -212 56 -204 73
rect -279 37 -204 56
rect -118 73 -43 81
rect -118 56 -110 73
rect -51 56 -43 73
rect -118 37 -43 56
rect 43 73 118 81
rect 43 56 51 73
rect 110 56 118 73
rect 43 37 118 56
rect 204 73 279 81
rect 204 56 212 73
rect 271 56 279 73
rect 204 37 279 56
rect 365 73 440 81
rect 365 56 373 73
rect 432 56 440 73
rect 365 37 440 56
rect -440 -81 -365 -68
rect -279 -81 -204 -68
rect -118 -81 -43 -68
rect 43 -81 118 -68
rect 204 -81 279 -68
rect 365 -81 440 -68
<< polycont >>
rect -432 56 -373 73
rect -271 56 -212 73
rect -110 56 -51 73
rect 51 56 110 73
rect 212 56 271 73
rect 373 56 432 73
<< locali >>
rect -440 56 -432 73
rect -373 56 -365 73
rect -279 56 -271 73
rect -212 56 -204 73
rect -118 56 -110 73
rect -51 56 -43 73
rect 43 56 51 73
rect 110 56 118 73
rect 204 56 212 73
rect 271 56 279 73
rect 365 56 373 73
rect 432 56 440 73
rect -463 31 -446 39
rect -463 -70 -446 -62
rect -359 31 -342 39
rect -359 -70 -342 -62
rect -302 31 -285 39
rect -302 -70 -285 -62
rect -198 31 -181 39
rect -198 -70 -181 -62
rect -141 31 -124 39
rect -141 -70 -124 -62
rect -37 31 -20 39
rect -37 -70 -20 -62
rect 20 31 37 39
rect 20 -70 37 -62
rect 124 31 141 39
rect 124 -70 141 -62
rect 181 31 198 39
rect 181 -70 198 -62
rect 285 31 302 39
rect 285 -70 302 -62
rect 342 31 359 39
rect 342 -70 359 -62
rect 446 31 463 39
rect 446 -70 463 -62
<< viali >>
rect -432 56 -373 73
rect -271 56 -212 73
rect -110 56 -51 73
rect 51 56 110 73
rect 212 56 271 73
rect 373 56 432 73
rect -463 -62 -446 31
rect -359 -62 -342 31
rect -302 -62 -285 31
rect -198 -62 -181 31
rect -141 -62 -124 31
rect -37 -62 -20 31
rect 20 -62 37 31
rect 124 -62 141 31
rect 181 -62 198 31
rect 285 -62 302 31
rect 342 -62 359 31
rect 446 -62 463 31
<< metal1 >>
rect -438 73 -367 76
rect -438 56 -432 73
rect -373 56 -367 73
rect -438 53 -367 56
rect -277 73 -206 76
rect -277 56 -271 73
rect -212 56 -206 73
rect -277 53 -206 56
rect -116 73 -45 76
rect -116 56 -110 73
rect -51 56 -45 73
rect -116 53 -45 56
rect 45 73 116 76
rect 45 56 51 73
rect 110 56 116 73
rect 45 53 116 56
rect 206 73 277 76
rect 206 56 212 73
rect 271 56 277 73
rect 206 53 277 56
rect 367 73 438 76
rect 367 56 373 73
rect 432 56 438 73
rect 367 53 438 56
rect -466 31 -443 37
rect -466 -62 -463 31
rect -446 -62 -443 31
rect -466 -68 -443 -62
rect -362 31 -339 37
rect -362 -62 -359 31
rect -342 -62 -339 31
rect -362 -68 -339 -62
rect -305 31 -282 37
rect -305 -62 -302 31
rect -285 -62 -282 31
rect -305 -68 -282 -62
rect -201 31 -178 37
rect -201 -62 -198 31
rect -181 -62 -178 31
rect -201 -68 -178 -62
rect -144 31 -121 37
rect -144 -62 -141 31
rect -124 -62 -121 31
rect -144 -68 -121 -62
rect -40 31 -17 37
rect -40 -62 -37 31
rect -20 -62 -17 31
rect -40 -68 -17 -62
rect 17 31 40 37
rect 17 -62 20 31
rect 37 -62 40 31
rect 17 -68 40 -62
rect 121 31 144 37
rect 121 -62 124 31
rect 141 -62 144 31
rect 121 -68 144 -62
rect 178 31 201 37
rect 178 -62 181 31
rect 198 -62 201 31
rect 178 -68 201 -62
rect 282 31 305 37
rect 282 -62 285 31
rect 302 -62 305 31
rect 282 -68 305 -62
rect 339 31 362 37
rect 339 -62 342 31
rect 359 -62 362 31
rect 339 -68 362 -62
rect 443 31 466 37
rect 443 -62 446 31
rect 463 -62 466 31
rect 443 -68 466 -62
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.05 l 0.75 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
