magic
tech sky130A
magscale 1 2
timestamp 1769616064
<< nwell >>
rect -845 -540 845 540
<< mvpmos >>
rect -587 -243 -337 243
rect -279 -243 -29 243
rect 29 -243 279 243
rect 337 -243 587 243
<< mvpdiff >>
rect -645 231 -587 243
rect -645 -231 -633 231
rect -599 -231 -587 231
rect -645 -243 -587 -231
rect -337 231 -279 243
rect -337 -231 -325 231
rect -291 -231 -279 231
rect -337 -243 -279 -231
rect -29 231 29 243
rect -29 -231 -17 231
rect 17 -231 29 231
rect -29 -243 29 -231
rect 279 231 337 243
rect 279 -231 291 231
rect 325 -231 337 231
rect 279 -243 337 -231
rect 587 231 645 243
rect 587 -231 599 231
rect 633 -231 645 231
rect 587 -243 645 -231
<< mvpdiffc >>
rect -633 -231 -599 231
rect -325 -231 -291 231
rect -17 -231 17 231
rect 291 -231 325 231
rect 599 -231 633 231
<< mvnsubdiff >>
rect -779 462 779 474
rect -779 428 -671 462
rect 671 428 779 462
rect -779 416 779 428
rect -779 366 -721 416
rect -779 -366 -767 366
rect -733 -366 -721 366
rect 721 366 779 416
rect -779 -416 -721 -366
rect 721 -366 733 366
rect 767 -366 779 366
rect 721 -416 779 -366
rect -779 -428 779 -416
rect -779 -462 -671 -428
rect 671 -462 779 -428
rect -779 -474 779 -462
<< mvnsubdiffcont >>
rect -671 428 671 462
rect -767 -366 -733 366
rect 733 -366 767 366
rect -671 -462 671 -428
<< poly >>
rect -587 324 -337 340
rect -587 290 -571 324
rect -353 290 -337 324
rect -587 243 -337 290
rect -279 324 -29 340
rect -279 290 -263 324
rect -45 290 -29 324
rect -279 243 -29 290
rect 29 324 279 340
rect 29 290 45 324
rect 263 290 279 324
rect 29 243 279 290
rect 337 324 587 340
rect 337 290 353 324
rect 571 290 587 324
rect 337 243 587 290
rect -587 -290 -337 -243
rect -587 -324 -571 -290
rect -353 -324 -337 -290
rect -587 -340 -337 -324
rect -279 -290 -29 -243
rect -279 -324 -263 -290
rect -45 -324 -29 -290
rect -279 -340 -29 -324
rect 29 -290 279 -243
rect 29 -324 45 -290
rect 263 -324 279 -290
rect 29 -340 279 -324
rect 337 -290 587 -243
rect 337 -324 353 -290
rect 571 -324 587 -290
rect 337 -340 587 -324
<< polycont >>
rect -571 290 -353 324
rect -263 290 -45 324
rect 45 290 263 324
rect 353 290 571 324
rect -571 -324 -353 -290
rect -263 -324 -45 -290
rect 45 -324 263 -290
rect 353 -324 571 -290
<< locali >>
rect -767 428 -671 462
rect 671 428 767 462
rect -767 366 -733 428
rect 733 366 767 428
rect -587 290 -571 324
rect -353 290 -337 324
rect -279 290 -263 324
rect -45 290 -29 324
rect 29 290 45 324
rect 263 290 279 324
rect 337 290 353 324
rect 571 290 587 324
rect -633 231 -599 247
rect -633 -247 -599 -231
rect -325 231 -291 247
rect -325 -247 -291 -231
rect -17 231 17 247
rect -17 -247 17 -231
rect 291 231 325 247
rect 291 -247 325 -231
rect 599 231 633 247
rect 599 -247 633 -231
rect -587 -324 -571 -290
rect -353 -324 -337 -290
rect -279 -324 -263 -290
rect -45 -324 -29 -290
rect 29 -324 45 -290
rect 263 -324 279 -290
rect 337 -324 353 -290
rect 571 -324 587 -290
rect -767 -428 -733 -366
rect 733 -428 767 -366
rect -767 -462 -671 -428
rect 671 -462 767 -428
<< viali >>
rect -571 290 -353 324
rect -263 290 -45 324
rect 45 290 263 324
rect 353 290 571 324
rect -633 -231 -599 231
rect -325 -231 -291 231
rect -17 -231 17 231
rect 291 -231 325 231
rect 599 -231 633 231
rect -571 -324 -353 -290
rect -263 -324 -45 -290
rect 45 -324 263 -290
rect 353 -324 571 -290
<< metal1 >>
rect -583 324 -341 330
rect -583 290 -571 324
rect -353 290 -341 324
rect -583 284 -341 290
rect -275 324 -33 330
rect -275 290 -263 324
rect -45 290 -33 324
rect -275 284 -33 290
rect 33 324 275 330
rect 33 290 45 324
rect 263 290 275 324
rect 33 284 275 290
rect 341 324 583 330
rect 341 290 353 324
rect 571 290 583 324
rect 341 284 583 290
rect -639 231 -593 243
rect -639 -231 -633 231
rect -599 -231 -593 231
rect -639 -243 -593 -231
rect -331 231 -285 243
rect -331 -231 -325 231
rect -291 -231 -285 231
rect -331 -243 -285 -231
rect -23 231 23 243
rect -23 -231 -17 231
rect 17 -231 23 231
rect -23 -243 23 -231
rect 285 231 331 243
rect 285 -231 291 231
rect 325 -231 331 231
rect 285 -243 331 -231
rect 593 231 639 243
rect 593 -231 599 231
rect 633 -231 639 231
rect 593 -243 639 -231
rect -583 -290 -341 -284
rect -583 -324 -571 -290
rect -353 -324 -341 -290
rect -583 -330 -341 -324
rect -275 -290 -33 -284
rect -275 -324 -263 -290
rect -45 -324 -33 -290
rect -275 -330 -33 -324
rect 33 -290 275 -284
rect 33 -324 45 -290
rect 263 -324 275 -290
rect 33 -330 275 -324
rect 341 -290 583 -284
rect 341 -324 353 -290
rect 571 -324 583 -290
rect 341 -330 583 -324
<< properties >>
string FIXED_BBOX -750 -445 750 445
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.425 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
