magic
tech sky130A
magscale 1 2
timestamp 1769931968
<< mvnmos >>
rect -287 -450 -187 450
rect -129 -450 -29 450
rect 29 -450 129 450
rect 187 -450 287 450
<< mvndiff >>
rect -345 438 -287 450
rect -345 -438 -333 438
rect -299 -438 -287 438
rect -345 -450 -287 -438
rect -187 438 -129 450
rect -187 -438 -175 438
rect -141 -438 -129 438
rect -187 -450 -129 -438
rect -29 438 29 450
rect -29 -438 -17 438
rect 17 -438 29 438
rect -29 -450 29 -438
rect 129 438 187 450
rect 129 -438 141 438
rect 175 -438 187 438
rect 129 -450 187 -438
rect 287 438 345 450
rect 287 -438 299 438
rect 333 -438 345 438
rect 287 -450 345 -438
<< mvndiffc >>
rect -333 -438 -299 438
rect -175 -438 -141 438
rect -17 -438 17 438
rect 141 -438 175 438
rect 299 -438 333 438
<< poly >>
rect -287 522 -187 538
rect -287 488 -271 522
rect -203 488 -187 522
rect -287 450 -187 488
rect -129 522 -29 538
rect -129 488 -113 522
rect -45 488 -29 522
rect -129 450 -29 488
rect 29 522 129 538
rect 29 488 45 522
rect 113 488 129 522
rect 29 450 129 488
rect 187 522 287 538
rect 187 488 203 522
rect 271 488 287 522
rect 187 450 287 488
rect -287 -488 -187 -450
rect -287 -522 -271 -488
rect -203 -522 -187 -488
rect -287 -538 -187 -522
rect -129 -488 -29 -450
rect -129 -522 -113 -488
rect -45 -522 -29 -488
rect -129 -538 -29 -522
rect 29 -488 129 -450
rect 29 -522 45 -488
rect 113 -522 129 -488
rect 29 -538 129 -522
rect 187 -488 287 -450
rect 187 -522 203 -488
rect 271 -522 287 -488
rect 187 -538 287 -522
<< polycont >>
rect -271 488 -203 522
rect -113 488 -45 522
rect 45 488 113 522
rect 203 488 271 522
rect -271 -522 -203 -488
rect -113 -522 -45 -488
rect 45 -522 113 -488
rect 203 -522 271 -488
<< locali >>
rect -287 488 -271 522
rect -203 488 -187 522
rect -129 488 -113 522
rect -45 488 -29 522
rect 29 488 45 522
rect 113 488 129 522
rect 187 488 203 522
rect 271 488 287 522
rect -333 438 -299 454
rect -333 -454 -299 -438
rect -175 438 -141 454
rect -175 -454 -141 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 141 438 175 454
rect 141 -454 175 -438
rect 299 438 333 454
rect 299 -454 333 -438
rect -287 -522 -271 -488
rect -203 -522 -187 -488
rect -129 -522 -113 -488
rect -45 -522 -29 -488
rect 29 -522 45 -488
rect 113 -522 129 -488
rect 187 -522 203 -488
rect 271 -522 287 -488
<< viali >>
rect -271 488 -203 522
rect -113 488 -45 522
rect 45 488 113 522
rect 203 488 271 522
rect -333 -438 -299 438
rect -175 -438 -141 438
rect -17 -438 17 438
rect 141 -438 175 438
rect 299 -438 333 438
rect -271 -522 -203 -488
rect -113 -522 -45 -488
rect 45 -522 113 -488
rect 203 -522 271 -488
<< metal1 >>
rect -283 522 -191 528
rect -283 488 -271 522
rect -203 488 -191 522
rect -283 482 -191 488
rect -125 522 -33 528
rect -125 488 -113 522
rect -45 488 -33 522
rect -125 482 -33 488
rect 33 522 125 528
rect 33 488 45 522
rect 113 488 125 522
rect 33 482 125 488
rect 191 522 283 528
rect 191 488 203 522
rect 271 488 283 522
rect 191 482 283 488
rect -339 438 -293 450
rect -339 -438 -333 438
rect -299 -438 -293 438
rect -339 -450 -293 -438
rect -181 438 -135 450
rect -181 -438 -175 438
rect -141 -438 -135 438
rect -181 -450 -135 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 135 438 181 450
rect 135 -438 141 438
rect 175 -438 181 438
rect 135 -450 181 -438
rect 293 438 339 450
rect 293 -438 299 438
rect 333 -438 339 438
rect 293 -450 339 -438
rect -283 -488 -191 -482
rect -283 -522 -271 -488
rect -203 -522 -191 -488
rect -283 -528 -191 -522
rect -125 -488 -33 -482
rect -125 -522 -113 -488
rect -45 -522 -33 -488
rect -125 -528 -33 -522
rect 33 -488 125 -482
rect 33 -522 45 -488
rect 113 -522 125 -488
rect 33 -528 125 -522
rect 191 -488 283 -482
rect 191 -522 203 -488
rect 271 -522 283 -488
rect 191 -528 283 -522
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
