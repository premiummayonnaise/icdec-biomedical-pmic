magic
tech sky130A
magscale 1 2
timestamp 1770370310
<< nwell >>
rect -5285 -1328 5285 1328
<< mvpmos >>
rect -5027 -1031 -4927 1031
rect -4869 -1031 -4769 1031
rect -4711 -1031 -4611 1031
rect -4553 -1031 -4453 1031
rect -4395 -1031 -4295 1031
rect -4237 -1031 -4137 1031
rect -4079 -1031 -3979 1031
rect -3921 -1031 -3821 1031
rect -3763 -1031 -3663 1031
rect -3605 -1031 -3505 1031
rect -3447 -1031 -3347 1031
rect -3289 -1031 -3189 1031
rect -3131 -1031 -3031 1031
rect -2973 -1031 -2873 1031
rect -2815 -1031 -2715 1031
rect -2657 -1031 -2557 1031
rect -2499 -1031 -2399 1031
rect -2341 -1031 -2241 1031
rect -2183 -1031 -2083 1031
rect -2025 -1031 -1925 1031
rect -1867 -1031 -1767 1031
rect -1709 -1031 -1609 1031
rect -1551 -1031 -1451 1031
rect -1393 -1031 -1293 1031
rect -1235 -1031 -1135 1031
rect -1077 -1031 -977 1031
rect -919 -1031 -819 1031
rect -761 -1031 -661 1031
rect -603 -1031 -503 1031
rect -445 -1031 -345 1031
rect -287 -1031 -187 1031
rect -129 -1031 -29 1031
rect 29 -1031 129 1031
rect 187 -1031 287 1031
rect 345 -1031 445 1031
rect 503 -1031 603 1031
rect 661 -1031 761 1031
rect 819 -1031 919 1031
rect 977 -1031 1077 1031
rect 1135 -1031 1235 1031
rect 1293 -1031 1393 1031
rect 1451 -1031 1551 1031
rect 1609 -1031 1709 1031
rect 1767 -1031 1867 1031
rect 1925 -1031 2025 1031
rect 2083 -1031 2183 1031
rect 2241 -1031 2341 1031
rect 2399 -1031 2499 1031
rect 2557 -1031 2657 1031
rect 2715 -1031 2815 1031
rect 2873 -1031 2973 1031
rect 3031 -1031 3131 1031
rect 3189 -1031 3289 1031
rect 3347 -1031 3447 1031
rect 3505 -1031 3605 1031
rect 3663 -1031 3763 1031
rect 3821 -1031 3921 1031
rect 3979 -1031 4079 1031
rect 4137 -1031 4237 1031
rect 4295 -1031 4395 1031
rect 4453 -1031 4553 1031
rect 4611 -1031 4711 1031
rect 4769 -1031 4869 1031
rect 4927 -1031 5027 1031
<< mvpdiff >>
rect -5085 1019 -5027 1031
rect -5085 -1019 -5073 1019
rect -5039 -1019 -5027 1019
rect -5085 -1031 -5027 -1019
rect -4927 1019 -4869 1031
rect -4927 -1019 -4915 1019
rect -4881 -1019 -4869 1019
rect -4927 -1031 -4869 -1019
rect -4769 1019 -4711 1031
rect -4769 -1019 -4757 1019
rect -4723 -1019 -4711 1019
rect -4769 -1031 -4711 -1019
rect -4611 1019 -4553 1031
rect -4611 -1019 -4599 1019
rect -4565 -1019 -4553 1019
rect -4611 -1031 -4553 -1019
rect -4453 1019 -4395 1031
rect -4453 -1019 -4441 1019
rect -4407 -1019 -4395 1019
rect -4453 -1031 -4395 -1019
rect -4295 1019 -4237 1031
rect -4295 -1019 -4283 1019
rect -4249 -1019 -4237 1019
rect -4295 -1031 -4237 -1019
rect -4137 1019 -4079 1031
rect -4137 -1019 -4125 1019
rect -4091 -1019 -4079 1019
rect -4137 -1031 -4079 -1019
rect -3979 1019 -3921 1031
rect -3979 -1019 -3967 1019
rect -3933 -1019 -3921 1019
rect -3979 -1031 -3921 -1019
rect -3821 1019 -3763 1031
rect -3821 -1019 -3809 1019
rect -3775 -1019 -3763 1019
rect -3821 -1031 -3763 -1019
rect -3663 1019 -3605 1031
rect -3663 -1019 -3651 1019
rect -3617 -1019 -3605 1019
rect -3663 -1031 -3605 -1019
rect -3505 1019 -3447 1031
rect -3505 -1019 -3493 1019
rect -3459 -1019 -3447 1019
rect -3505 -1031 -3447 -1019
rect -3347 1019 -3289 1031
rect -3347 -1019 -3335 1019
rect -3301 -1019 -3289 1019
rect -3347 -1031 -3289 -1019
rect -3189 1019 -3131 1031
rect -3189 -1019 -3177 1019
rect -3143 -1019 -3131 1019
rect -3189 -1031 -3131 -1019
rect -3031 1019 -2973 1031
rect -3031 -1019 -3019 1019
rect -2985 -1019 -2973 1019
rect -3031 -1031 -2973 -1019
rect -2873 1019 -2815 1031
rect -2873 -1019 -2861 1019
rect -2827 -1019 -2815 1019
rect -2873 -1031 -2815 -1019
rect -2715 1019 -2657 1031
rect -2715 -1019 -2703 1019
rect -2669 -1019 -2657 1019
rect -2715 -1031 -2657 -1019
rect -2557 1019 -2499 1031
rect -2557 -1019 -2545 1019
rect -2511 -1019 -2499 1019
rect -2557 -1031 -2499 -1019
rect -2399 1019 -2341 1031
rect -2399 -1019 -2387 1019
rect -2353 -1019 -2341 1019
rect -2399 -1031 -2341 -1019
rect -2241 1019 -2183 1031
rect -2241 -1019 -2229 1019
rect -2195 -1019 -2183 1019
rect -2241 -1031 -2183 -1019
rect -2083 1019 -2025 1031
rect -2083 -1019 -2071 1019
rect -2037 -1019 -2025 1019
rect -2083 -1031 -2025 -1019
rect -1925 1019 -1867 1031
rect -1925 -1019 -1913 1019
rect -1879 -1019 -1867 1019
rect -1925 -1031 -1867 -1019
rect -1767 1019 -1709 1031
rect -1767 -1019 -1755 1019
rect -1721 -1019 -1709 1019
rect -1767 -1031 -1709 -1019
rect -1609 1019 -1551 1031
rect -1609 -1019 -1597 1019
rect -1563 -1019 -1551 1019
rect -1609 -1031 -1551 -1019
rect -1451 1019 -1393 1031
rect -1451 -1019 -1439 1019
rect -1405 -1019 -1393 1019
rect -1451 -1031 -1393 -1019
rect -1293 1019 -1235 1031
rect -1293 -1019 -1281 1019
rect -1247 -1019 -1235 1019
rect -1293 -1031 -1235 -1019
rect -1135 1019 -1077 1031
rect -1135 -1019 -1123 1019
rect -1089 -1019 -1077 1019
rect -1135 -1031 -1077 -1019
rect -977 1019 -919 1031
rect -977 -1019 -965 1019
rect -931 -1019 -919 1019
rect -977 -1031 -919 -1019
rect -819 1019 -761 1031
rect -819 -1019 -807 1019
rect -773 -1019 -761 1019
rect -819 -1031 -761 -1019
rect -661 1019 -603 1031
rect -661 -1019 -649 1019
rect -615 -1019 -603 1019
rect -661 -1031 -603 -1019
rect -503 1019 -445 1031
rect -503 -1019 -491 1019
rect -457 -1019 -445 1019
rect -503 -1031 -445 -1019
rect -345 1019 -287 1031
rect -345 -1019 -333 1019
rect -299 -1019 -287 1019
rect -345 -1031 -287 -1019
rect -187 1019 -129 1031
rect -187 -1019 -175 1019
rect -141 -1019 -129 1019
rect -187 -1031 -129 -1019
rect -29 1019 29 1031
rect -29 -1019 -17 1019
rect 17 -1019 29 1019
rect -29 -1031 29 -1019
rect 129 1019 187 1031
rect 129 -1019 141 1019
rect 175 -1019 187 1019
rect 129 -1031 187 -1019
rect 287 1019 345 1031
rect 287 -1019 299 1019
rect 333 -1019 345 1019
rect 287 -1031 345 -1019
rect 445 1019 503 1031
rect 445 -1019 457 1019
rect 491 -1019 503 1019
rect 445 -1031 503 -1019
rect 603 1019 661 1031
rect 603 -1019 615 1019
rect 649 -1019 661 1019
rect 603 -1031 661 -1019
rect 761 1019 819 1031
rect 761 -1019 773 1019
rect 807 -1019 819 1019
rect 761 -1031 819 -1019
rect 919 1019 977 1031
rect 919 -1019 931 1019
rect 965 -1019 977 1019
rect 919 -1031 977 -1019
rect 1077 1019 1135 1031
rect 1077 -1019 1089 1019
rect 1123 -1019 1135 1019
rect 1077 -1031 1135 -1019
rect 1235 1019 1293 1031
rect 1235 -1019 1247 1019
rect 1281 -1019 1293 1019
rect 1235 -1031 1293 -1019
rect 1393 1019 1451 1031
rect 1393 -1019 1405 1019
rect 1439 -1019 1451 1019
rect 1393 -1031 1451 -1019
rect 1551 1019 1609 1031
rect 1551 -1019 1563 1019
rect 1597 -1019 1609 1019
rect 1551 -1031 1609 -1019
rect 1709 1019 1767 1031
rect 1709 -1019 1721 1019
rect 1755 -1019 1767 1019
rect 1709 -1031 1767 -1019
rect 1867 1019 1925 1031
rect 1867 -1019 1879 1019
rect 1913 -1019 1925 1019
rect 1867 -1031 1925 -1019
rect 2025 1019 2083 1031
rect 2025 -1019 2037 1019
rect 2071 -1019 2083 1019
rect 2025 -1031 2083 -1019
rect 2183 1019 2241 1031
rect 2183 -1019 2195 1019
rect 2229 -1019 2241 1019
rect 2183 -1031 2241 -1019
rect 2341 1019 2399 1031
rect 2341 -1019 2353 1019
rect 2387 -1019 2399 1019
rect 2341 -1031 2399 -1019
rect 2499 1019 2557 1031
rect 2499 -1019 2511 1019
rect 2545 -1019 2557 1019
rect 2499 -1031 2557 -1019
rect 2657 1019 2715 1031
rect 2657 -1019 2669 1019
rect 2703 -1019 2715 1019
rect 2657 -1031 2715 -1019
rect 2815 1019 2873 1031
rect 2815 -1019 2827 1019
rect 2861 -1019 2873 1019
rect 2815 -1031 2873 -1019
rect 2973 1019 3031 1031
rect 2973 -1019 2985 1019
rect 3019 -1019 3031 1019
rect 2973 -1031 3031 -1019
rect 3131 1019 3189 1031
rect 3131 -1019 3143 1019
rect 3177 -1019 3189 1019
rect 3131 -1031 3189 -1019
rect 3289 1019 3347 1031
rect 3289 -1019 3301 1019
rect 3335 -1019 3347 1019
rect 3289 -1031 3347 -1019
rect 3447 1019 3505 1031
rect 3447 -1019 3459 1019
rect 3493 -1019 3505 1019
rect 3447 -1031 3505 -1019
rect 3605 1019 3663 1031
rect 3605 -1019 3617 1019
rect 3651 -1019 3663 1019
rect 3605 -1031 3663 -1019
rect 3763 1019 3821 1031
rect 3763 -1019 3775 1019
rect 3809 -1019 3821 1019
rect 3763 -1031 3821 -1019
rect 3921 1019 3979 1031
rect 3921 -1019 3933 1019
rect 3967 -1019 3979 1019
rect 3921 -1031 3979 -1019
rect 4079 1019 4137 1031
rect 4079 -1019 4091 1019
rect 4125 -1019 4137 1019
rect 4079 -1031 4137 -1019
rect 4237 1019 4295 1031
rect 4237 -1019 4249 1019
rect 4283 -1019 4295 1019
rect 4237 -1031 4295 -1019
rect 4395 1019 4453 1031
rect 4395 -1019 4407 1019
rect 4441 -1019 4453 1019
rect 4395 -1031 4453 -1019
rect 4553 1019 4611 1031
rect 4553 -1019 4565 1019
rect 4599 -1019 4611 1019
rect 4553 -1031 4611 -1019
rect 4711 1019 4769 1031
rect 4711 -1019 4723 1019
rect 4757 -1019 4769 1019
rect 4711 -1031 4769 -1019
rect 4869 1019 4927 1031
rect 4869 -1019 4881 1019
rect 4915 -1019 4927 1019
rect 4869 -1031 4927 -1019
rect 5027 1019 5085 1031
rect 5027 -1019 5039 1019
rect 5073 -1019 5085 1019
rect 5027 -1031 5085 -1019
<< mvpdiffc >>
rect -5073 -1019 -5039 1019
rect -4915 -1019 -4881 1019
rect -4757 -1019 -4723 1019
rect -4599 -1019 -4565 1019
rect -4441 -1019 -4407 1019
rect -4283 -1019 -4249 1019
rect -4125 -1019 -4091 1019
rect -3967 -1019 -3933 1019
rect -3809 -1019 -3775 1019
rect -3651 -1019 -3617 1019
rect -3493 -1019 -3459 1019
rect -3335 -1019 -3301 1019
rect -3177 -1019 -3143 1019
rect -3019 -1019 -2985 1019
rect -2861 -1019 -2827 1019
rect -2703 -1019 -2669 1019
rect -2545 -1019 -2511 1019
rect -2387 -1019 -2353 1019
rect -2229 -1019 -2195 1019
rect -2071 -1019 -2037 1019
rect -1913 -1019 -1879 1019
rect -1755 -1019 -1721 1019
rect -1597 -1019 -1563 1019
rect -1439 -1019 -1405 1019
rect -1281 -1019 -1247 1019
rect -1123 -1019 -1089 1019
rect -965 -1019 -931 1019
rect -807 -1019 -773 1019
rect -649 -1019 -615 1019
rect -491 -1019 -457 1019
rect -333 -1019 -299 1019
rect -175 -1019 -141 1019
rect -17 -1019 17 1019
rect 141 -1019 175 1019
rect 299 -1019 333 1019
rect 457 -1019 491 1019
rect 615 -1019 649 1019
rect 773 -1019 807 1019
rect 931 -1019 965 1019
rect 1089 -1019 1123 1019
rect 1247 -1019 1281 1019
rect 1405 -1019 1439 1019
rect 1563 -1019 1597 1019
rect 1721 -1019 1755 1019
rect 1879 -1019 1913 1019
rect 2037 -1019 2071 1019
rect 2195 -1019 2229 1019
rect 2353 -1019 2387 1019
rect 2511 -1019 2545 1019
rect 2669 -1019 2703 1019
rect 2827 -1019 2861 1019
rect 2985 -1019 3019 1019
rect 3143 -1019 3177 1019
rect 3301 -1019 3335 1019
rect 3459 -1019 3493 1019
rect 3617 -1019 3651 1019
rect 3775 -1019 3809 1019
rect 3933 -1019 3967 1019
rect 4091 -1019 4125 1019
rect 4249 -1019 4283 1019
rect 4407 -1019 4441 1019
rect 4565 -1019 4599 1019
rect 4723 -1019 4757 1019
rect 4881 -1019 4915 1019
rect 5039 -1019 5073 1019
<< mvnsubdiff >>
rect -5219 1250 5219 1262
rect -5219 1216 -5111 1250
rect 5111 1216 5219 1250
rect -5219 1204 5219 1216
rect -5219 1154 -5161 1204
rect -5219 -1154 -5207 1154
rect -5173 -1154 -5161 1154
rect 5161 1154 5219 1204
rect -5219 -1204 -5161 -1154
rect 5161 -1154 5173 1154
rect 5207 -1154 5219 1154
rect 5161 -1204 5219 -1154
rect -5219 -1216 5219 -1204
rect -5219 -1250 -5111 -1216
rect 5111 -1250 5219 -1216
rect -5219 -1262 5219 -1250
<< mvnsubdiffcont >>
rect -5111 1216 5111 1250
rect -5207 -1154 -5173 1154
rect 5173 -1154 5207 1154
rect -5111 -1250 5111 -1216
<< poly >>
rect -5027 1112 -4927 1128
rect -5027 1078 -5011 1112
rect -4943 1078 -4927 1112
rect -5027 1031 -4927 1078
rect -4869 1112 -4769 1128
rect -4869 1078 -4853 1112
rect -4785 1078 -4769 1112
rect -4869 1031 -4769 1078
rect -4711 1112 -4611 1128
rect -4711 1078 -4695 1112
rect -4627 1078 -4611 1112
rect -4711 1031 -4611 1078
rect -4553 1112 -4453 1128
rect -4553 1078 -4537 1112
rect -4469 1078 -4453 1112
rect -4553 1031 -4453 1078
rect -4395 1112 -4295 1128
rect -4395 1078 -4379 1112
rect -4311 1078 -4295 1112
rect -4395 1031 -4295 1078
rect -4237 1112 -4137 1128
rect -4237 1078 -4221 1112
rect -4153 1078 -4137 1112
rect -4237 1031 -4137 1078
rect -4079 1112 -3979 1128
rect -4079 1078 -4063 1112
rect -3995 1078 -3979 1112
rect -4079 1031 -3979 1078
rect -3921 1112 -3821 1128
rect -3921 1078 -3905 1112
rect -3837 1078 -3821 1112
rect -3921 1031 -3821 1078
rect -3763 1112 -3663 1128
rect -3763 1078 -3747 1112
rect -3679 1078 -3663 1112
rect -3763 1031 -3663 1078
rect -3605 1112 -3505 1128
rect -3605 1078 -3589 1112
rect -3521 1078 -3505 1112
rect -3605 1031 -3505 1078
rect -3447 1112 -3347 1128
rect -3447 1078 -3431 1112
rect -3363 1078 -3347 1112
rect -3447 1031 -3347 1078
rect -3289 1112 -3189 1128
rect -3289 1078 -3273 1112
rect -3205 1078 -3189 1112
rect -3289 1031 -3189 1078
rect -3131 1112 -3031 1128
rect -3131 1078 -3115 1112
rect -3047 1078 -3031 1112
rect -3131 1031 -3031 1078
rect -2973 1112 -2873 1128
rect -2973 1078 -2957 1112
rect -2889 1078 -2873 1112
rect -2973 1031 -2873 1078
rect -2815 1112 -2715 1128
rect -2815 1078 -2799 1112
rect -2731 1078 -2715 1112
rect -2815 1031 -2715 1078
rect -2657 1112 -2557 1128
rect -2657 1078 -2641 1112
rect -2573 1078 -2557 1112
rect -2657 1031 -2557 1078
rect -2499 1112 -2399 1128
rect -2499 1078 -2483 1112
rect -2415 1078 -2399 1112
rect -2499 1031 -2399 1078
rect -2341 1112 -2241 1128
rect -2341 1078 -2325 1112
rect -2257 1078 -2241 1112
rect -2341 1031 -2241 1078
rect -2183 1112 -2083 1128
rect -2183 1078 -2167 1112
rect -2099 1078 -2083 1112
rect -2183 1031 -2083 1078
rect -2025 1112 -1925 1128
rect -2025 1078 -2009 1112
rect -1941 1078 -1925 1112
rect -2025 1031 -1925 1078
rect -1867 1112 -1767 1128
rect -1867 1078 -1851 1112
rect -1783 1078 -1767 1112
rect -1867 1031 -1767 1078
rect -1709 1112 -1609 1128
rect -1709 1078 -1693 1112
rect -1625 1078 -1609 1112
rect -1709 1031 -1609 1078
rect -1551 1112 -1451 1128
rect -1551 1078 -1535 1112
rect -1467 1078 -1451 1112
rect -1551 1031 -1451 1078
rect -1393 1112 -1293 1128
rect -1393 1078 -1377 1112
rect -1309 1078 -1293 1112
rect -1393 1031 -1293 1078
rect -1235 1112 -1135 1128
rect -1235 1078 -1219 1112
rect -1151 1078 -1135 1112
rect -1235 1031 -1135 1078
rect -1077 1112 -977 1128
rect -1077 1078 -1061 1112
rect -993 1078 -977 1112
rect -1077 1031 -977 1078
rect -919 1112 -819 1128
rect -919 1078 -903 1112
rect -835 1078 -819 1112
rect -919 1031 -819 1078
rect -761 1112 -661 1128
rect -761 1078 -745 1112
rect -677 1078 -661 1112
rect -761 1031 -661 1078
rect -603 1112 -503 1128
rect -603 1078 -587 1112
rect -519 1078 -503 1112
rect -603 1031 -503 1078
rect -445 1112 -345 1128
rect -445 1078 -429 1112
rect -361 1078 -345 1112
rect -445 1031 -345 1078
rect -287 1112 -187 1128
rect -287 1078 -271 1112
rect -203 1078 -187 1112
rect -287 1031 -187 1078
rect -129 1112 -29 1128
rect -129 1078 -113 1112
rect -45 1078 -29 1112
rect -129 1031 -29 1078
rect 29 1112 129 1128
rect 29 1078 45 1112
rect 113 1078 129 1112
rect 29 1031 129 1078
rect 187 1112 287 1128
rect 187 1078 203 1112
rect 271 1078 287 1112
rect 187 1031 287 1078
rect 345 1112 445 1128
rect 345 1078 361 1112
rect 429 1078 445 1112
rect 345 1031 445 1078
rect 503 1112 603 1128
rect 503 1078 519 1112
rect 587 1078 603 1112
rect 503 1031 603 1078
rect 661 1112 761 1128
rect 661 1078 677 1112
rect 745 1078 761 1112
rect 661 1031 761 1078
rect 819 1112 919 1128
rect 819 1078 835 1112
rect 903 1078 919 1112
rect 819 1031 919 1078
rect 977 1112 1077 1128
rect 977 1078 993 1112
rect 1061 1078 1077 1112
rect 977 1031 1077 1078
rect 1135 1112 1235 1128
rect 1135 1078 1151 1112
rect 1219 1078 1235 1112
rect 1135 1031 1235 1078
rect 1293 1112 1393 1128
rect 1293 1078 1309 1112
rect 1377 1078 1393 1112
rect 1293 1031 1393 1078
rect 1451 1112 1551 1128
rect 1451 1078 1467 1112
rect 1535 1078 1551 1112
rect 1451 1031 1551 1078
rect 1609 1112 1709 1128
rect 1609 1078 1625 1112
rect 1693 1078 1709 1112
rect 1609 1031 1709 1078
rect 1767 1112 1867 1128
rect 1767 1078 1783 1112
rect 1851 1078 1867 1112
rect 1767 1031 1867 1078
rect 1925 1112 2025 1128
rect 1925 1078 1941 1112
rect 2009 1078 2025 1112
rect 1925 1031 2025 1078
rect 2083 1112 2183 1128
rect 2083 1078 2099 1112
rect 2167 1078 2183 1112
rect 2083 1031 2183 1078
rect 2241 1112 2341 1128
rect 2241 1078 2257 1112
rect 2325 1078 2341 1112
rect 2241 1031 2341 1078
rect 2399 1112 2499 1128
rect 2399 1078 2415 1112
rect 2483 1078 2499 1112
rect 2399 1031 2499 1078
rect 2557 1112 2657 1128
rect 2557 1078 2573 1112
rect 2641 1078 2657 1112
rect 2557 1031 2657 1078
rect 2715 1112 2815 1128
rect 2715 1078 2731 1112
rect 2799 1078 2815 1112
rect 2715 1031 2815 1078
rect 2873 1112 2973 1128
rect 2873 1078 2889 1112
rect 2957 1078 2973 1112
rect 2873 1031 2973 1078
rect 3031 1112 3131 1128
rect 3031 1078 3047 1112
rect 3115 1078 3131 1112
rect 3031 1031 3131 1078
rect 3189 1112 3289 1128
rect 3189 1078 3205 1112
rect 3273 1078 3289 1112
rect 3189 1031 3289 1078
rect 3347 1112 3447 1128
rect 3347 1078 3363 1112
rect 3431 1078 3447 1112
rect 3347 1031 3447 1078
rect 3505 1112 3605 1128
rect 3505 1078 3521 1112
rect 3589 1078 3605 1112
rect 3505 1031 3605 1078
rect 3663 1112 3763 1128
rect 3663 1078 3679 1112
rect 3747 1078 3763 1112
rect 3663 1031 3763 1078
rect 3821 1112 3921 1128
rect 3821 1078 3837 1112
rect 3905 1078 3921 1112
rect 3821 1031 3921 1078
rect 3979 1112 4079 1128
rect 3979 1078 3995 1112
rect 4063 1078 4079 1112
rect 3979 1031 4079 1078
rect 4137 1112 4237 1128
rect 4137 1078 4153 1112
rect 4221 1078 4237 1112
rect 4137 1031 4237 1078
rect 4295 1112 4395 1128
rect 4295 1078 4311 1112
rect 4379 1078 4395 1112
rect 4295 1031 4395 1078
rect 4453 1112 4553 1128
rect 4453 1078 4469 1112
rect 4537 1078 4553 1112
rect 4453 1031 4553 1078
rect 4611 1112 4711 1128
rect 4611 1078 4627 1112
rect 4695 1078 4711 1112
rect 4611 1031 4711 1078
rect 4769 1112 4869 1128
rect 4769 1078 4785 1112
rect 4853 1078 4869 1112
rect 4769 1031 4869 1078
rect 4927 1112 5027 1128
rect 4927 1078 4943 1112
rect 5011 1078 5027 1112
rect 4927 1031 5027 1078
rect -5027 -1078 -4927 -1031
rect -5027 -1112 -5011 -1078
rect -4943 -1112 -4927 -1078
rect -5027 -1128 -4927 -1112
rect -4869 -1078 -4769 -1031
rect -4869 -1112 -4853 -1078
rect -4785 -1112 -4769 -1078
rect -4869 -1128 -4769 -1112
rect -4711 -1078 -4611 -1031
rect -4711 -1112 -4695 -1078
rect -4627 -1112 -4611 -1078
rect -4711 -1128 -4611 -1112
rect -4553 -1078 -4453 -1031
rect -4553 -1112 -4537 -1078
rect -4469 -1112 -4453 -1078
rect -4553 -1128 -4453 -1112
rect -4395 -1078 -4295 -1031
rect -4395 -1112 -4379 -1078
rect -4311 -1112 -4295 -1078
rect -4395 -1128 -4295 -1112
rect -4237 -1078 -4137 -1031
rect -4237 -1112 -4221 -1078
rect -4153 -1112 -4137 -1078
rect -4237 -1128 -4137 -1112
rect -4079 -1078 -3979 -1031
rect -4079 -1112 -4063 -1078
rect -3995 -1112 -3979 -1078
rect -4079 -1128 -3979 -1112
rect -3921 -1078 -3821 -1031
rect -3921 -1112 -3905 -1078
rect -3837 -1112 -3821 -1078
rect -3921 -1128 -3821 -1112
rect -3763 -1078 -3663 -1031
rect -3763 -1112 -3747 -1078
rect -3679 -1112 -3663 -1078
rect -3763 -1128 -3663 -1112
rect -3605 -1078 -3505 -1031
rect -3605 -1112 -3589 -1078
rect -3521 -1112 -3505 -1078
rect -3605 -1128 -3505 -1112
rect -3447 -1078 -3347 -1031
rect -3447 -1112 -3431 -1078
rect -3363 -1112 -3347 -1078
rect -3447 -1128 -3347 -1112
rect -3289 -1078 -3189 -1031
rect -3289 -1112 -3273 -1078
rect -3205 -1112 -3189 -1078
rect -3289 -1128 -3189 -1112
rect -3131 -1078 -3031 -1031
rect -3131 -1112 -3115 -1078
rect -3047 -1112 -3031 -1078
rect -3131 -1128 -3031 -1112
rect -2973 -1078 -2873 -1031
rect -2973 -1112 -2957 -1078
rect -2889 -1112 -2873 -1078
rect -2973 -1128 -2873 -1112
rect -2815 -1078 -2715 -1031
rect -2815 -1112 -2799 -1078
rect -2731 -1112 -2715 -1078
rect -2815 -1128 -2715 -1112
rect -2657 -1078 -2557 -1031
rect -2657 -1112 -2641 -1078
rect -2573 -1112 -2557 -1078
rect -2657 -1128 -2557 -1112
rect -2499 -1078 -2399 -1031
rect -2499 -1112 -2483 -1078
rect -2415 -1112 -2399 -1078
rect -2499 -1128 -2399 -1112
rect -2341 -1078 -2241 -1031
rect -2341 -1112 -2325 -1078
rect -2257 -1112 -2241 -1078
rect -2341 -1128 -2241 -1112
rect -2183 -1078 -2083 -1031
rect -2183 -1112 -2167 -1078
rect -2099 -1112 -2083 -1078
rect -2183 -1128 -2083 -1112
rect -2025 -1078 -1925 -1031
rect -2025 -1112 -2009 -1078
rect -1941 -1112 -1925 -1078
rect -2025 -1128 -1925 -1112
rect -1867 -1078 -1767 -1031
rect -1867 -1112 -1851 -1078
rect -1783 -1112 -1767 -1078
rect -1867 -1128 -1767 -1112
rect -1709 -1078 -1609 -1031
rect -1709 -1112 -1693 -1078
rect -1625 -1112 -1609 -1078
rect -1709 -1128 -1609 -1112
rect -1551 -1078 -1451 -1031
rect -1551 -1112 -1535 -1078
rect -1467 -1112 -1451 -1078
rect -1551 -1128 -1451 -1112
rect -1393 -1078 -1293 -1031
rect -1393 -1112 -1377 -1078
rect -1309 -1112 -1293 -1078
rect -1393 -1128 -1293 -1112
rect -1235 -1078 -1135 -1031
rect -1235 -1112 -1219 -1078
rect -1151 -1112 -1135 -1078
rect -1235 -1128 -1135 -1112
rect -1077 -1078 -977 -1031
rect -1077 -1112 -1061 -1078
rect -993 -1112 -977 -1078
rect -1077 -1128 -977 -1112
rect -919 -1078 -819 -1031
rect -919 -1112 -903 -1078
rect -835 -1112 -819 -1078
rect -919 -1128 -819 -1112
rect -761 -1078 -661 -1031
rect -761 -1112 -745 -1078
rect -677 -1112 -661 -1078
rect -761 -1128 -661 -1112
rect -603 -1078 -503 -1031
rect -603 -1112 -587 -1078
rect -519 -1112 -503 -1078
rect -603 -1128 -503 -1112
rect -445 -1078 -345 -1031
rect -445 -1112 -429 -1078
rect -361 -1112 -345 -1078
rect -445 -1128 -345 -1112
rect -287 -1078 -187 -1031
rect -287 -1112 -271 -1078
rect -203 -1112 -187 -1078
rect -287 -1128 -187 -1112
rect -129 -1078 -29 -1031
rect -129 -1112 -113 -1078
rect -45 -1112 -29 -1078
rect -129 -1128 -29 -1112
rect 29 -1078 129 -1031
rect 29 -1112 45 -1078
rect 113 -1112 129 -1078
rect 29 -1128 129 -1112
rect 187 -1078 287 -1031
rect 187 -1112 203 -1078
rect 271 -1112 287 -1078
rect 187 -1128 287 -1112
rect 345 -1078 445 -1031
rect 345 -1112 361 -1078
rect 429 -1112 445 -1078
rect 345 -1128 445 -1112
rect 503 -1078 603 -1031
rect 503 -1112 519 -1078
rect 587 -1112 603 -1078
rect 503 -1128 603 -1112
rect 661 -1078 761 -1031
rect 661 -1112 677 -1078
rect 745 -1112 761 -1078
rect 661 -1128 761 -1112
rect 819 -1078 919 -1031
rect 819 -1112 835 -1078
rect 903 -1112 919 -1078
rect 819 -1128 919 -1112
rect 977 -1078 1077 -1031
rect 977 -1112 993 -1078
rect 1061 -1112 1077 -1078
rect 977 -1128 1077 -1112
rect 1135 -1078 1235 -1031
rect 1135 -1112 1151 -1078
rect 1219 -1112 1235 -1078
rect 1135 -1128 1235 -1112
rect 1293 -1078 1393 -1031
rect 1293 -1112 1309 -1078
rect 1377 -1112 1393 -1078
rect 1293 -1128 1393 -1112
rect 1451 -1078 1551 -1031
rect 1451 -1112 1467 -1078
rect 1535 -1112 1551 -1078
rect 1451 -1128 1551 -1112
rect 1609 -1078 1709 -1031
rect 1609 -1112 1625 -1078
rect 1693 -1112 1709 -1078
rect 1609 -1128 1709 -1112
rect 1767 -1078 1867 -1031
rect 1767 -1112 1783 -1078
rect 1851 -1112 1867 -1078
rect 1767 -1128 1867 -1112
rect 1925 -1078 2025 -1031
rect 1925 -1112 1941 -1078
rect 2009 -1112 2025 -1078
rect 1925 -1128 2025 -1112
rect 2083 -1078 2183 -1031
rect 2083 -1112 2099 -1078
rect 2167 -1112 2183 -1078
rect 2083 -1128 2183 -1112
rect 2241 -1078 2341 -1031
rect 2241 -1112 2257 -1078
rect 2325 -1112 2341 -1078
rect 2241 -1128 2341 -1112
rect 2399 -1078 2499 -1031
rect 2399 -1112 2415 -1078
rect 2483 -1112 2499 -1078
rect 2399 -1128 2499 -1112
rect 2557 -1078 2657 -1031
rect 2557 -1112 2573 -1078
rect 2641 -1112 2657 -1078
rect 2557 -1128 2657 -1112
rect 2715 -1078 2815 -1031
rect 2715 -1112 2731 -1078
rect 2799 -1112 2815 -1078
rect 2715 -1128 2815 -1112
rect 2873 -1078 2973 -1031
rect 2873 -1112 2889 -1078
rect 2957 -1112 2973 -1078
rect 2873 -1128 2973 -1112
rect 3031 -1078 3131 -1031
rect 3031 -1112 3047 -1078
rect 3115 -1112 3131 -1078
rect 3031 -1128 3131 -1112
rect 3189 -1078 3289 -1031
rect 3189 -1112 3205 -1078
rect 3273 -1112 3289 -1078
rect 3189 -1128 3289 -1112
rect 3347 -1078 3447 -1031
rect 3347 -1112 3363 -1078
rect 3431 -1112 3447 -1078
rect 3347 -1128 3447 -1112
rect 3505 -1078 3605 -1031
rect 3505 -1112 3521 -1078
rect 3589 -1112 3605 -1078
rect 3505 -1128 3605 -1112
rect 3663 -1078 3763 -1031
rect 3663 -1112 3679 -1078
rect 3747 -1112 3763 -1078
rect 3663 -1128 3763 -1112
rect 3821 -1078 3921 -1031
rect 3821 -1112 3837 -1078
rect 3905 -1112 3921 -1078
rect 3821 -1128 3921 -1112
rect 3979 -1078 4079 -1031
rect 3979 -1112 3995 -1078
rect 4063 -1112 4079 -1078
rect 3979 -1128 4079 -1112
rect 4137 -1078 4237 -1031
rect 4137 -1112 4153 -1078
rect 4221 -1112 4237 -1078
rect 4137 -1128 4237 -1112
rect 4295 -1078 4395 -1031
rect 4295 -1112 4311 -1078
rect 4379 -1112 4395 -1078
rect 4295 -1128 4395 -1112
rect 4453 -1078 4553 -1031
rect 4453 -1112 4469 -1078
rect 4537 -1112 4553 -1078
rect 4453 -1128 4553 -1112
rect 4611 -1078 4711 -1031
rect 4611 -1112 4627 -1078
rect 4695 -1112 4711 -1078
rect 4611 -1128 4711 -1112
rect 4769 -1078 4869 -1031
rect 4769 -1112 4785 -1078
rect 4853 -1112 4869 -1078
rect 4769 -1128 4869 -1112
rect 4927 -1078 5027 -1031
rect 4927 -1112 4943 -1078
rect 5011 -1112 5027 -1078
rect 4927 -1128 5027 -1112
<< polycont >>
rect -5011 1078 -4943 1112
rect -4853 1078 -4785 1112
rect -4695 1078 -4627 1112
rect -4537 1078 -4469 1112
rect -4379 1078 -4311 1112
rect -4221 1078 -4153 1112
rect -4063 1078 -3995 1112
rect -3905 1078 -3837 1112
rect -3747 1078 -3679 1112
rect -3589 1078 -3521 1112
rect -3431 1078 -3363 1112
rect -3273 1078 -3205 1112
rect -3115 1078 -3047 1112
rect -2957 1078 -2889 1112
rect -2799 1078 -2731 1112
rect -2641 1078 -2573 1112
rect -2483 1078 -2415 1112
rect -2325 1078 -2257 1112
rect -2167 1078 -2099 1112
rect -2009 1078 -1941 1112
rect -1851 1078 -1783 1112
rect -1693 1078 -1625 1112
rect -1535 1078 -1467 1112
rect -1377 1078 -1309 1112
rect -1219 1078 -1151 1112
rect -1061 1078 -993 1112
rect -903 1078 -835 1112
rect -745 1078 -677 1112
rect -587 1078 -519 1112
rect -429 1078 -361 1112
rect -271 1078 -203 1112
rect -113 1078 -45 1112
rect 45 1078 113 1112
rect 203 1078 271 1112
rect 361 1078 429 1112
rect 519 1078 587 1112
rect 677 1078 745 1112
rect 835 1078 903 1112
rect 993 1078 1061 1112
rect 1151 1078 1219 1112
rect 1309 1078 1377 1112
rect 1467 1078 1535 1112
rect 1625 1078 1693 1112
rect 1783 1078 1851 1112
rect 1941 1078 2009 1112
rect 2099 1078 2167 1112
rect 2257 1078 2325 1112
rect 2415 1078 2483 1112
rect 2573 1078 2641 1112
rect 2731 1078 2799 1112
rect 2889 1078 2957 1112
rect 3047 1078 3115 1112
rect 3205 1078 3273 1112
rect 3363 1078 3431 1112
rect 3521 1078 3589 1112
rect 3679 1078 3747 1112
rect 3837 1078 3905 1112
rect 3995 1078 4063 1112
rect 4153 1078 4221 1112
rect 4311 1078 4379 1112
rect 4469 1078 4537 1112
rect 4627 1078 4695 1112
rect 4785 1078 4853 1112
rect 4943 1078 5011 1112
rect -5011 -1112 -4943 -1078
rect -4853 -1112 -4785 -1078
rect -4695 -1112 -4627 -1078
rect -4537 -1112 -4469 -1078
rect -4379 -1112 -4311 -1078
rect -4221 -1112 -4153 -1078
rect -4063 -1112 -3995 -1078
rect -3905 -1112 -3837 -1078
rect -3747 -1112 -3679 -1078
rect -3589 -1112 -3521 -1078
rect -3431 -1112 -3363 -1078
rect -3273 -1112 -3205 -1078
rect -3115 -1112 -3047 -1078
rect -2957 -1112 -2889 -1078
rect -2799 -1112 -2731 -1078
rect -2641 -1112 -2573 -1078
rect -2483 -1112 -2415 -1078
rect -2325 -1112 -2257 -1078
rect -2167 -1112 -2099 -1078
rect -2009 -1112 -1941 -1078
rect -1851 -1112 -1783 -1078
rect -1693 -1112 -1625 -1078
rect -1535 -1112 -1467 -1078
rect -1377 -1112 -1309 -1078
rect -1219 -1112 -1151 -1078
rect -1061 -1112 -993 -1078
rect -903 -1112 -835 -1078
rect -745 -1112 -677 -1078
rect -587 -1112 -519 -1078
rect -429 -1112 -361 -1078
rect -271 -1112 -203 -1078
rect -113 -1112 -45 -1078
rect 45 -1112 113 -1078
rect 203 -1112 271 -1078
rect 361 -1112 429 -1078
rect 519 -1112 587 -1078
rect 677 -1112 745 -1078
rect 835 -1112 903 -1078
rect 993 -1112 1061 -1078
rect 1151 -1112 1219 -1078
rect 1309 -1112 1377 -1078
rect 1467 -1112 1535 -1078
rect 1625 -1112 1693 -1078
rect 1783 -1112 1851 -1078
rect 1941 -1112 2009 -1078
rect 2099 -1112 2167 -1078
rect 2257 -1112 2325 -1078
rect 2415 -1112 2483 -1078
rect 2573 -1112 2641 -1078
rect 2731 -1112 2799 -1078
rect 2889 -1112 2957 -1078
rect 3047 -1112 3115 -1078
rect 3205 -1112 3273 -1078
rect 3363 -1112 3431 -1078
rect 3521 -1112 3589 -1078
rect 3679 -1112 3747 -1078
rect 3837 -1112 3905 -1078
rect 3995 -1112 4063 -1078
rect 4153 -1112 4221 -1078
rect 4311 -1112 4379 -1078
rect 4469 -1112 4537 -1078
rect 4627 -1112 4695 -1078
rect 4785 -1112 4853 -1078
rect 4943 -1112 5011 -1078
<< locali >>
rect -5207 1216 -5111 1250
rect 5111 1216 5207 1250
rect -5207 1154 -5173 1216
rect 5173 1154 5207 1216
rect -5027 1078 -5011 1112
rect -4943 1078 -4927 1112
rect -4869 1078 -4853 1112
rect -4785 1078 -4769 1112
rect -4711 1078 -4695 1112
rect -4627 1078 -4611 1112
rect -4553 1078 -4537 1112
rect -4469 1078 -4453 1112
rect -4395 1078 -4379 1112
rect -4311 1078 -4295 1112
rect -4237 1078 -4221 1112
rect -4153 1078 -4137 1112
rect -4079 1078 -4063 1112
rect -3995 1078 -3979 1112
rect -3921 1078 -3905 1112
rect -3837 1078 -3821 1112
rect -3763 1078 -3747 1112
rect -3679 1078 -3663 1112
rect -3605 1078 -3589 1112
rect -3521 1078 -3505 1112
rect -3447 1078 -3431 1112
rect -3363 1078 -3347 1112
rect -3289 1078 -3273 1112
rect -3205 1078 -3189 1112
rect -3131 1078 -3115 1112
rect -3047 1078 -3031 1112
rect -2973 1078 -2957 1112
rect -2889 1078 -2873 1112
rect -2815 1078 -2799 1112
rect -2731 1078 -2715 1112
rect -2657 1078 -2641 1112
rect -2573 1078 -2557 1112
rect -2499 1078 -2483 1112
rect -2415 1078 -2399 1112
rect -2341 1078 -2325 1112
rect -2257 1078 -2241 1112
rect -2183 1078 -2167 1112
rect -2099 1078 -2083 1112
rect -2025 1078 -2009 1112
rect -1941 1078 -1925 1112
rect -1867 1078 -1851 1112
rect -1783 1078 -1767 1112
rect -1709 1078 -1693 1112
rect -1625 1078 -1609 1112
rect -1551 1078 -1535 1112
rect -1467 1078 -1451 1112
rect -1393 1078 -1377 1112
rect -1309 1078 -1293 1112
rect -1235 1078 -1219 1112
rect -1151 1078 -1135 1112
rect -1077 1078 -1061 1112
rect -993 1078 -977 1112
rect -919 1078 -903 1112
rect -835 1078 -819 1112
rect -761 1078 -745 1112
rect -677 1078 -661 1112
rect -603 1078 -587 1112
rect -519 1078 -503 1112
rect -445 1078 -429 1112
rect -361 1078 -345 1112
rect -287 1078 -271 1112
rect -203 1078 -187 1112
rect -129 1078 -113 1112
rect -45 1078 -29 1112
rect 29 1078 45 1112
rect 113 1078 129 1112
rect 187 1078 203 1112
rect 271 1078 287 1112
rect 345 1078 361 1112
rect 429 1078 445 1112
rect 503 1078 519 1112
rect 587 1078 603 1112
rect 661 1078 677 1112
rect 745 1078 761 1112
rect 819 1078 835 1112
rect 903 1078 919 1112
rect 977 1078 993 1112
rect 1061 1078 1077 1112
rect 1135 1078 1151 1112
rect 1219 1078 1235 1112
rect 1293 1078 1309 1112
rect 1377 1078 1393 1112
rect 1451 1078 1467 1112
rect 1535 1078 1551 1112
rect 1609 1078 1625 1112
rect 1693 1078 1709 1112
rect 1767 1078 1783 1112
rect 1851 1078 1867 1112
rect 1925 1078 1941 1112
rect 2009 1078 2025 1112
rect 2083 1078 2099 1112
rect 2167 1078 2183 1112
rect 2241 1078 2257 1112
rect 2325 1078 2341 1112
rect 2399 1078 2415 1112
rect 2483 1078 2499 1112
rect 2557 1078 2573 1112
rect 2641 1078 2657 1112
rect 2715 1078 2731 1112
rect 2799 1078 2815 1112
rect 2873 1078 2889 1112
rect 2957 1078 2973 1112
rect 3031 1078 3047 1112
rect 3115 1078 3131 1112
rect 3189 1078 3205 1112
rect 3273 1078 3289 1112
rect 3347 1078 3363 1112
rect 3431 1078 3447 1112
rect 3505 1078 3521 1112
rect 3589 1078 3605 1112
rect 3663 1078 3679 1112
rect 3747 1078 3763 1112
rect 3821 1078 3837 1112
rect 3905 1078 3921 1112
rect 3979 1078 3995 1112
rect 4063 1078 4079 1112
rect 4137 1078 4153 1112
rect 4221 1078 4237 1112
rect 4295 1078 4311 1112
rect 4379 1078 4395 1112
rect 4453 1078 4469 1112
rect 4537 1078 4553 1112
rect 4611 1078 4627 1112
rect 4695 1078 4711 1112
rect 4769 1078 4785 1112
rect 4853 1078 4869 1112
rect 4927 1078 4943 1112
rect 5011 1078 5027 1112
rect -5073 1019 -5039 1035
rect -5073 -1035 -5039 -1019
rect -4915 1019 -4881 1035
rect -4915 -1035 -4881 -1019
rect -4757 1019 -4723 1035
rect -4757 -1035 -4723 -1019
rect -4599 1019 -4565 1035
rect -4599 -1035 -4565 -1019
rect -4441 1019 -4407 1035
rect -4441 -1035 -4407 -1019
rect -4283 1019 -4249 1035
rect -4283 -1035 -4249 -1019
rect -4125 1019 -4091 1035
rect -4125 -1035 -4091 -1019
rect -3967 1019 -3933 1035
rect -3967 -1035 -3933 -1019
rect -3809 1019 -3775 1035
rect -3809 -1035 -3775 -1019
rect -3651 1019 -3617 1035
rect -3651 -1035 -3617 -1019
rect -3493 1019 -3459 1035
rect -3493 -1035 -3459 -1019
rect -3335 1019 -3301 1035
rect -3335 -1035 -3301 -1019
rect -3177 1019 -3143 1035
rect -3177 -1035 -3143 -1019
rect -3019 1019 -2985 1035
rect -3019 -1035 -2985 -1019
rect -2861 1019 -2827 1035
rect -2861 -1035 -2827 -1019
rect -2703 1019 -2669 1035
rect -2703 -1035 -2669 -1019
rect -2545 1019 -2511 1035
rect -2545 -1035 -2511 -1019
rect -2387 1019 -2353 1035
rect -2387 -1035 -2353 -1019
rect -2229 1019 -2195 1035
rect -2229 -1035 -2195 -1019
rect -2071 1019 -2037 1035
rect -2071 -1035 -2037 -1019
rect -1913 1019 -1879 1035
rect -1913 -1035 -1879 -1019
rect -1755 1019 -1721 1035
rect -1755 -1035 -1721 -1019
rect -1597 1019 -1563 1035
rect -1597 -1035 -1563 -1019
rect -1439 1019 -1405 1035
rect -1439 -1035 -1405 -1019
rect -1281 1019 -1247 1035
rect -1281 -1035 -1247 -1019
rect -1123 1019 -1089 1035
rect -1123 -1035 -1089 -1019
rect -965 1019 -931 1035
rect -965 -1035 -931 -1019
rect -807 1019 -773 1035
rect -807 -1035 -773 -1019
rect -649 1019 -615 1035
rect -649 -1035 -615 -1019
rect -491 1019 -457 1035
rect -491 -1035 -457 -1019
rect -333 1019 -299 1035
rect -333 -1035 -299 -1019
rect -175 1019 -141 1035
rect -175 -1035 -141 -1019
rect -17 1019 17 1035
rect -17 -1035 17 -1019
rect 141 1019 175 1035
rect 141 -1035 175 -1019
rect 299 1019 333 1035
rect 299 -1035 333 -1019
rect 457 1019 491 1035
rect 457 -1035 491 -1019
rect 615 1019 649 1035
rect 615 -1035 649 -1019
rect 773 1019 807 1035
rect 773 -1035 807 -1019
rect 931 1019 965 1035
rect 931 -1035 965 -1019
rect 1089 1019 1123 1035
rect 1089 -1035 1123 -1019
rect 1247 1019 1281 1035
rect 1247 -1035 1281 -1019
rect 1405 1019 1439 1035
rect 1405 -1035 1439 -1019
rect 1563 1019 1597 1035
rect 1563 -1035 1597 -1019
rect 1721 1019 1755 1035
rect 1721 -1035 1755 -1019
rect 1879 1019 1913 1035
rect 1879 -1035 1913 -1019
rect 2037 1019 2071 1035
rect 2037 -1035 2071 -1019
rect 2195 1019 2229 1035
rect 2195 -1035 2229 -1019
rect 2353 1019 2387 1035
rect 2353 -1035 2387 -1019
rect 2511 1019 2545 1035
rect 2511 -1035 2545 -1019
rect 2669 1019 2703 1035
rect 2669 -1035 2703 -1019
rect 2827 1019 2861 1035
rect 2827 -1035 2861 -1019
rect 2985 1019 3019 1035
rect 2985 -1035 3019 -1019
rect 3143 1019 3177 1035
rect 3143 -1035 3177 -1019
rect 3301 1019 3335 1035
rect 3301 -1035 3335 -1019
rect 3459 1019 3493 1035
rect 3459 -1035 3493 -1019
rect 3617 1019 3651 1035
rect 3617 -1035 3651 -1019
rect 3775 1019 3809 1035
rect 3775 -1035 3809 -1019
rect 3933 1019 3967 1035
rect 3933 -1035 3967 -1019
rect 4091 1019 4125 1035
rect 4091 -1035 4125 -1019
rect 4249 1019 4283 1035
rect 4249 -1035 4283 -1019
rect 4407 1019 4441 1035
rect 4407 -1035 4441 -1019
rect 4565 1019 4599 1035
rect 4565 -1035 4599 -1019
rect 4723 1019 4757 1035
rect 4723 -1035 4757 -1019
rect 4881 1019 4915 1035
rect 4881 -1035 4915 -1019
rect 5039 1019 5073 1035
rect 5039 -1035 5073 -1019
rect -5027 -1112 -5011 -1078
rect -4943 -1112 -4927 -1078
rect -4869 -1112 -4853 -1078
rect -4785 -1112 -4769 -1078
rect -4711 -1112 -4695 -1078
rect -4627 -1112 -4611 -1078
rect -4553 -1112 -4537 -1078
rect -4469 -1112 -4453 -1078
rect -4395 -1112 -4379 -1078
rect -4311 -1112 -4295 -1078
rect -4237 -1112 -4221 -1078
rect -4153 -1112 -4137 -1078
rect -4079 -1112 -4063 -1078
rect -3995 -1112 -3979 -1078
rect -3921 -1112 -3905 -1078
rect -3837 -1112 -3821 -1078
rect -3763 -1112 -3747 -1078
rect -3679 -1112 -3663 -1078
rect -3605 -1112 -3589 -1078
rect -3521 -1112 -3505 -1078
rect -3447 -1112 -3431 -1078
rect -3363 -1112 -3347 -1078
rect -3289 -1112 -3273 -1078
rect -3205 -1112 -3189 -1078
rect -3131 -1112 -3115 -1078
rect -3047 -1112 -3031 -1078
rect -2973 -1112 -2957 -1078
rect -2889 -1112 -2873 -1078
rect -2815 -1112 -2799 -1078
rect -2731 -1112 -2715 -1078
rect -2657 -1112 -2641 -1078
rect -2573 -1112 -2557 -1078
rect -2499 -1112 -2483 -1078
rect -2415 -1112 -2399 -1078
rect -2341 -1112 -2325 -1078
rect -2257 -1112 -2241 -1078
rect -2183 -1112 -2167 -1078
rect -2099 -1112 -2083 -1078
rect -2025 -1112 -2009 -1078
rect -1941 -1112 -1925 -1078
rect -1867 -1112 -1851 -1078
rect -1783 -1112 -1767 -1078
rect -1709 -1112 -1693 -1078
rect -1625 -1112 -1609 -1078
rect -1551 -1112 -1535 -1078
rect -1467 -1112 -1451 -1078
rect -1393 -1112 -1377 -1078
rect -1309 -1112 -1293 -1078
rect -1235 -1112 -1219 -1078
rect -1151 -1112 -1135 -1078
rect -1077 -1112 -1061 -1078
rect -993 -1112 -977 -1078
rect -919 -1112 -903 -1078
rect -835 -1112 -819 -1078
rect -761 -1112 -745 -1078
rect -677 -1112 -661 -1078
rect -603 -1112 -587 -1078
rect -519 -1112 -503 -1078
rect -445 -1112 -429 -1078
rect -361 -1112 -345 -1078
rect -287 -1112 -271 -1078
rect -203 -1112 -187 -1078
rect -129 -1112 -113 -1078
rect -45 -1112 -29 -1078
rect 29 -1112 45 -1078
rect 113 -1112 129 -1078
rect 187 -1112 203 -1078
rect 271 -1112 287 -1078
rect 345 -1112 361 -1078
rect 429 -1112 445 -1078
rect 503 -1112 519 -1078
rect 587 -1112 603 -1078
rect 661 -1112 677 -1078
rect 745 -1112 761 -1078
rect 819 -1112 835 -1078
rect 903 -1112 919 -1078
rect 977 -1112 993 -1078
rect 1061 -1112 1077 -1078
rect 1135 -1112 1151 -1078
rect 1219 -1112 1235 -1078
rect 1293 -1112 1309 -1078
rect 1377 -1112 1393 -1078
rect 1451 -1112 1467 -1078
rect 1535 -1112 1551 -1078
rect 1609 -1112 1625 -1078
rect 1693 -1112 1709 -1078
rect 1767 -1112 1783 -1078
rect 1851 -1112 1867 -1078
rect 1925 -1112 1941 -1078
rect 2009 -1112 2025 -1078
rect 2083 -1112 2099 -1078
rect 2167 -1112 2183 -1078
rect 2241 -1112 2257 -1078
rect 2325 -1112 2341 -1078
rect 2399 -1112 2415 -1078
rect 2483 -1112 2499 -1078
rect 2557 -1112 2573 -1078
rect 2641 -1112 2657 -1078
rect 2715 -1112 2731 -1078
rect 2799 -1112 2815 -1078
rect 2873 -1112 2889 -1078
rect 2957 -1112 2973 -1078
rect 3031 -1112 3047 -1078
rect 3115 -1112 3131 -1078
rect 3189 -1112 3205 -1078
rect 3273 -1112 3289 -1078
rect 3347 -1112 3363 -1078
rect 3431 -1112 3447 -1078
rect 3505 -1112 3521 -1078
rect 3589 -1112 3605 -1078
rect 3663 -1112 3679 -1078
rect 3747 -1112 3763 -1078
rect 3821 -1112 3837 -1078
rect 3905 -1112 3921 -1078
rect 3979 -1112 3995 -1078
rect 4063 -1112 4079 -1078
rect 4137 -1112 4153 -1078
rect 4221 -1112 4237 -1078
rect 4295 -1112 4311 -1078
rect 4379 -1112 4395 -1078
rect 4453 -1112 4469 -1078
rect 4537 -1112 4553 -1078
rect 4611 -1112 4627 -1078
rect 4695 -1112 4711 -1078
rect 4769 -1112 4785 -1078
rect 4853 -1112 4869 -1078
rect 4927 -1112 4943 -1078
rect 5011 -1112 5027 -1078
rect -5207 -1216 -5173 -1154
rect 5173 -1216 5207 -1154
rect -5207 -1250 -5111 -1216
rect 5111 -1250 5207 -1216
<< viali >>
rect -5011 1078 -4943 1112
rect -4853 1078 -4785 1112
rect -4695 1078 -4627 1112
rect -4537 1078 -4469 1112
rect -4379 1078 -4311 1112
rect -4221 1078 -4153 1112
rect -4063 1078 -3995 1112
rect -3905 1078 -3837 1112
rect -3747 1078 -3679 1112
rect -3589 1078 -3521 1112
rect -3431 1078 -3363 1112
rect -3273 1078 -3205 1112
rect -3115 1078 -3047 1112
rect -2957 1078 -2889 1112
rect -2799 1078 -2731 1112
rect -2641 1078 -2573 1112
rect -2483 1078 -2415 1112
rect -2325 1078 -2257 1112
rect -2167 1078 -2099 1112
rect -2009 1078 -1941 1112
rect -1851 1078 -1783 1112
rect -1693 1078 -1625 1112
rect -1535 1078 -1467 1112
rect -1377 1078 -1309 1112
rect -1219 1078 -1151 1112
rect -1061 1078 -993 1112
rect -903 1078 -835 1112
rect -745 1078 -677 1112
rect -587 1078 -519 1112
rect -429 1078 -361 1112
rect -271 1078 -203 1112
rect -113 1078 -45 1112
rect 45 1078 113 1112
rect 203 1078 271 1112
rect 361 1078 429 1112
rect 519 1078 587 1112
rect 677 1078 745 1112
rect 835 1078 903 1112
rect 993 1078 1061 1112
rect 1151 1078 1219 1112
rect 1309 1078 1377 1112
rect 1467 1078 1535 1112
rect 1625 1078 1693 1112
rect 1783 1078 1851 1112
rect 1941 1078 2009 1112
rect 2099 1078 2167 1112
rect 2257 1078 2325 1112
rect 2415 1078 2483 1112
rect 2573 1078 2641 1112
rect 2731 1078 2799 1112
rect 2889 1078 2957 1112
rect 3047 1078 3115 1112
rect 3205 1078 3273 1112
rect 3363 1078 3431 1112
rect 3521 1078 3589 1112
rect 3679 1078 3747 1112
rect 3837 1078 3905 1112
rect 3995 1078 4063 1112
rect 4153 1078 4221 1112
rect 4311 1078 4379 1112
rect 4469 1078 4537 1112
rect 4627 1078 4695 1112
rect 4785 1078 4853 1112
rect 4943 1078 5011 1112
rect -5073 -1019 -5039 1019
rect -4915 -1019 -4881 1019
rect -4757 -1019 -4723 1019
rect -4599 -1019 -4565 1019
rect -4441 -1019 -4407 1019
rect -4283 -1019 -4249 1019
rect -4125 -1019 -4091 1019
rect -3967 -1019 -3933 1019
rect -3809 -1019 -3775 1019
rect -3651 -1019 -3617 1019
rect -3493 -1019 -3459 1019
rect -3335 -1019 -3301 1019
rect -3177 -1019 -3143 1019
rect -3019 -1019 -2985 1019
rect -2861 -1019 -2827 1019
rect -2703 -1019 -2669 1019
rect -2545 -1019 -2511 1019
rect -2387 -1019 -2353 1019
rect -2229 -1019 -2195 1019
rect -2071 -1019 -2037 1019
rect -1913 -1019 -1879 1019
rect -1755 -1019 -1721 1019
rect -1597 -1019 -1563 1019
rect -1439 -1019 -1405 1019
rect -1281 -1019 -1247 1019
rect -1123 -1019 -1089 1019
rect -965 -1019 -931 1019
rect -807 -1019 -773 1019
rect -649 -1019 -615 1019
rect -491 -1019 -457 1019
rect -333 -1019 -299 1019
rect -175 -1019 -141 1019
rect -17 -1019 17 1019
rect 141 -1019 175 1019
rect 299 -1019 333 1019
rect 457 -1019 491 1019
rect 615 -1019 649 1019
rect 773 -1019 807 1019
rect 931 -1019 965 1019
rect 1089 -1019 1123 1019
rect 1247 -1019 1281 1019
rect 1405 -1019 1439 1019
rect 1563 -1019 1597 1019
rect 1721 -1019 1755 1019
rect 1879 -1019 1913 1019
rect 2037 -1019 2071 1019
rect 2195 -1019 2229 1019
rect 2353 -1019 2387 1019
rect 2511 -1019 2545 1019
rect 2669 -1019 2703 1019
rect 2827 -1019 2861 1019
rect 2985 -1019 3019 1019
rect 3143 -1019 3177 1019
rect 3301 -1019 3335 1019
rect 3459 -1019 3493 1019
rect 3617 -1019 3651 1019
rect 3775 -1019 3809 1019
rect 3933 -1019 3967 1019
rect 4091 -1019 4125 1019
rect 4249 -1019 4283 1019
rect 4407 -1019 4441 1019
rect 4565 -1019 4599 1019
rect 4723 -1019 4757 1019
rect 4881 -1019 4915 1019
rect 5039 -1019 5073 1019
rect -5011 -1112 -4943 -1078
rect -4853 -1112 -4785 -1078
rect -4695 -1112 -4627 -1078
rect -4537 -1112 -4469 -1078
rect -4379 -1112 -4311 -1078
rect -4221 -1112 -4153 -1078
rect -4063 -1112 -3995 -1078
rect -3905 -1112 -3837 -1078
rect -3747 -1112 -3679 -1078
rect -3589 -1112 -3521 -1078
rect -3431 -1112 -3363 -1078
rect -3273 -1112 -3205 -1078
rect -3115 -1112 -3047 -1078
rect -2957 -1112 -2889 -1078
rect -2799 -1112 -2731 -1078
rect -2641 -1112 -2573 -1078
rect -2483 -1112 -2415 -1078
rect -2325 -1112 -2257 -1078
rect -2167 -1112 -2099 -1078
rect -2009 -1112 -1941 -1078
rect -1851 -1112 -1783 -1078
rect -1693 -1112 -1625 -1078
rect -1535 -1112 -1467 -1078
rect -1377 -1112 -1309 -1078
rect -1219 -1112 -1151 -1078
rect -1061 -1112 -993 -1078
rect -903 -1112 -835 -1078
rect -745 -1112 -677 -1078
rect -587 -1112 -519 -1078
rect -429 -1112 -361 -1078
rect -271 -1112 -203 -1078
rect -113 -1112 -45 -1078
rect 45 -1112 113 -1078
rect 203 -1112 271 -1078
rect 361 -1112 429 -1078
rect 519 -1112 587 -1078
rect 677 -1112 745 -1078
rect 835 -1112 903 -1078
rect 993 -1112 1061 -1078
rect 1151 -1112 1219 -1078
rect 1309 -1112 1377 -1078
rect 1467 -1112 1535 -1078
rect 1625 -1112 1693 -1078
rect 1783 -1112 1851 -1078
rect 1941 -1112 2009 -1078
rect 2099 -1112 2167 -1078
rect 2257 -1112 2325 -1078
rect 2415 -1112 2483 -1078
rect 2573 -1112 2641 -1078
rect 2731 -1112 2799 -1078
rect 2889 -1112 2957 -1078
rect 3047 -1112 3115 -1078
rect 3205 -1112 3273 -1078
rect 3363 -1112 3431 -1078
rect 3521 -1112 3589 -1078
rect 3679 -1112 3747 -1078
rect 3837 -1112 3905 -1078
rect 3995 -1112 4063 -1078
rect 4153 -1112 4221 -1078
rect 4311 -1112 4379 -1078
rect 4469 -1112 4537 -1078
rect 4627 -1112 4695 -1078
rect 4785 -1112 4853 -1078
rect 4943 -1112 5011 -1078
<< metal1 >>
rect -5023 1112 -4931 1118
rect -5023 1078 -5011 1112
rect -4943 1078 -4931 1112
rect -5023 1072 -4931 1078
rect -4865 1112 -4773 1118
rect -4865 1078 -4853 1112
rect -4785 1078 -4773 1112
rect -4865 1072 -4773 1078
rect -4707 1112 -4615 1118
rect -4707 1078 -4695 1112
rect -4627 1078 -4615 1112
rect -4707 1072 -4615 1078
rect -4549 1112 -4457 1118
rect -4549 1078 -4537 1112
rect -4469 1078 -4457 1112
rect -4549 1072 -4457 1078
rect -4391 1112 -4299 1118
rect -4391 1078 -4379 1112
rect -4311 1078 -4299 1112
rect -4391 1072 -4299 1078
rect -4233 1112 -4141 1118
rect -4233 1078 -4221 1112
rect -4153 1078 -4141 1112
rect -4233 1072 -4141 1078
rect -4075 1112 -3983 1118
rect -4075 1078 -4063 1112
rect -3995 1078 -3983 1112
rect -4075 1072 -3983 1078
rect -3917 1112 -3825 1118
rect -3917 1078 -3905 1112
rect -3837 1078 -3825 1112
rect -3917 1072 -3825 1078
rect -3759 1112 -3667 1118
rect -3759 1078 -3747 1112
rect -3679 1078 -3667 1112
rect -3759 1072 -3667 1078
rect -3601 1112 -3509 1118
rect -3601 1078 -3589 1112
rect -3521 1078 -3509 1112
rect -3601 1072 -3509 1078
rect -3443 1112 -3351 1118
rect -3443 1078 -3431 1112
rect -3363 1078 -3351 1112
rect -3443 1072 -3351 1078
rect -3285 1112 -3193 1118
rect -3285 1078 -3273 1112
rect -3205 1078 -3193 1112
rect -3285 1072 -3193 1078
rect -3127 1112 -3035 1118
rect -3127 1078 -3115 1112
rect -3047 1078 -3035 1112
rect -3127 1072 -3035 1078
rect -2969 1112 -2877 1118
rect -2969 1078 -2957 1112
rect -2889 1078 -2877 1112
rect -2969 1072 -2877 1078
rect -2811 1112 -2719 1118
rect -2811 1078 -2799 1112
rect -2731 1078 -2719 1112
rect -2811 1072 -2719 1078
rect -2653 1112 -2561 1118
rect -2653 1078 -2641 1112
rect -2573 1078 -2561 1112
rect -2653 1072 -2561 1078
rect -2495 1112 -2403 1118
rect -2495 1078 -2483 1112
rect -2415 1078 -2403 1112
rect -2495 1072 -2403 1078
rect -2337 1112 -2245 1118
rect -2337 1078 -2325 1112
rect -2257 1078 -2245 1112
rect -2337 1072 -2245 1078
rect -2179 1112 -2087 1118
rect -2179 1078 -2167 1112
rect -2099 1078 -2087 1112
rect -2179 1072 -2087 1078
rect -2021 1112 -1929 1118
rect -2021 1078 -2009 1112
rect -1941 1078 -1929 1112
rect -2021 1072 -1929 1078
rect -1863 1112 -1771 1118
rect -1863 1078 -1851 1112
rect -1783 1078 -1771 1112
rect -1863 1072 -1771 1078
rect -1705 1112 -1613 1118
rect -1705 1078 -1693 1112
rect -1625 1078 -1613 1112
rect -1705 1072 -1613 1078
rect -1547 1112 -1455 1118
rect -1547 1078 -1535 1112
rect -1467 1078 -1455 1112
rect -1547 1072 -1455 1078
rect -1389 1112 -1297 1118
rect -1389 1078 -1377 1112
rect -1309 1078 -1297 1112
rect -1389 1072 -1297 1078
rect -1231 1112 -1139 1118
rect -1231 1078 -1219 1112
rect -1151 1078 -1139 1112
rect -1231 1072 -1139 1078
rect -1073 1112 -981 1118
rect -1073 1078 -1061 1112
rect -993 1078 -981 1112
rect -1073 1072 -981 1078
rect -915 1112 -823 1118
rect -915 1078 -903 1112
rect -835 1078 -823 1112
rect -915 1072 -823 1078
rect -757 1112 -665 1118
rect -757 1078 -745 1112
rect -677 1078 -665 1112
rect -757 1072 -665 1078
rect -599 1112 -507 1118
rect -599 1078 -587 1112
rect -519 1078 -507 1112
rect -599 1072 -507 1078
rect -441 1112 -349 1118
rect -441 1078 -429 1112
rect -361 1078 -349 1112
rect -441 1072 -349 1078
rect -283 1112 -191 1118
rect -283 1078 -271 1112
rect -203 1078 -191 1112
rect -283 1072 -191 1078
rect -125 1112 -33 1118
rect -125 1078 -113 1112
rect -45 1078 -33 1112
rect -125 1072 -33 1078
rect 33 1112 125 1118
rect 33 1078 45 1112
rect 113 1078 125 1112
rect 33 1072 125 1078
rect 191 1112 283 1118
rect 191 1078 203 1112
rect 271 1078 283 1112
rect 191 1072 283 1078
rect 349 1112 441 1118
rect 349 1078 361 1112
rect 429 1078 441 1112
rect 349 1072 441 1078
rect 507 1112 599 1118
rect 507 1078 519 1112
rect 587 1078 599 1112
rect 507 1072 599 1078
rect 665 1112 757 1118
rect 665 1078 677 1112
rect 745 1078 757 1112
rect 665 1072 757 1078
rect 823 1112 915 1118
rect 823 1078 835 1112
rect 903 1078 915 1112
rect 823 1072 915 1078
rect 981 1112 1073 1118
rect 981 1078 993 1112
rect 1061 1078 1073 1112
rect 981 1072 1073 1078
rect 1139 1112 1231 1118
rect 1139 1078 1151 1112
rect 1219 1078 1231 1112
rect 1139 1072 1231 1078
rect 1297 1112 1389 1118
rect 1297 1078 1309 1112
rect 1377 1078 1389 1112
rect 1297 1072 1389 1078
rect 1455 1112 1547 1118
rect 1455 1078 1467 1112
rect 1535 1078 1547 1112
rect 1455 1072 1547 1078
rect 1613 1112 1705 1118
rect 1613 1078 1625 1112
rect 1693 1078 1705 1112
rect 1613 1072 1705 1078
rect 1771 1112 1863 1118
rect 1771 1078 1783 1112
rect 1851 1078 1863 1112
rect 1771 1072 1863 1078
rect 1929 1112 2021 1118
rect 1929 1078 1941 1112
rect 2009 1078 2021 1112
rect 1929 1072 2021 1078
rect 2087 1112 2179 1118
rect 2087 1078 2099 1112
rect 2167 1078 2179 1112
rect 2087 1072 2179 1078
rect 2245 1112 2337 1118
rect 2245 1078 2257 1112
rect 2325 1078 2337 1112
rect 2245 1072 2337 1078
rect 2403 1112 2495 1118
rect 2403 1078 2415 1112
rect 2483 1078 2495 1112
rect 2403 1072 2495 1078
rect 2561 1112 2653 1118
rect 2561 1078 2573 1112
rect 2641 1078 2653 1112
rect 2561 1072 2653 1078
rect 2719 1112 2811 1118
rect 2719 1078 2731 1112
rect 2799 1078 2811 1112
rect 2719 1072 2811 1078
rect 2877 1112 2969 1118
rect 2877 1078 2889 1112
rect 2957 1078 2969 1112
rect 2877 1072 2969 1078
rect 3035 1112 3127 1118
rect 3035 1078 3047 1112
rect 3115 1078 3127 1112
rect 3035 1072 3127 1078
rect 3193 1112 3285 1118
rect 3193 1078 3205 1112
rect 3273 1078 3285 1112
rect 3193 1072 3285 1078
rect 3351 1112 3443 1118
rect 3351 1078 3363 1112
rect 3431 1078 3443 1112
rect 3351 1072 3443 1078
rect 3509 1112 3601 1118
rect 3509 1078 3521 1112
rect 3589 1078 3601 1112
rect 3509 1072 3601 1078
rect 3667 1112 3759 1118
rect 3667 1078 3679 1112
rect 3747 1078 3759 1112
rect 3667 1072 3759 1078
rect 3825 1112 3917 1118
rect 3825 1078 3837 1112
rect 3905 1078 3917 1112
rect 3825 1072 3917 1078
rect 3983 1112 4075 1118
rect 3983 1078 3995 1112
rect 4063 1078 4075 1112
rect 3983 1072 4075 1078
rect 4141 1112 4233 1118
rect 4141 1078 4153 1112
rect 4221 1078 4233 1112
rect 4141 1072 4233 1078
rect 4299 1112 4391 1118
rect 4299 1078 4311 1112
rect 4379 1078 4391 1112
rect 4299 1072 4391 1078
rect 4457 1112 4549 1118
rect 4457 1078 4469 1112
rect 4537 1078 4549 1112
rect 4457 1072 4549 1078
rect 4615 1112 4707 1118
rect 4615 1078 4627 1112
rect 4695 1078 4707 1112
rect 4615 1072 4707 1078
rect 4773 1112 4865 1118
rect 4773 1078 4785 1112
rect 4853 1078 4865 1112
rect 4773 1072 4865 1078
rect 4931 1112 5023 1118
rect 4931 1078 4943 1112
rect 5011 1078 5023 1112
rect 4931 1072 5023 1078
rect -5079 1019 -5033 1031
rect -5079 -1019 -5073 1019
rect -5039 -1019 -5033 1019
rect -5079 -1031 -5033 -1019
rect -4921 1019 -4875 1031
rect -4921 -1019 -4915 1019
rect -4881 -1019 -4875 1019
rect -4921 -1031 -4875 -1019
rect -4763 1019 -4717 1031
rect -4763 -1019 -4757 1019
rect -4723 -1019 -4717 1019
rect -4763 -1031 -4717 -1019
rect -4605 1019 -4559 1031
rect -4605 -1019 -4599 1019
rect -4565 -1019 -4559 1019
rect -4605 -1031 -4559 -1019
rect -4447 1019 -4401 1031
rect -4447 -1019 -4441 1019
rect -4407 -1019 -4401 1019
rect -4447 -1031 -4401 -1019
rect -4289 1019 -4243 1031
rect -4289 -1019 -4283 1019
rect -4249 -1019 -4243 1019
rect -4289 -1031 -4243 -1019
rect -4131 1019 -4085 1031
rect -4131 -1019 -4125 1019
rect -4091 -1019 -4085 1019
rect -4131 -1031 -4085 -1019
rect -3973 1019 -3927 1031
rect -3973 -1019 -3967 1019
rect -3933 -1019 -3927 1019
rect -3973 -1031 -3927 -1019
rect -3815 1019 -3769 1031
rect -3815 -1019 -3809 1019
rect -3775 -1019 -3769 1019
rect -3815 -1031 -3769 -1019
rect -3657 1019 -3611 1031
rect -3657 -1019 -3651 1019
rect -3617 -1019 -3611 1019
rect -3657 -1031 -3611 -1019
rect -3499 1019 -3453 1031
rect -3499 -1019 -3493 1019
rect -3459 -1019 -3453 1019
rect -3499 -1031 -3453 -1019
rect -3341 1019 -3295 1031
rect -3341 -1019 -3335 1019
rect -3301 -1019 -3295 1019
rect -3341 -1031 -3295 -1019
rect -3183 1019 -3137 1031
rect -3183 -1019 -3177 1019
rect -3143 -1019 -3137 1019
rect -3183 -1031 -3137 -1019
rect -3025 1019 -2979 1031
rect -3025 -1019 -3019 1019
rect -2985 -1019 -2979 1019
rect -3025 -1031 -2979 -1019
rect -2867 1019 -2821 1031
rect -2867 -1019 -2861 1019
rect -2827 -1019 -2821 1019
rect -2867 -1031 -2821 -1019
rect -2709 1019 -2663 1031
rect -2709 -1019 -2703 1019
rect -2669 -1019 -2663 1019
rect -2709 -1031 -2663 -1019
rect -2551 1019 -2505 1031
rect -2551 -1019 -2545 1019
rect -2511 -1019 -2505 1019
rect -2551 -1031 -2505 -1019
rect -2393 1019 -2347 1031
rect -2393 -1019 -2387 1019
rect -2353 -1019 -2347 1019
rect -2393 -1031 -2347 -1019
rect -2235 1019 -2189 1031
rect -2235 -1019 -2229 1019
rect -2195 -1019 -2189 1019
rect -2235 -1031 -2189 -1019
rect -2077 1019 -2031 1031
rect -2077 -1019 -2071 1019
rect -2037 -1019 -2031 1019
rect -2077 -1031 -2031 -1019
rect -1919 1019 -1873 1031
rect -1919 -1019 -1913 1019
rect -1879 -1019 -1873 1019
rect -1919 -1031 -1873 -1019
rect -1761 1019 -1715 1031
rect -1761 -1019 -1755 1019
rect -1721 -1019 -1715 1019
rect -1761 -1031 -1715 -1019
rect -1603 1019 -1557 1031
rect -1603 -1019 -1597 1019
rect -1563 -1019 -1557 1019
rect -1603 -1031 -1557 -1019
rect -1445 1019 -1399 1031
rect -1445 -1019 -1439 1019
rect -1405 -1019 -1399 1019
rect -1445 -1031 -1399 -1019
rect -1287 1019 -1241 1031
rect -1287 -1019 -1281 1019
rect -1247 -1019 -1241 1019
rect -1287 -1031 -1241 -1019
rect -1129 1019 -1083 1031
rect -1129 -1019 -1123 1019
rect -1089 -1019 -1083 1019
rect -1129 -1031 -1083 -1019
rect -971 1019 -925 1031
rect -971 -1019 -965 1019
rect -931 -1019 -925 1019
rect -971 -1031 -925 -1019
rect -813 1019 -767 1031
rect -813 -1019 -807 1019
rect -773 -1019 -767 1019
rect -813 -1031 -767 -1019
rect -655 1019 -609 1031
rect -655 -1019 -649 1019
rect -615 -1019 -609 1019
rect -655 -1031 -609 -1019
rect -497 1019 -451 1031
rect -497 -1019 -491 1019
rect -457 -1019 -451 1019
rect -497 -1031 -451 -1019
rect -339 1019 -293 1031
rect -339 -1019 -333 1019
rect -299 -1019 -293 1019
rect -339 -1031 -293 -1019
rect -181 1019 -135 1031
rect -181 -1019 -175 1019
rect -141 -1019 -135 1019
rect -181 -1031 -135 -1019
rect -23 1019 23 1031
rect -23 -1019 -17 1019
rect 17 -1019 23 1019
rect -23 -1031 23 -1019
rect 135 1019 181 1031
rect 135 -1019 141 1019
rect 175 -1019 181 1019
rect 135 -1031 181 -1019
rect 293 1019 339 1031
rect 293 -1019 299 1019
rect 333 -1019 339 1019
rect 293 -1031 339 -1019
rect 451 1019 497 1031
rect 451 -1019 457 1019
rect 491 -1019 497 1019
rect 451 -1031 497 -1019
rect 609 1019 655 1031
rect 609 -1019 615 1019
rect 649 -1019 655 1019
rect 609 -1031 655 -1019
rect 767 1019 813 1031
rect 767 -1019 773 1019
rect 807 -1019 813 1019
rect 767 -1031 813 -1019
rect 925 1019 971 1031
rect 925 -1019 931 1019
rect 965 -1019 971 1019
rect 925 -1031 971 -1019
rect 1083 1019 1129 1031
rect 1083 -1019 1089 1019
rect 1123 -1019 1129 1019
rect 1083 -1031 1129 -1019
rect 1241 1019 1287 1031
rect 1241 -1019 1247 1019
rect 1281 -1019 1287 1019
rect 1241 -1031 1287 -1019
rect 1399 1019 1445 1031
rect 1399 -1019 1405 1019
rect 1439 -1019 1445 1019
rect 1399 -1031 1445 -1019
rect 1557 1019 1603 1031
rect 1557 -1019 1563 1019
rect 1597 -1019 1603 1019
rect 1557 -1031 1603 -1019
rect 1715 1019 1761 1031
rect 1715 -1019 1721 1019
rect 1755 -1019 1761 1019
rect 1715 -1031 1761 -1019
rect 1873 1019 1919 1031
rect 1873 -1019 1879 1019
rect 1913 -1019 1919 1019
rect 1873 -1031 1919 -1019
rect 2031 1019 2077 1031
rect 2031 -1019 2037 1019
rect 2071 -1019 2077 1019
rect 2031 -1031 2077 -1019
rect 2189 1019 2235 1031
rect 2189 -1019 2195 1019
rect 2229 -1019 2235 1019
rect 2189 -1031 2235 -1019
rect 2347 1019 2393 1031
rect 2347 -1019 2353 1019
rect 2387 -1019 2393 1019
rect 2347 -1031 2393 -1019
rect 2505 1019 2551 1031
rect 2505 -1019 2511 1019
rect 2545 -1019 2551 1019
rect 2505 -1031 2551 -1019
rect 2663 1019 2709 1031
rect 2663 -1019 2669 1019
rect 2703 -1019 2709 1019
rect 2663 -1031 2709 -1019
rect 2821 1019 2867 1031
rect 2821 -1019 2827 1019
rect 2861 -1019 2867 1019
rect 2821 -1031 2867 -1019
rect 2979 1019 3025 1031
rect 2979 -1019 2985 1019
rect 3019 -1019 3025 1019
rect 2979 -1031 3025 -1019
rect 3137 1019 3183 1031
rect 3137 -1019 3143 1019
rect 3177 -1019 3183 1019
rect 3137 -1031 3183 -1019
rect 3295 1019 3341 1031
rect 3295 -1019 3301 1019
rect 3335 -1019 3341 1019
rect 3295 -1031 3341 -1019
rect 3453 1019 3499 1031
rect 3453 -1019 3459 1019
rect 3493 -1019 3499 1019
rect 3453 -1031 3499 -1019
rect 3611 1019 3657 1031
rect 3611 -1019 3617 1019
rect 3651 -1019 3657 1019
rect 3611 -1031 3657 -1019
rect 3769 1019 3815 1031
rect 3769 -1019 3775 1019
rect 3809 -1019 3815 1019
rect 3769 -1031 3815 -1019
rect 3927 1019 3973 1031
rect 3927 -1019 3933 1019
rect 3967 -1019 3973 1019
rect 3927 -1031 3973 -1019
rect 4085 1019 4131 1031
rect 4085 -1019 4091 1019
rect 4125 -1019 4131 1019
rect 4085 -1031 4131 -1019
rect 4243 1019 4289 1031
rect 4243 -1019 4249 1019
rect 4283 -1019 4289 1019
rect 4243 -1031 4289 -1019
rect 4401 1019 4447 1031
rect 4401 -1019 4407 1019
rect 4441 -1019 4447 1019
rect 4401 -1031 4447 -1019
rect 4559 1019 4605 1031
rect 4559 -1019 4565 1019
rect 4599 -1019 4605 1019
rect 4559 -1031 4605 -1019
rect 4717 1019 4763 1031
rect 4717 -1019 4723 1019
rect 4757 -1019 4763 1019
rect 4717 -1031 4763 -1019
rect 4875 1019 4921 1031
rect 4875 -1019 4881 1019
rect 4915 -1019 4921 1019
rect 4875 -1031 4921 -1019
rect 5033 1019 5079 1031
rect 5033 -1019 5039 1019
rect 5073 -1019 5079 1019
rect 5033 -1031 5079 -1019
rect -5023 -1078 -4931 -1072
rect -5023 -1112 -5011 -1078
rect -4943 -1112 -4931 -1078
rect -5023 -1118 -4931 -1112
rect -4865 -1078 -4773 -1072
rect -4865 -1112 -4853 -1078
rect -4785 -1112 -4773 -1078
rect -4865 -1118 -4773 -1112
rect -4707 -1078 -4615 -1072
rect -4707 -1112 -4695 -1078
rect -4627 -1112 -4615 -1078
rect -4707 -1118 -4615 -1112
rect -4549 -1078 -4457 -1072
rect -4549 -1112 -4537 -1078
rect -4469 -1112 -4457 -1078
rect -4549 -1118 -4457 -1112
rect -4391 -1078 -4299 -1072
rect -4391 -1112 -4379 -1078
rect -4311 -1112 -4299 -1078
rect -4391 -1118 -4299 -1112
rect -4233 -1078 -4141 -1072
rect -4233 -1112 -4221 -1078
rect -4153 -1112 -4141 -1078
rect -4233 -1118 -4141 -1112
rect -4075 -1078 -3983 -1072
rect -4075 -1112 -4063 -1078
rect -3995 -1112 -3983 -1078
rect -4075 -1118 -3983 -1112
rect -3917 -1078 -3825 -1072
rect -3917 -1112 -3905 -1078
rect -3837 -1112 -3825 -1078
rect -3917 -1118 -3825 -1112
rect -3759 -1078 -3667 -1072
rect -3759 -1112 -3747 -1078
rect -3679 -1112 -3667 -1078
rect -3759 -1118 -3667 -1112
rect -3601 -1078 -3509 -1072
rect -3601 -1112 -3589 -1078
rect -3521 -1112 -3509 -1078
rect -3601 -1118 -3509 -1112
rect -3443 -1078 -3351 -1072
rect -3443 -1112 -3431 -1078
rect -3363 -1112 -3351 -1078
rect -3443 -1118 -3351 -1112
rect -3285 -1078 -3193 -1072
rect -3285 -1112 -3273 -1078
rect -3205 -1112 -3193 -1078
rect -3285 -1118 -3193 -1112
rect -3127 -1078 -3035 -1072
rect -3127 -1112 -3115 -1078
rect -3047 -1112 -3035 -1078
rect -3127 -1118 -3035 -1112
rect -2969 -1078 -2877 -1072
rect -2969 -1112 -2957 -1078
rect -2889 -1112 -2877 -1078
rect -2969 -1118 -2877 -1112
rect -2811 -1078 -2719 -1072
rect -2811 -1112 -2799 -1078
rect -2731 -1112 -2719 -1078
rect -2811 -1118 -2719 -1112
rect -2653 -1078 -2561 -1072
rect -2653 -1112 -2641 -1078
rect -2573 -1112 -2561 -1078
rect -2653 -1118 -2561 -1112
rect -2495 -1078 -2403 -1072
rect -2495 -1112 -2483 -1078
rect -2415 -1112 -2403 -1078
rect -2495 -1118 -2403 -1112
rect -2337 -1078 -2245 -1072
rect -2337 -1112 -2325 -1078
rect -2257 -1112 -2245 -1078
rect -2337 -1118 -2245 -1112
rect -2179 -1078 -2087 -1072
rect -2179 -1112 -2167 -1078
rect -2099 -1112 -2087 -1078
rect -2179 -1118 -2087 -1112
rect -2021 -1078 -1929 -1072
rect -2021 -1112 -2009 -1078
rect -1941 -1112 -1929 -1078
rect -2021 -1118 -1929 -1112
rect -1863 -1078 -1771 -1072
rect -1863 -1112 -1851 -1078
rect -1783 -1112 -1771 -1078
rect -1863 -1118 -1771 -1112
rect -1705 -1078 -1613 -1072
rect -1705 -1112 -1693 -1078
rect -1625 -1112 -1613 -1078
rect -1705 -1118 -1613 -1112
rect -1547 -1078 -1455 -1072
rect -1547 -1112 -1535 -1078
rect -1467 -1112 -1455 -1078
rect -1547 -1118 -1455 -1112
rect -1389 -1078 -1297 -1072
rect -1389 -1112 -1377 -1078
rect -1309 -1112 -1297 -1078
rect -1389 -1118 -1297 -1112
rect -1231 -1078 -1139 -1072
rect -1231 -1112 -1219 -1078
rect -1151 -1112 -1139 -1078
rect -1231 -1118 -1139 -1112
rect -1073 -1078 -981 -1072
rect -1073 -1112 -1061 -1078
rect -993 -1112 -981 -1078
rect -1073 -1118 -981 -1112
rect -915 -1078 -823 -1072
rect -915 -1112 -903 -1078
rect -835 -1112 -823 -1078
rect -915 -1118 -823 -1112
rect -757 -1078 -665 -1072
rect -757 -1112 -745 -1078
rect -677 -1112 -665 -1078
rect -757 -1118 -665 -1112
rect -599 -1078 -507 -1072
rect -599 -1112 -587 -1078
rect -519 -1112 -507 -1078
rect -599 -1118 -507 -1112
rect -441 -1078 -349 -1072
rect -441 -1112 -429 -1078
rect -361 -1112 -349 -1078
rect -441 -1118 -349 -1112
rect -283 -1078 -191 -1072
rect -283 -1112 -271 -1078
rect -203 -1112 -191 -1078
rect -283 -1118 -191 -1112
rect -125 -1078 -33 -1072
rect -125 -1112 -113 -1078
rect -45 -1112 -33 -1078
rect -125 -1118 -33 -1112
rect 33 -1078 125 -1072
rect 33 -1112 45 -1078
rect 113 -1112 125 -1078
rect 33 -1118 125 -1112
rect 191 -1078 283 -1072
rect 191 -1112 203 -1078
rect 271 -1112 283 -1078
rect 191 -1118 283 -1112
rect 349 -1078 441 -1072
rect 349 -1112 361 -1078
rect 429 -1112 441 -1078
rect 349 -1118 441 -1112
rect 507 -1078 599 -1072
rect 507 -1112 519 -1078
rect 587 -1112 599 -1078
rect 507 -1118 599 -1112
rect 665 -1078 757 -1072
rect 665 -1112 677 -1078
rect 745 -1112 757 -1078
rect 665 -1118 757 -1112
rect 823 -1078 915 -1072
rect 823 -1112 835 -1078
rect 903 -1112 915 -1078
rect 823 -1118 915 -1112
rect 981 -1078 1073 -1072
rect 981 -1112 993 -1078
rect 1061 -1112 1073 -1078
rect 981 -1118 1073 -1112
rect 1139 -1078 1231 -1072
rect 1139 -1112 1151 -1078
rect 1219 -1112 1231 -1078
rect 1139 -1118 1231 -1112
rect 1297 -1078 1389 -1072
rect 1297 -1112 1309 -1078
rect 1377 -1112 1389 -1078
rect 1297 -1118 1389 -1112
rect 1455 -1078 1547 -1072
rect 1455 -1112 1467 -1078
rect 1535 -1112 1547 -1078
rect 1455 -1118 1547 -1112
rect 1613 -1078 1705 -1072
rect 1613 -1112 1625 -1078
rect 1693 -1112 1705 -1078
rect 1613 -1118 1705 -1112
rect 1771 -1078 1863 -1072
rect 1771 -1112 1783 -1078
rect 1851 -1112 1863 -1078
rect 1771 -1118 1863 -1112
rect 1929 -1078 2021 -1072
rect 1929 -1112 1941 -1078
rect 2009 -1112 2021 -1078
rect 1929 -1118 2021 -1112
rect 2087 -1078 2179 -1072
rect 2087 -1112 2099 -1078
rect 2167 -1112 2179 -1078
rect 2087 -1118 2179 -1112
rect 2245 -1078 2337 -1072
rect 2245 -1112 2257 -1078
rect 2325 -1112 2337 -1078
rect 2245 -1118 2337 -1112
rect 2403 -1078 2495 -1072
rect 2403 -1112 2415 -1078
rect 2483 -1112 2495 -1078
rect 2403 -1118 2495 -1112
rect 2561 -1078 2653 -1072
rect 2561 -1112 2573 -1078
rect 2641 -1112 2653 -1078
rect 2561 -1118 2653 -1112
rect 2719 -1078 2811 -1072
rect 2719 -1112 2731 -1078
rect 2799 -1112 2811 -1078
rect 2719 -1118 2811 -1112
rect 2877 -1078 2969 -1072
rect 2877 -1112 2889 -1078
rect 2957 -1112 2969 -1078
rect 2877 -1118 2969 -1112
rect 3035 -1078 3127 -1072
rect 3035 -1112 3047 -1078
rect 3115 -1112 3127 -1078
rect 3035 -1118 3127 -1112
rect 3193 -1078 3285 -1072
rect 3193 -1112 3205 -1078
rect 3273 -1112 3285 -1078
rect 3193 -1118 3285 -1112
rect 3351 -1078 3443 -1072
rect 3351 -1112 3363 -1078
rect 3431 -1112 3443 -1078
rect 3351 -1118 3443 -1112
rect 3509 -1078 3601 -1072
rect 3509 -1112 3521 -1078
rect 3589 -1112 3601 -1078
rect 3509 -1118 3601 -1112
rect 3667 -1078 3759 -1072
rect 3667 -1112 3679 -1078
rect 3747 -1112 3759 -1078
rect 3667 -1118 3759 -1112
rect 3825 -1078 3917 -1072
rect 3825 -1112 3837 -1078
rect 3905 -1112 3917 -1078
rect 3825 -1118 3917 -1112
rect 3983 -1078 4075 -1072
rect 3983 -1112 3995 -1078
rect 4063 -1112 4075 -1078
rect 3983 -1118 4075 -1112
rect 4141 -1078 4233 -1072
rect 4141 -1112 4153 -1078
rect 4221 -1112 4233 -1078
rect 4141 -1118 4233 -1112
rect 4299 -1078 4391 -1072
rect 4299 -1112 4311 -1078
rect 4379 -1112 4391 -1078
rect 4299 -1118 4391 -1112
rect 4457 -1078 4549 -1072
rect 4457 -1112 4469 -1078
rect 4537 -1112 4549 -1078
rect 4457 -1118 4549 -1112
rect 4615 -1078 4707 -1072
rect 4615 -1112 4627 -1078
rect 4695 -1112 4707 -1078
rect 4615 -1118 4707 -1112
rect 4773 -1078 4865 -1072
rect 4773 -1112 4785 -1078
rect 4853 -1112 4865 -1078
rect 4773 -1118 4865 -1112
rect 4931 -1078 5023 -1072
rect 4931 -1112 4943 -1078
rect 5011 -1112 5023 -1078
rect 4931 -1118 5023 -1112
<< properties >>
string FIXED_BBOX -5190 -1233 5190 1233
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.3125 l 0.5 m 1 nf 64 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
