magic
tech sky130A
magscale 1 2
timestamp 1770370310
<< pwell >>
rect -201 -2932 201 2932
<< psubdiff >>
rect -165 2862 -69 2896
rect 69 2862 165 2896
rect -165 2800 -131 2862
rect 131 2800 165 2862
rect -165 -2862 -131 -2800
rect 131 -2862 165 -2800
rect -165 -2896 -69 -2862
rect 69 -2896 165 -2862
<< psubdiffcont >>
rect -69 2862 69 2896
rect -165 -2800 -131 2800
rect 131 -2800 165 2800
rect -69 -2896 69 -2862
<< xpolycontact >>
rect -35 2334 35 2766
rect -35 -2766 35 -2334
<< ppolyres >>
rect -35 -2334 35 2334
<< locali >>
rect -165 2862 -69 2896
rect 69 2862 165 2896
rect -165 2800 -131 2862
rect 131 2800 165 2862
rect -165 -2862 -131 -2800
rect 131 -2862 165 -2800
rect -165 -2896 -69 -2862
rect 69 -2896 165 -2862
<< viali >>
rect -19 2351 19 2748
rect -19 -2748 19 -2351
<< metal1 >>
rect -25 2748 25 2760
rect -25 2351 -19 2748
rect 19 2351 25 2748
rect -25 2339 25 2351
rect -25 -2351 25 -2339
rect -25 -2748 -19 -2351
rect 19 -2748 25 -2351
rect -25 -2760 25 -2748
<< properties >>
string FIXED_BBOX -148 -2879 148 2879
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 23.5 m 1 nx 1 wmin 0.350 lmin 0.50 class resistor rho 319.8 val 22.585k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0 mult 1
<< end >>
