magic
tech sky130A
magscale 1 2
timestamp 1770112220
<< metal3 >>
rect -22328 21132 -16956 21160
rect -22328 16108 -17040 21132
rect -16976 16108 -16956 21132
rect -22328 16080 -16956 16108
rect -16716 21132 -11344 21160
rect -16716 16108 -11428 21132
rect -11364 16108 -11344 21132
rect -16716 16080 -11344 16108
rect -11104 21132 -5732 21160
rect -11104 16108 -5816 21132
rect -5752 16108 -5732 21132
rect -11104 16080 -5732 16108
rect -5492 21132 -120 21160
rect -5492 16108 -204 21132
rect -140 16108 -120 21132
rect -5492 16080 -120 16108
rect 120 21132 5492 21160
rect 120 16108 5408 21132
rect 5472 16108 5492 21132
rect 120 16080 5492 16108
rect 5732 21132 11104 21160
rect 5732 16108 11020 21132
rect 11084 16108 11104 21132
rect 5732 16080 11104 16108
rect 11344 21132 16716 21160
rect 11344 16108 16632 21132
rect 16696 16108 16716 21132
rect 11344 16080 16716 16108
rect 16956 21132 22328 21160
rect 16956 16108 22244 21132
rect 22308 16108 22328 21132
rect 16956 16080 22328 16108
rect -22328 15812 -16956 15840
rect -22328 10788 -17040 15812
rect -16976 10788 -16956 15812
rect -22328 10760 -16956 10788
rect -16716 15812 -11344 15840
rect -16716 10788 -11428 15812
rect -11364 10788 -11344 15812
rect -16716 10760 -11344 10788
rect -11104 15812 -5732 15840
rect -11104 10788 -5816 15812
rect -5752 10788 -5732 15812
rect -11104 10760 -5732 10788
rect -5492 15812 -120 15840
rect -5492 10788 -204 15812
rect -140 10788 -120 15812
rect -5492 10760 -120 10788
rect 120 15812 5492 15840
rect 120 10788 5408 15812
rect 5472 10788 5492 15812
rect 120 10760 5492 10788
rect 5732 15812 11104 15840
rect 5732 10788 11020 15812
rect 11084 10788 11104 15812
rect 5732 10760 11104 10788
rect 11344 15812 16716 15840
rect 11344 10788 16632 15812
rect 16696 10788 16716 15812
rect 11344 10760 16716 10788
rect 16956 15812 22328 15840
rect 16956 10788 22244 15812
rect 22308 10788 22328 15812
rect 16956 10760 22328 10788
rect -22328 10492 -16956 10520
rect -22328 5468 -17040 10492
rect -16976 5468 -16956 10492
rect -22328 5440 -16956 5468
rect -16716 10492 -11344 10520
rect -16716 5468 -11428 10492
rect -11364 5468 -11344 10492
rect -16716 5440 -11344 5468
rect -11104 10492 -5732 10520
rect -11104 5468 -5816 10492
rect -5752 5468 -5732 10492
rect -11104 5440 -5732 5468
rect -5492 10492 -120 10520
rect -5492 5468 -204 10492
rect -140 5468 -120 10492
rect -5492 5440 -120 5468
rect 120 10492 5492 10520
rect 120 5468 5408 10492
rect 5472 5468 5492 10492
rect 120 5440 5492 5468
rect 5732 10492 11104 10520
rect 5732 5468 11020 10492
rect 11084 5468 11104 10492
rect 5732 5440 11104 5468
rect 11344 10492 16716 10520
rect 11344 5468 16632 10492
rect 16696 5468 16716 10492
rect 11344 5440 16716 5468
rect 16956 10492 22328 10520
rect 16956 5468 22244 10492
rect 22308 5468 22328 10492
rect 16956 5440 22328 5468
rect -22328 5172 -16956 5200
rect -22328 148 -17040 5172
rect -16976 148 -16956 5172
rect -22328 120 -16956 148
rect -16716 5172 -11344 5200
rect -16716 148 -11428 5172
rect -11364 148 -11344 5172
rect -16716 120 -11344 148
rect -11104 5172 -5732 5200
rect -11104 148 -5816 5172
rect -5752 148 -5732 5172
rect -11104 120 -5732 148
rect -5492 5172 -120 5200
rect -5492 148 -204 5172
rect -140 148 -120 5172
rect -5492 120 -120 148
rect 120 5172 5492 5200
rect 120 148 5408 5172
rect 5472 148 5492 5172
rect 120 120 5492 148
rect 5732 5172 11104 5200
rect 5732 148 11020 5172
rect 11084 148 11104 5172
rect 5732 120 11104 148
rect 11344 5172 16716 5200
rect 11344 148 16632 5172
rect 16696 148 16716 5172
rect 11344 120 16716 148
rect 16956 5172 22328 5200
rect 16956 148 22244 5172
rect 22308 148 22328 5172
rect 16956 120 22328 148
rect -22328 -148 -16956 -120
rect -22328 -5172 -17040 -148
rect -16976 -5172 -16956 -148
rect -22328 -5200 -16956 -5172
rect -16716 -148 -11344 -120
rect -16716 -5172 -11428 -148
rect -11364 -5172 -11344 -148
rect -16716 -5200 -11344 -5172
rect -11104 -148 -5732 -120
rect -11104 -5172 -5816 -148
rect -5752 -5172 -5732 -148
rect -11104 -5200 -5732 -5172
rect -5492 -148 -120 -120
rect -5492 -5172 -204 -148
rect -140 -5172 -120 -148
rect -5492 -5200 -120 -5172
rect 120 -148 5492 -120
rect 120 -5172 5408 -148
rect 5472 -5172 5492 -148
rect 120 -5200 5492 -5172
rect 5732 -148 11104 -120
rect 5732 -5172 11020 -148
rect 11084 -5172 11104 -148
rect 5732 -5200 11104 -5172
rect 11344 -148 16716 -120
rect 11344 -5172 16632 -148
rect 16696 -5172 16716 -148
rect 11344 -5200 16716 -5172
rect 16956 -148 22328 -120
rect 16956 -5172 22244 -148
rect 22308 -5172 22328 -148
rect 16956 -5200 22328 -5172
rect -22328 -5468 -16956 -5440
rect -22328 -10492 -17040 -5468
rect -16976 -10492 -16956 -5468
rect -22328 -10520 -16956 -10492
rect -16716 -5468 -11344 -5440
rect -16716 -10492 -11428 -5468
rect -11364 -10492 -11344 -5468
rect -16716 -10520 -11344 -10492
rect -11104 -5468 -5732 -5440
rect -11104 -10492 -5816 -5468
rect -5752 -10492 -5732 -5468
rect -11104 -10520 -5732 -10492
rect -5492 -5468 -120 -5440
rect -5492 -10492 -204 -5468
rect -140 -10492 -120 -5468
rect -5492 -10520 -120 -10492
rect 120 -5468 5492 -5440
rect 120 -10492 5408 -5468
rect 5472 -10492 5492 -5468
rect 120 -10520 5492 -10492
rect 5732 -5468 11104 -5440
rect 5732 -10492 11020 -5468
rect 11084 -10492 11104 -5468
rect 5732 -10520 11104 -10492
rect 11344 -5468 16716 -5440
rect 11344 -10492 16632 -5468
rect 16696 -10492 16716 -5468
rect 11344 -10520 16716 -10492
rect 16956 -5468 22328 -5440
rect 16956 -10492 22244 -5468
rect 22308 -10492 22328 -5468
rect 16956 -10520 22328 -10492
rect -22328 -10788 -16956 -10760
rect -22328 -15812 -17040 -10788
rect -16976 -15812 -16956 -10788
rect -22328 -15840 -16956 -15812
rect -16716 -10788 -11344 -10760
rect -16716 -15812 -11428 -10788
rect -11364 -15812 -11344 -10788
rect -16716 -15840 -11344 -15812
rect -11104 -10788 -5732 -10760
rect -11104 -15812 -5816 -10788
rect -5752 -15812 -5732 -10788
rect -11104 -15840 -5732 -15812
rect -5492 -10788 -120 -10760
rect -5492 -15812 -204 -10788
rect -140 -15812 -120 -10788
rect -5492 -15840 -120 -15812
rect 120 -10788 5492 -10760
rect 120 -15812 5408 -10788
rect 5472 -15812 5492 -10788
rect 120 -15840 5492 -15812
rect 5732 -10788 11104 -10760
rect 5732 -15812 11020 -10788
rect 11084 -15812 11104 -10788
rect 5732 -15840 11104 -15812
rect 11344 -10788 16716 -10760
rect 11344 -15812 16632 -10788
rect 16696 -15812 16716 -10788
rect 11344 -15840 16716 -15812
rect 16956 -10788 22328 -10760
rect 16956 -15812 22244 -10788
rect 22308 -15812 22328 -10788
rect 16956 -15840 22328 -15812
rect -22328 -16108 -16956 -16080
rect -22328 -21132 -17040 -16108
rect -16976 -21132 -16956 -16108
rect -22328 -21160 -16956 -21132
rect -16716 -16108 -11344 -16080
rect -16716 -21132 -11428 -16108
rect -11364 -21132 -11344 -16108
rect -16716 -21160 -11344 -21132
rect -11104 -16108 -5732 -16080
rect -11104 -21132 -5816 -16108
rect -5752 -21132 -5732 -16108
rect -11104 -21160 -5732 -21132
rect -5492 -16108 -120 -16080
rect -5492 -21132 -204 -16108
rect -140 -21132 -120 -16108
rect -5492 -21160 -120 -21132
rect 120 -16108 5492 -16080
rect 120 -21132 5408 -16108
rect 5472 -21132 5492 -16108
rect 120 -21160 5492 -21132
rect 5732 -16108 11104 -16080
rect 5732 -21132 11020 -16108
rect 11084 -21132 11104 -16108
rect 5732 -21160 11104 -21132
rect 11344 -16108 16716 -16080
rect 11344 -21132 16632 -16108
rect 16696 -21132 16716 -16108
rect 11344 -21160 16716 -21132
rect 16956 -16108 22328 -16080
rect 16956 -21132 22244 -16108
rect 22308 -21132 22328 -16108
rect 16956 -21160 22328 -21132
<< via3 >>
rect -17040 16108 -16976 21132
rect -11428 16108 -11364 21132
rect -5816 16108 -5752 21132
rect -204 16108 -140 21132
rect 5408 16108 5472 21132
rect 11020 16108 11084 21132
rect 16632 16108 16696 21132
rect 22244 16108 22308 21132
rect -17040 10788 -16976 15812
rect -11428 10788 -11364 15812
rect -5816 10788 -5752 15812
rect -204 10788 -140 15812
rect 5408 10788 5472 15812
rect 11020 10788 11084 15812
rect 16632 10788 16696 15812
rect 22244 10788 22308 15812
rect -17040 5468 -16976 10492
rect -11428 5468 -11364 10492
rect -5816 5468 -5752 10492
rect -204 5468 -140 10492
rect 5408 5468 5472 10492
rect 11020 5468 11084 10492
rect 16632 5468 16696 10492
rect 22244 5468 22308 10492
rect -17040 148 -16976 5172
rect -11428 148 -11364 5172
rect -5816 148 -5752 5172
rect -204 148 -140 5172
rect 5408 148 5472 5172
rect 11020 148 11084 5172
rect 16632 148 16696 5172
rect 22244 148 22308 5172
rect -17040 -5172 -16976 -148
rect -11428 -5172 -11364 -148
rect -5816 -5172 -5752 -148
rect -204 -5172 -140 -148
rect 5408 -5172 5472 -148
rect 11020 -5172 11084 -148
rect 16632 -5172 16696 -148
rect 22244 -5172 22308 -148
rect -17040 -10492 -16976 -5468
rect -11428 -10492 -11364 -5468
rect -5816 -10492 -5752 -5468
rect -204 -10492 -140 -5468
rect 5408 -10492 5472 -5468
rect 11020 -10492 11084 -5468
rect 16632 -10492 16696 -5468
rect 22244 -10492 22308 -5468
rect -17040 -15812 -16976 -10788
rect -11428 -15812 -11364 -10788
rect -5816 -15812 -5752 -10788
rect -204 -15812 -140 -10788
rect 5408 -15812 5472 -10788
rect 11020 -15812 11084 -10788
rect 16632 -15812 16696 -10788
rect 22244 -15812 22308 -10788
rect -17040 -21132 -16976 -16108
rect -11428 -21132 -11364 -16108
rect -5816 -21132 -5752 -16108
rect -204 -21132 -140 -16108
rect 5408 -21132 5472 -16108
rect 11020 -21132 11084 -16108
rect 16632 -21132 16696 -16108
rect 22244 -21132 22308 -16108
<< mimcap >>
rect -22288 21080 -17288 21120
rect -22288 16160 -22248 21080
rect -17328 16160 -17288 21080
rect -22288 16120 -17288 16160
rect -16676 21080 -11676 21120
rect -16676 16160 -16636 21080
rect -11716 16160 -11676 21080
rect -16676 16120 -11676 16160
rect -11064 21080 -6064 21120
rect -11064 16160 -11024 21080
rect -6104 16160 -6064 21080
rect -11064 16120 -6064 16160
rect -5452 21080 -452 21120
rect -5452 16160 -5412 21080
rect -492 16160 -452 21080
rect -5452 16120 -452 16160
rect 160 21080 5160 21120
rect 160 16160 200 21080
rect 5120 16160 5160 21080
rect 160 16120 5160 16160
rect 5772 21080 10772 21120
rect 5772 16160 5812 21080
rect 10732 16160 10772 21080
rect 5772 16120 10772 16160
rect 11384 21080 16384 21120
rect 11384 16160 11424 21080
rect 16344 16160 16384 21080
rect 11384 16120 16384 16160
rect 16996 21080 21996 21120
rect 16996 16160 17036 21080
rect 21956 16160 21996 21080
rect 16996 16120 21996 16160
rect -22288 15760 -17288 15800
rect -22288 10840 -22248 15760
rect -17328 10840 -17288 15760
rect -22288 10800 -17288 10840
rect -16676 15760 -11676 15800
rect -16676 10840 -16636 15760
rect -11716 10840 -11676 15760
rect -16676 10800 -11676 10840
rect -11064 15760 -6064 15800
rect -11064 10840 -11024 15760
rect -6104 10840 -6064 15760
rect -11064 10800 -6064 10840
rect -5452 15760 -452 15800
rect -5452 10840 -5412 15760
rect -492 10840 -452 15760
rect -5452 10800 -452 10840
rect 160 15760 5160 15800
rect 160 10840 200 15760
rect 5120 10840 5160 15760
rect 160 10800 5160 10840
rect 5772 15760 10772 15800
rect 5772 10840 5812 15760
rect 10732 10840 10772 15760
rect 5772 10800 10772 10840
rect 11384 15760 16384 15800
rect 11384 10840 11424 15760
rect 16344 10840 16384 15760
rect 11384 10800 16384 10840
rect 16996 15760 21996 15800
rect 16996 10840 17036 15760
rect 21956 10840 21996 15760
rect 16996 10800 21996 10840
rect -22288 10440 -17288 10480
rect -22288 5520 -22248 10440
rect -17328 5520 -17288 10440
rect -22288 5480 -17288 5520
rect -16676 10440 -11676 10480
rect -16676 5520 -16636 10440
rect -11716 5520 -11676 10440
rect -16676 5480 -11676 5520
rect -11064 10440 -6064 10480
rect -11064 5520 -11024 10440
rect -6104 5520 -6064 10440
rect -11064 5480 -6064 5520
rect -5452 10440 -452 10480
rect -5452 5520 -5412 10440
rect -492 5520 -452 10440
rect -5452 5480 -452 5520
rect 160 10440 5160 10480
rect 160 5520 200 10440
rect 5120 5520 5160 10440
rect 160 5480 5160 5520
rect 5772 10440 10772 10480
rect 5772 5520 5812 10440
rect 10732 5520 10772 10440
rect 5772 5480 10772 5520
rect 11384 10440 16384 10480
rect 11384 5520 11424 10440
rect 16344 5520 16384 10440
rect 11384 5480 16384 5520
rect 16996 10440 21996 10480
rect 16996 5520 17036 10440
rect 21956 5520 21996 10440
rect 16996 5480 21996 5520
rect -22288 5120 -17288 5160
rect -22288 200 -22248 5120
rect -17328 200 -17288 5120
rect -22288 160 -17288 200
rect -16676 5120 -11676 5160
rect -16676 200 -16636 5120
rect -11716 200 -11676 5120
rect -16676 160 -11676 200
rect -11064 5120 -6064 5160
rect -11064 200 -11024 5120
rect -6104 200 -6064 5120
rect -11064 160 -6064 200
rect -5452 5120 -452 5160
rect -5452 200 -5412 5120
rect -492 200 -452 5120
rect -5452 160 -452 200
rect 160 5120 5160 5160
rect 160 200 200 5120
rect 5120 200 5160 5120
rect 160 160 5160 200
rect 5772 5120 10772 5160
rect 5772 200 5812 5120
rect 10732 200 10772 5120
rect 5772 160 10772 200
rect 11384 5120 16384 5160
rect 11384 200 11424 5120
rect 16344 200 16384 5120
rect 11384 160 16384 200
rect 16996 5120 21996 5160
rect 16996 200 17036 5120
rect 21956 200 21996 5120
rect 16996 160 21996 200
rect -22288 -200 -17288 -160
rect -22288 -5120 -22248 -200
rect -17328 -5120 -17288 -200
rect -22288 -5160 -17288 -5120
rect -16676 -200 -11676 -160
rect -16676 -5120 -16636 -200
rect -11716 -5120 -11676 -200
rect -16676 -5160 -11676 -5120
rect -11064 -200 -6064 -160
rect -11064 -5120 -11024 -200
rect -6104 -5120 -6064 -200
rect -11064 -5160 -6064 -5120
rect -5452 -200 -452 -160
rect -5452 -5120 -5412 -200
rect -492 -5120 -452 -200
rect -5452 -5160 -452 -5120
rect 160 -200 5160 -160
rect 160 -5120 200 -200
rect 5120 -5120 5160 -200
rect 160 -5160 5160 -5120
rect 5772 -200 10772 -160
rect 5772 -5120 5812 -200
rect 10732 -5120 10772 -200
rect 5772 -5160 10772 -5120
rect 11384 -200 16384 -160
rect 11384 -5120 11424 -200
rect 16344 -5120 16384 -200
rect 11384 -5160 16384 -5120
rect 16996 -200 21996 -160
rect 16996 -5120 17036 -200
rect 21956 -5120 21996 -200
rect 16996 -5160 21996 -5120
rect -22288 -5520 -17288 -5480
rect -22288 -10440 -22248 -5520
rect -17328 -10440 -17288 -5520
rect -22288 -10480 -17288 -10440
rect -16676 -5520 -11676 -5480
rect -16676 -10440 -16636 -5520
rect -11716 -10440 -11676 -5520
rect -16676 -10480 -11676 -10440
rect -11064 -5520 -6064 -5480
rect -11064 -10440 -11024 -5520
rect -6104 -10440 -6064 -5520
rect -11064 -10480 -6064 -10440
rect -5452 -5520 -452 -5480
rect -5452 -10440 -5412 -5520
rect -492 -10440 -452 -5520
rect -5452 -10480 -452 -10440
rect 160 -5520 5160 -5480
rect 160 -10440 200 -5520
rect 5120 -10440 5160 -5520
rect 160 -10480 5160 -10440
rect 5772 -5520 10772 -5480
rect 5772 -10440 5812 -5520
rect 10732 -10440 10772 -5520
rect 5772 -10480 10772 -10440
rect 11384 -5520 16384 -5480
rect 11384 -10440 11424 -5520
rect 16344 -10440 16384 -5520
rect 11384 -10480 16384 -10440
rect 16996 -5520 21996 -5480
rect 16996 -10440 17036 -5520
rect 21956 -10440 21996 -5520
rect 16996 -10480 21996 -10440
rect -22288 -10840 -17288 -10800
rect -22288 -15760 -22248 -10840
rect -17328 -15760 -17288 -10840
rect -22288 -15800 -17288 -15760
rect -16676 -10840 -11676 -10800
rect -16676 -15760 -16636 -10840
rect -11716 -15760 -11676 -10840
rect -16676 -15800 -11676 -15760
rect -11064 -10840 -6064 -10800
rect -11064 -15760 -11024 -10840
rect -6104 -15760 -6064 -10840
rect -11064 -15800 -6064 -15760
rect -5452 -10840 -452 -10800
rect -5452 -15760 -5412 -10840
rect -492 -15760 -452 -10840
rect -5452 -15800 -452 -15760
rect 160 -10840 5160 -10800
rect 160 -15760 200 -10840
rect 5120 -15760 5160 -10840
rect 160 -15800 5160 -15760
rect 5772 -10840 10772 -10800
rect 5772 -15760 5812 -10840
rect 10732 -15760 10772 -10840
rect 5772 -15800 10772 -15760
rect 11384 -10840 16384 -10800
rect 11384 -15760 11424 -10840
rect 16344 -15760 16384 -10840
rect 11384 -15800 16384 -15760
rect 16996 -10840 21996 -10800
rect 16996 -15760 17036 -10840
rect 21956 -15760 21996 -10840
rect 16996 -15800 21996 -15760
rect -22288 -16160 -17288 -16120
rect -22288 -21080 -22248 -16160
rect -17328 -21080 -17288 -16160
rect -22288 -21120 -17288 -21080
rect -16676 -16160 -11676 -16120
rect -16676 -21080 -16636 -16160
rect -11716 -21080 -11676 -16160
rect -16676 -21120 -11676 -21080
rect -11064 -16160 -6064 -16120
rect -11064 -21080 -11024 -16160
rect -6104 -21080 -6064 -16160
rect -11064 -21120 -6064 -21080
rect -5452 -16160 -452 -16120
rect -5452 -21080 -5412 -16160
rect -492 -21080 -452 -16160
rect -5452 -21120 -452 -21080
rect 160 -16160 5160 -16120
rect 160 -21080 200 -16160
rect 5120 -21080 5160 -16160
rect 160 -21120 5160 -21080
rect 5772 -16160 10772 -16120
rect 5772 -21080 5812 -16160
rect 10732 -21080 10772 -16160
rect 5772 -21120 10772 -21080
rect 11384 -16160 16384 -16120
rect 11384 -21080 11424 -16160
rect 16344 -21080 16384 -16160
rect 11384 -21120 16384 -21080
rect 16996 -16160 21996 -16120
rect 16996 -21080 17036 -16160
rect 21956 -21080 21996 -16160
rect 16996 -21120 21996 -21080
<< mimcapcontact >>
rect -22248 16160 -17328 21080
rect -16636 16160 -11716 21080
rect -11024 16160 -6104 21080
rect -5412 16160 -492 21080
rect 200 16160 5120 21080
rect 5812 16160 10732 21080
rect 11424 16160 16344 21080
rect 17036 16160 21956 21080
rect -22248 10840 -17328 15760
rect -16636 10840 -11716 15760
rect -11024 10840 -6104 15760
rect -5412 10840 -492 15760
rect 200 10840 5120 15760
rect 5812 10840 10732 15760
rect 11424 10840 16344 15760
rect 17036 10840 21956 15760
rect -22248 5520 -17328 10440
rect -16636 5520 -11716 10440
rect -11024 5520 -6104 10440
rect -5412 5520 -492 10440
rect 200 5520 5120 10440
rect 5812 5520 10732 10440
rect 11424 5520 16344 10440
rect 17036 5520 21956 10440
rect -22248 200 -17328 5120
rect -16636 200 -11716 5120
rect -11024 200 -6104 5120
rect -5412 200 -492 5120
rect 200 200 5120 5120
rect 5812 200 10732 5120
rect 11424 200 16344 5120
rect 17036 200 21956 5120
rect -22248 -5120 -17328 -200
rect -16636 -5120 -11716 -200
rect -11024 -5120 -6104 -200
rect -5412 -5120 -492 -200
rect 200 -5120 5120 -200
rect 5812 -5120 10732 -200
rect 11424 -5120 16344 -200
rect 17036 -5120 21956 -200
rect -22248 -10440 -17328 -5520
rect -16636 -10440 -11716 -5520
rect -11024 -10440 -6104 -5520
rect -5412 -10440 -492 -5520
rect 200 -10440 5120 -5520
rect 5812 -10440 10732 -5520
rect 11424 -10440 16344 -5520
rect 17036 -10440 21956 -5520
rect -22248 -15760 -17328 -10840
rect -16636 -15760 -11716 -10840
rect -11024 -15760 -6104 -10840
rect -5412 -15760 -492 -10840
rect 200 -15760 5120 -10840
rect 5812 -15760 10732 -10840
rect 11424 -15760 16344 -10840
rect 17036 -15760 21956 -10840
rect -22248 -21080 -17328 -16160
rect -16636 -21080 -11716 -16160
rect -11024 -21080 -6104 -16160
rect -5412 -21080 -492 -16160
rect 200 -21080 5120 -16160
rect 5812 -21080 10732 -16160
rect 11424 -21080 16344 -16160
rect 17036 -21080 21956 -16160
<< metal4 >>
rect -19840 21081 -19736 21280
rect -17060 21132 -16956 21280
rect -22249 21080 -17327 21081
rect -22249 16160 -22248 21080
rect -17328 16160 -17327 21080
rect -22249 16159 -17327 16160
rect -19840 15761 -19736 16159
rect -17060 16108 -17040 21132
rect -16976 16108 -16956 21132
rect -14228 21081 -14124 21280
rect -11448 21132 -11344 21280
rect -16637 21080 -11715 21081
rect -16637 16160 -16636 21080
rect -11716 16160 -11715 21080
rect -16637 16159 -11715 16160
rect -17060 15812 -16956 16108
rect -22249 15760 -17327 15761
rect -22249 10840 -22248 15760
rect -17328 10840 -17327 15760
rect -22249 10839 -17327 10840
rect -19840 10441 -19736 10839
rect -17060 10788 -17040 15812
rect -16976 10788 -16956 15812
rect -14228 15761 -14124 16159
rect -11448 16108 -11428 21132
rect -11364 16108 -11344 21132
rect -8616 21081 -8512 21280
rect -5836 21132 -5732 21280
rect -11025 21080 -6103 21081
rect -11025 16160 -11024 21080
rect -6104 16160 -6103 21080
rect -11025 16159 -6103 16160
rect -11448 15812 -11344 16108
rect -16637 15760 -11715 15761
rect -16637 10840 -16636 15760
rect -11716 10840 -11715 15760
rect -16637 10839 -11715 10840
rect -17060 10492 -16956 10788
rect -22249 10440 -17327 10441
rect -22249 5520 -22248 10440
rect -17328 5520 -17327 10440
rect -22249 5519 -17327 5520
rect -19840 5121 -19736 5519
rect -17060 5468 -17040 10492
rect -16976 5468 -16956 10492
rect -14228 10441 -14124 10839
rect -11448 10788 -11428 15812
rect -11364 10788 -11344 15812
rect -8616 15761 -8512 16159
rect -5836 16108 -5816 21132
rect -5752 16108 -5732 21132
rect -3004 21081 -2900 21280
rect -224 21132 -120 21280
rect -5413 21080 -491 21081
rect -5413 16160 -5412 21080
rect -492 16160 -491 21080
rect -5413 16159 -491 16160
rect -5836 15812 -5732 16108
rect -11025 15760 -6103 15761
rect -11025 10840 -11024 15760
rect -6104 10840 -6103 15760
rect -11025 10839 -6103 10840
rect -11448 10492 -11344 10788
rect -16637 10440 -11715 10441
rect -16637 5520 -16636 10440
rect -11716 5520 -11715 10440
rect -16637 5519 -11715 5520
rect -17060 5172 -16956 5468
rect -22249 5120 -17327 5121
rect -22249 200 -22248 5120
rect -17328 200 -17327 5120
rect -22249 199 -17327 200
rect -19840 -199 -19736 199
rect -17060 148 -17040 5172
rect -16976 148 -16956 5172
rect -14228 5121 -14124 5519
rect -11448 5468 -11428 10492
rect -11364 5468 -11344 10492
rect -8616 10441 -8512 10839
rect -5836 10788 -5816 15812
rect -5752 10788 -5732 15812
rect -3004 15761 -2900 16159
rect -224 16108 -204 21132
rect -140 16108 -120 21132
rect 2608 21081 2712 21280
rect 5388 21132 5492 21280
rect 199 21080 5121 21081
rect 199 16160 200 21080
rect 5120 16160 5121 21080
rect 199 16159 5121 16160
rect -224 15812 -120 16108
rect -5413 15760 -491 15761
rect -5413 10840 -5412 15760
rect -492 10840 -491 15760
rect -5413 10839 -491 10840
rect -5836 10492 -5732 10788
rect -11025 10440 -6103 10441
rect -11025 5520 -11024 10440
rect -6104 5520 -6103 10440
rect -11025 5519 -6103 5520
rect -11448 5172 -11344 5468
rect -16637 5120 -11715 5121
rect -16637 200 -16636 5120
rect -11716 200 -11715 5120
rect -16637 199 -11715 200
rect -17060 -148 -16956 148
rect -22249 -200 -17327 -199
rect -22249 -5120 -22248 -200
rect -17328 -5120 -17327 -200
rect -22249 -5121 -17327 -5120
rect -19840 -5519 -19736 -5121
rect -17060 -5172 -17040 -148
rect -16976 -5172 -16956 -148
rect -14228 -199 -14124 199
rect -11448 148 -11428 5172
rect -11364 148 -11344 5172
rect -8616 5121 -8512 5519
rect -5836 5468 -5816 10492
rect -5752 5468 -5732 10492
rect -3004 10441 -2900 10839
rect -224 10788 -204 15812
rect -140 10788 -120 15812
rect 2608 15761 2712 16159
rect 5388 16108 5408 21132
rect 5472 16108 5492 21132
rect 8220 21081 8324 21280
rect 11000 21132 11104 21280
rect 5811 21080 10733 21081
rect 5811 16160 5812 21080
rect 10732 16160 10733 21080
rect 5811 16159 10733 16160
rect 5388 15812 5492 16108
rect 199 15760 5121 15761
rect 199 10840 200 15760
rect 5120 10840 5121 15760
rect 199 10839 5121 10840
rect -224 10492 -120 10788
rect -5413 10440 -491 10441
rect -5413 5520 -5412 10440
rect -492 5520 -491 10440
rect -5413 5519 -491 5520
rect -5836 5172 -5732 5468
rect -11025 5120 -6103 5121
rect -11025 200 -11024 5120
rect -6104 200 -6103 5120
rect -11025 199 -6103 200
rect -11448 -148 -11344 148
rect -16637 -200 -11715 -199
rect -16637 -5120 -16636 -200
rect -11716 -5120 -11715 -200
rect -16637 -5121 -11715 -5120
rect -17060 -5468 -16956 -5172
rect -22249 -5520 -17327 -5519
rect -22249 -10440 -22248 -5520
rect -17328 -10440 -17327 -5520
rect -22249 -10441 -17327 -10440
rect -19840 -10839 -19736 -10441
rect -17060 -10492 -17040 -5468
rect -16976 -10492 -16956 -5468
rect -14228 -5519 -14124 -5121
rect -11448 -5172 -11428 -148
rect -11364 -5172 -11344 -148
rect -8616 -199 -8512 199
rect -5836 148 -5816 5172
rect -5752 148 -5732 5172
rect -3004 5121 -2900 5519
rect -224 5468 -204 10492
rect -140 5468 -120 10492
rect 2608 10441 2712 10839
rect 5388 10788 5408 15812
rect 5472 10788 5492 15812
rect 8220 15761 8324 16159
rect 11000 16108 11020 21132
rect 11084 16108 11104 21132
rect 13832 21081 13936 21280
rect 16612 21132 16716 21280
rect 11423 21080 16345 21081
rect 11423 16160 11424 21080
rect 16344 16160 16345 21080
rect 11423 16159 16345 16160
rect 11000 15812 11104 16108
rect 5811 15760 10733 15761
rect 5811 10840 5812 15760
rect 10732 10840 10733 15760
rect 5811 10839 10733 10840
rect 5388 10492 5492 10788
rect 199 10440 5121 10441
rect 199 5520 200 10440
rect 5120 5520 5121 10440
rect 199 5519 5121 5520
rect -224 5172 -120 5468
rect -5413 5120 -491 5121
rect -5413 200 -5412 5120
rect -492 200 -491 5120
rect -5413 199 -491 200
rect -5836 -148 -5732 148
rect -11025 -200 -6103 -199
rect -11025 -5120 -11024 -200
rect -6104 -5120 -6103 -200
rect -11025 -5121 -6103 -5120
rect -11448 -5468 -11344 -5172
rect -16637 -5520 -11715 -5519
rect -16637 -10440 -16636 -5520
rect -11716 -10440 -11715 -5520
rect -16637 -10441 -11715 -10440
rect -17060 -10788 -16956 -10492
rect -22249 -10840 -17327 -10839
rect -22249 -15760 -22248 -10840
rect -17328 -15760 -17327 -10840
rect -22249 -15761 -17327 -15760
rect -19840 -16159 -19736 -15761
rect -17060 -15812 -17040 -10788
rect -16976 -15812 -16956 -10788
rect -14228 -10839 -14124 -10441
rect -11448 -10492 -11428 -5468
rect -11364 -10492 -11344 -5468
rect -8616 -5519 -8512 -5121
rect -5836 -5172 -5816 -148
rect -5752 -5172 -5732 -148
rect -3004 -199 -2900 199
rect -224 148 -204 5172
rect -140 148 -120 5172
rect 2608 5121 2712 5519
rect 5388 5468 5408 10492
rect 5472 5468 5492 10492
rect 8220 10441 8324 10839
rect 11000 10788 11020 15812
rect 11084 10788 11104 15812
rect 13832 15761 13936 16159
rect 16612 16108 16632 21132
rect 16696 16108 16716 21132
rect 19444 21081 19548 21280
rect 22224 21132 22328 21280
rect 17035 21080 21957 21081
rect 17035 16160 17036 21080
rect 21956 16160 21957 21080
rect 17035 16159 21957 16160
rect 16612 15812 16716 16108
rect 11423 15760 16345 15761
rect 11423 10840 11424 15760
rect 16344 10840 16345 15760
rect 11423 10839 16345 10840
rect 11000 10492 11104 10788
rect 5811 10440 10733 10441
rect 5811 5520 5812 10440
rect 10732 5520 10733 10440
rect 5811 5519 10733 5520
rect 5388 5172 5492 5468
rect 199 5120 5121 5121
rect 199 200 200 5120
rect 5120 200 5121 5120
rect 199 199 5121 200
rect -224 -148 -120 148
rect -5413 -200 -491 -199
rect -5413 -5120 -5412 -200
rect -492 -5120 -491 -200
rect -5413 -5121 -491 -5120
rect -5836 -5468 -5732 -5172
rect -11025 -5520 -6103 -5519
rect -11025 -10440 -11024 -5520
rect -6104 -10440 -6103 -5520
rect -11025 -10441 -6103 -10440
rect -11448 -10788 -11344 -10492
rect -16637 -10840 -11715 -10839
rect -16637 -15760 -16636 -10840
rect -11716 -15760 -11715 -10840
rect -16637 -15761 -11715 -15760
rect -17060 -16108 -16956 -15812
rect -22249 -16160 -17327 -16159
rect -22249 -21080 -22248 -16160
rect -17328 -21080 -17327 -16160
rect -22249 -21081 -17327 -21080
rect -19840 -21280 -19736 -21081
rect -17060 -21132 -17040 -16108
rect -16976 -21132 -16956 -16108
rect -14228 -16159 -14124 -15761
rect -11448 -15812 -11428 -10788
rect -11364 -15812 -11344 -10788
rect -8616 -10839 -8512 -10441
rect -5836 -10492 -5816 -5468
rect -5752 -10492 -5732 -5468
rect -3004 -5519 -2900 -5121
rect -224 -5172 -204 -148
rect -140 -5172 -120 -148
rect 2608 -199 2712 199
rect 5388 148 5408 5172
rect 5472 148 5492 5172
rect 8220 5121 8324 5519
rect 11000 5468 11020 10492
rect 11084 5468 11104 10492
rect 13832 10441 13936 10839
rect 16612 10788 16632 15812
rect 16696 10788 16716 15812
rect 19444 15761 19548 16159
rect 22224 16108 22244 21132
rect 22308 16108 22328 21132
rect 22224 15812 22328 16108
rect 17035 15760 21957 15761
rect 17035 10840 17036 15760
rect 21956 10840 21957 15760
rect 17035 10839 21957 10840
rect 16612 10492 16716 10788
rect 11423 10440 16345 10441
rect 11423 5520 11424 10440
rect 16344 5520 16345 10440
rect 11423 5519 16345 5520
rect 11000 5172 11104 5468
rect 5811 5120 10733 5121
rect 5811 200 5812 5120
rect 10732 200 10733 5120
rect 5811 199 10733 200
rect 5388 -148 5492 148
rect 199 -200 5121 -199
rect 199 -5120 200 -200
rect 5120 -5120 5121 -200
rect 199 -5121 5121 -5120
rect -224 -5468 -120 -5172
rect -5413 -5520 -491 -5519
rect -5413 -10440 -5412 -5520
rect -492 -10440 -491 -5520
rect -5413 -10441 -491 -10440
rect -5836 -10788 -5732 -10492
rect -11025 -10840 -6103 -10839
rect -11025 -15760 -11024 -10840
rect -6104 -15760 -6103 -10840
rect -11025 -15761 -6103 -15760
rect -11448 -16108 -11344 -15812
rect -16637 -16160 -11715 -16159
rect -16637 -21080 -16636 -16160
rect -11716 -21080 -11715 -16160
rect -16637 -21081 -11715 -21080
rect -17060 -21280 -16956 -21132
rect -14228 -21280 -14124 -21081
rect -11448 -21132 -11428 -16108
rect -11364 -21132 -11344 -16108
rect -8616 -16159 -8512 -15761
rect -5836 -15812 -5816 -10788
rect -5752 -15812 -5732 -10788
rect -3004 -10839 -2900 -10441
rect -224 -10492 -204 -5468
rect -140 -10492 -120 -5468
rect 2608 -5519 2712 -5121
rect 5388 -5172 5408 -148
rect 5472 -5172 5492 -148
rect 8220 -199 8324 199
rect 11000 148 11020 5172
rect 11084 148 11104 5172
rect 13832 5121 13936 5519
rect 16612 5468 16632 10492
rect 16696 5468 16716 10492
rect 19444 10441 19548 10839
rect 22224 10788 22244 15812
rect 22308 10788 22328 15812
rect 22224 10492 22328 10788
rect 17035 10440 21957 10441
rect 17035 5520 17036 10440
rect 21956 5520 21957 10440
rect 17035 5519 21957 5520
rect 16612 5172 16716 5468
rect 11423 5120 16345 5121
rect 11423 200 11424 5120
rect 16344 200 16345 5120
rect 11423 199 16345 200
rect 11000 -148 11104 148
rect 5811 -200 10733 -199
rect 5811 -5120 5812 -200
rect 10732 -5120 10733 -200
rect 5811 -5121 10733 -5120
rect 5388 -5468 5492 -5172
rect 199 -5520 5121 -5519
rect 199 -10440 200 -5520
rect 5120 -10440 5121 -5520
rect 199 -10441 5121 -10440
rect -224 -10788 -120 -10492
rect -5413 -10840 -491 -10839
rect -5413 -15760 -5412 -10840
rect -492 -15760 -491 -10840
rect -5413 -15761 -491 -15760
rect -5836 -16108 -5732 -15812
rect -11025 -16160 -6103 -16159
rect -11025 -21080 -11024 -16160
rect -6104 -21080 -6103 -16160
rect -11025 -21081 -6103 -21080
rect -11448 -21280 -11344 -21132
rect -8616 -21280 -8512 -21081
rect -5836 -21132 -5816 -16108
rect -5752 -21132 -5732 -16108
rect -3004 -16159 -2900 -15761
rect -224 -15812 -204 -10788
rect -140 -15812 -120 -10788
rect 2608 -10839 2712 -10441
rect 5388 -10492 5408 -5468
rect 5472 -10492 5492 -5468
rect 8220 -5519 8324 -5121
rect 11000 -5172 11020 -148
rect 11084 -5172 11104 -148
rect 13832 -199 13936 199
rect 16612 148 16632 5172
rect 16696 148 16716 5172
rect 19444 5121 19548 5519
rect 22224 5468 22244 10492
rect 22308 5468 22328 10492
rect 22224 5172 22328 5468
rect 17035 5120 21957 5121
rect 17035 200 17036 5120
rect 21956 200 21957 5120
rect 17035 199 21957 200
rect 16612 -148 16716 148
rect 11423 -200 16345 -199
rect 11423 -5120 11424 -200
rect 16344 -5120 16345 -200
rect 11423 -5121 16345 -5120
rect 11000 -5468 11104 -5172
rect 5811 -5520 10733 -5519
rect 5811 -10440 5812 -5520
rect 10732 -10440 10733 -5520
rect 5811 -10441 10733 -10440
rect 5388 -10788 5492 -10492
rect 199 -10840 5121 -10839
rect 199 -15760 200 -10840
rect 5120 -15760 5121 -10840
rect 199 -15761 5121 -15760
rect -224 -16108 -120 -15812
rect -5413 -16160 -491 -16159
rect -5413 -21080 -5412 -16160
rect -492 -21080 -491 -16160
rect -5413 -21081 -491 -21080
rect -5836 -21280 -5732 -21132
rect -3004 -21280 -2900 -21081
rect -224 -21132 -204 -16108
rect -140 -21132 -120 -16108
rect 2608 -16159 2712 -15761
rect 5388 -15812 5408 -10788
rect 5472 -15812 5492 -10788
rect 8220 -10839 8324 -10441
rect 11000 -10492 11020 -5468
rect 11084 -10492 11104 -5468
rect 13832 -5519 13936 -5121
rect 16612 -5172 16632 -148
rect 16696 -5172 16716 -148
rect 19444 -199 19548 199
rect 22224 148 22244 5172
rect 22308 148 22328 5172
rect 22224 -148 22328 148
rect 17035 -200 21957 -199
rect 17035 -5120 17036 -200
rect 21956 -5120 21957 -200
rect 17035 -5121 21957 -5120
rect 16612 -5468 16716 -5172
rect 11423 -5520 16345 -5519
rect 11423 -10440 11424 -5520
rect 16344 -10440 16345 -5520
rect 11423 -10441 16345 -10440
rect 11000 -10788 11104 -10492
rect 5811 -10840 10733 -10839
rect 5811 -15760 5812 -10840
rect 10732 -15760 10733 -10840
rect 5811 -15761 10733 -15760
rect 5388 -16108 5492 -15812
rect 199 -16160 5121 -16159
rect 199 -21080 200 -16160
rect 5120 -21080 5121 -16160
rect 199 -21081 5121 -21080
rect -224 -21280 -120 -21132
rect 2608 -21280 2712 -21081
rect 5388 -21132 5408 -16108
rect 5472 -21132 5492 -16108
rect 8220 -16159 8324 -15761
rect 11000 -15812 11020 -10788
rect 11084 -15812 11104 -10788
rect 13832 -10839 13936 -10441
rect 16612 -10492 16632 -5468
rect 16696 -10492 16716 -5468
rect 19444 -5519 19548 -5121
rect 22224 -5172 22244 -148
rect 22308 -5172 22328 -148
rect 22224 -5468 22328 -5172
rect 17035 -5520 21957 -5519
rect 17035 -10440 17036 -5520
rect 21956 -10440 21957 -5520
rect 17035 -10441 21957 -10440
rect 16612 -10788 16716 -10492
rect 11423 -10840 16345 -10839
rect 11423 -15760 11424 -10840
rect 16344 -15760 16345 -10840
rect 11423 -15761 16345 -15760
rect 11000 -16108 11104 -15812
rect 5811 -16160 10733 -16159
rect 5811 -21080 5812 -16160
rect 10732 -21080 10733 -16160
rect 5811 -21081 10733 -21080
rect 5388 -21280 5492 -21132
rect 8220 -21280 8324 -21081
rect 11000 -21132 11020 -16108
rect 11084 -21132 11104 -16108
rect 13832 -16159 13936 -15761
rect 16612 -15812 16632 -10788
rect 16696 -15812 16716 -10788
rect 19444 -10839 19548 -10441
rect 22224 -10492 22244 -5468
rect 22308 -10492 22328 -5468
rect 22224 -10788 22328 -10492
rect 17035 -10840 21957 -10839
rect 17035 -15760 17036 -10840
rect 21956 -15760 21957 -10840
rect 17035 -15761 21957 -15760
rect 16612 -16108 16716 -15812
rect 11423 -16160 16345 -16159
rect 11423 -21080 11424 -16160
rect 16344 -21080 16345 -16160
rect 11423 -21081 16345 -21080
rect 11000 -21280 11104 -21132
rect 13832 -21280 13936 -21081
rect 16612 -21132 16632 -16108
rect 16696 -21132 16716 -16108
rect 19444 -16159 19548 -15761
rect 22224 -15812 22244 -10788
rect 22308 -15812 22328 -10788
rect 22224 -16108 22328 -15812
rect 17035 -16160 21957 -16159
rect 17035 -21080 17036 -16160
rect 21956 -21080 21957 -16160
rect 17035 -21081 21957 -21080
rect 16612 -21280 16716 -21132
rect 19444 -21280 19548 -21081
rect 22224 -21132 22244 -16108
rect 22308 -21132 22328 -16108
rect 22224 -21280 22328 -21132
<< properties >>
string FIXED_BBOX 16956 16080 22036 21160
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 25.0 val 1.269k carea 2.00 cperi 0.19 class capacitor nx 8 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
