magic
tech sky130A
magscale 1 2
timestamp 1769172933
<< error_p >>
rect -1747 568 1747 572
rect -1747 -500 -1717 568
rect -1681 502 -1315 506
rect -1253 502 -887 506
rect -825 502 -459 506
rect -397 502 -31 506
rect 31 502 397 506
rect 459 502 825 506
rect 887 502 1253 506
rect 1315 502 1681 506
rect -1681 -434 -1651 502
rect 1651 -434 1681 502
rect 1717 -500 1747 568
<< nwell >>
rect -1717 -534 1717 568
<< mvpmos >>
rect -1623 -434 -1373 506
rect -1195 -434 -945 506
rect -767 -434 -517 506
rect -339 -434 -89 506
rect 89 -434 339 506
rect 517 -434 767 506
rect 945 -434 1195 506
rect 1373 -434 1623 506
<< mvpdiff >>
rect -1681 494 -1623 506
rect -1681 -422 -1669 494
rect -1635 -422 -1623 494
rect -1681 -434 -1623 -422
rect -1373 494 -1315 506
rect -1373 -422 -1361 494
rect -1327 -422 -1315 494
rect -1373 -434 -1315 -422
rect -1253 494 -1195 506
rect -1253 -422 -1241 494
rect -1207 -422 -1195 494
rect -1253 -434 -1195 -422
rect -945 494 -887 506
rect -945 -422 -933 494
rect -899 -422 -887 494
rect -945 -434 -887 -422
rect -825 494 -767 506
rect -825 -422 -813 494
rect -779 -422 -767 494
rect -825 -434 -767 -422
rect -517 494 -459 506
rect -517 -422 -505 494
rect -471 -422 -459 494
rect -517 -434 -459 -422
rect -397 494 -339 506
rect -397 -422 -385 494
rect -351 -422 -339 494
rect -397 -434 -339 -422
rect -89 494 -31 506
rect -89 -422 -77 494
rect -43 -422 -31 494
rect -89 -434 -31 -422
rect 31 494 89 506
rect 31 -422 43 494
rect 77 -422 89 494
rect 31 -434 89 -422
rect 339 494 397 506
rect 339 -422 351 494
rect 385 -422 397 494
rect 339 -434 397 -422
rect 459 494 517 506
rect 459 -422 471 494
rect 505 -422 517 494
rect 459 -434 517 -422
rect 767 494 825 506
rect 767 -422 779 494
rect 813 -422 825 494
rect 767 -434 825 -422
rect 887 494 945 506
rect 887 -422 899 494
rect 933 -422 945 494
rect 887 -434 945 -422
rect 1195 494 1253 506
rect 1195 -422 1207 494
rect 1241 -422 1253 494
rect 1195 -434 1253 -422
rect 1315 494 1373 506
rect 1315 -422 1327 494
rect 1361 -422 1373 494
rect 1315 -434 1373 -422
rect 1623 494 1681 506
rect 1623 -422 1635 494
rect 1669 -422 1681 494
rect 1623 -434 1681 -422
<< mvpdiffc >>
rect -1669 -422 -1635 494
rect -1361 -422 -1327 494
rect -1241 -422 -1207 494
rect -933 -422 -899 494
rect -813 -422 -779 494
rect -505 -422 -471 494
rect -385 -422 -351 494
rect -77 -422 -43 494
rect 43 -422 77 494
rect 351 -422 385 494
rect 471 -422 505 494
rect 779 -422 813 494
rect 899 -422 933 494
rect 1207 -422 1241 494
rect 1327 -422 1361 494
rect 1635 -422 1669 494
<< poly >>
rect -1623 506 -1373 532
rect -1195 506 -945 532
rect -767 506 -517 532
rect -339 506 -89 532
rect 89 506 339 532
rect 517 506 767 532
rect 945 506 1195 532
rect 1373 506 1623 532
rect -1623 -481 -1373 -434
rect -1623 -515 -1607 -481
rect -1389 -515 -1373 -481
rect -1623 -531 -1373 -515
rect -1195 -481 -945 -434
rect -1195 -515 -1179 -481
rect -961 -515 -945 -481
rect -1195 -531 -945 -515
rect -767 -481 -517 -434
rect -767 -515 -751 -481
rect -533 -515 -517 -481
rect -767 -531 -517 -515
rect -339 -481 -89 -434
rect -339 -515 -323 -481
rect -105 -515 -89 -481
rect -339 -531 -89 -515
rect 89 -481 339 -434
rect 89 -515 105 -481
rect 323 -515 339 -481
rect 89 -531 339 -515
rect 517 -481 767 -434
rect 517 -515 533 -481
rect 751 -515 767 -481
rect 517 -531 767 -515
rect 945 -481 1195 -434
rect 945 -515 961 -481
rect 1179 -515 1195 -481
rect 945 -531 1195 -515
rect 1373 -481 1623 -434
rect 1373 -515 1389 -481
rect 1607 -515 1623 -481
rect 1373 -531 1623 -515
<< polycont >>
rect -1607 -515 -1389 -481
rect -1179 -515 -961 -481
rect -751 -515 -533 -481
rect -323 -515 -105 -481
rect 105 -515 323 -481
rect 533 -515 751 -481
rect 961 -515 1179 -481
rect 1389 -515 1607 -481
<< locali >>
rect -1669 494 -1635 510
rect -1669 -438 -1635 -422
rect -1361 494 -1327 510
rect -1361 -438 -1327 -422
rect -1241 494 -1207 510
rect -1241 -438 -1207 -422
rect -933 494 -899 510
rect -933 -438 -899 -422
rect -813 494 -779 510
rect -813 -438 -779 -422
rect -505 494 -471 510
rect -505 -438 -471 -422
rect -385 494 -351 510
rect -385 -438 -351 -422
rect -77 494 -43 510
rect -77 -438 -43 -422
rect 43 494 77 510
rect 43 -438 77 -422
rect 351 494 385 510
rect 351 -438 385 -422
rect 471 494 505 510
rect 471 -438 505 -422
rect 779 494 813 510
rect 779 -438 813 -422
rect 899 494 933 510
rect 899 -438 933 -422
rect 1207 494 1241 510
rect 1207 -438 1241 -422
rect 1327 494 1361 510
rect 1327 -438 1361 -422
rect 1635 494 1669 510
rect 1635 -438 1669 -422
rect -1623 -515 -1607 -481
rect -1389 -515 -1373 -481
rect -1195 -515 -1179 -481
rect -961 -515 -945 -481
rect -767 -515 -751 -481
rect -533 -515 -517 -481
rect -339 -515 -323 -481
rect -105 -515 -89 -481
rect 89 -515 105 -481
rect 323 -515 339 -481
rect 517 -515 533 -481
rect 751 -515 767 -481
rect 945 -515 961 -481
rect 1179 -515 1195 -481
rect 1373 -515 1389 -481
rect 1607 -515 1623 -481
<< viali >>
rect -1669 -422 -1635 494
rect -1361 -422 -1327 494
rect -1241 -422 -1207 494
rect -933 -422 -899 494
rect -813 -422 -779 494
rect -505 -422 -471 494
rect -385 -422 -351 494
rect -77 -422 -43 494
rect 43 -422 77 494
rect 351 -422 385 494
rect 471 -422 505 494
rect 779 -422 813 494
rect 899 -422 933 494
rect 1207 -422 1241 494
rect 1327 -422 1361 494
rect 1635 -422 1669 494
rect -1607 -515 -1389 -481
rect -1179 -515 -961 -481
rect -751 -515 -533 -481
rect -323 -515 -105 -481
rect 105 -515 323 -481
rect 533 -515 751 -481
rect 961 -515 1179 -481
rect 1389 -515 1607 -481
<< metal1 >>
rect -1675 494 -1629 506
rect -1675 -422 -1669 494
rect -1635 -422 -1629 494
rect -1675 -434 -1629 -422
rect -1367 494 -1321 506
rect -1367 -422 -1361 494
rect -1327 -422 -1321 494
rect -1367 -434 -1321 -422
rect -1247 494 -1201 506
rect -1247 -422 -1241 494
rect -1207 -422 -1201 494
rect -1247 -434 -1201 -422
rect -939 494 -893 506
rect -939 -422 -933 494
rect -899 -422 -893 494
rect -939 -434 -893 -422
rect -819 494 -773 506
rect -819 -422 -813 494
rect -779 -422 -773 494
rect -819 -434 -773 -422
rect -511 494 -465 506
rect -511 -422 -505 494
rect -471 -422 -465 494
rect -511 -434 -465 -422
rect -391 494 -345 506
rect -391 -422 -385 494
rect -351 -422 -345 494
rect -391 -434 -345 -422
rect -83 494 -37 506
rect -83 -422 -77 494
rect -43 -422 -37 494
rect -83 -434 -37 -422
rect 37 494 83 506
rect 37 -422 43 494
rect 77 -422 83 494
rect 37 -434 83 -422
rect 345 494 391 506
rect 345 -422 351 494
rect 385 -422 391 494
rect 345 -434 391 -422
rect 465 494 511 506
rect 465 -422 471 494
rect 505 -422 511 494
rect 465 -434 511 -422
rect 773 494 819 506
rect 773 -422 779 494
rect 813 -422 819 494
rect 773 -434 819 -422
rect 893 494 939 506
rect 893 -422 899 494
rect 933 -422 939 494
rect 893 -434 939 -422
rect 1201 494 1247 506
rect 1201 -422 1207 494
rect 1241 -422 1247 494
rect 1201 -434 1247 -422
rect 1321 494 1367 506
rect 1321 -422 1327 494
rect 1361 -422 1367 494
rect 1321 -434 1367 -422
rect 1629 494 1675 506
rect 1629 -422 1635 494
rect 1669 -422 1675 494
rect 1629 -434 1675 -422
rect -1619 -481 -1377 -475
rect -1619 -515 -1607 -481
rect -1389 -515 -1377 -481
rect -1619 -521 -1377 -515
rect -1191 -481 -949 -475
rect -1191 -515 -1179 -481
rect -961 -515 -949 -481
rect -1191 -521 -949 -515
rect -763 -481 -521 -475
rect -763 -515 -751 -481
rect -533 -515 -521 -481
rect -763 -521 -521 -515
rect -335 -481 -93 -475
rect -335 -515 -323 -481
rect -105 -515 -93 -481
rect -335 -521 -93 -515
rect 93 -481 335 -475
rect 93 -515 105 -481
rect 323 -515 335 -481
rect 93 -521 335 -515
rect 521 -481 763 -475
rect 521 -515 533 -481
rect 751 -515 763 -481
rect 521 -521 763 -515
rect 949 -481 1191 -475
rect 949 -515 961 -481
rect 1179 -515 1191 -481
rect 949 -521 1191 -515
rect 1377 -481 1619 -475
rect 1377 -515 1389 -481
rect 1607 -515 1619 -481
rect 1377 -521 1619 -515
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.7 l 1.25 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
