magic
tech sky130A
magscale 1 2
timestamp 1769529800
<< pwell >>
rect -515 -729 515 729
<< mvnmos >>
rect -287 -471 -187 471
rect -129 -471 -29 471
rect 29 -471 129 471
rect 187 -471 287 471
<< mvndiff >>
rect -345 459 -287 471
rect -345 -459 -333 459
rect -299 -459 -287 459
rect -345 -471 -287 -459
rect -187 459 -129 471
rect -187 -459 -175 459
rect -141 -459 -129 459
rect -187 -471 -129 -459
rect -29 459 29 471
rect -29 -459 -17 459
rect 17 -459 29 459
rect -29 -471 29 -459
rect 129 459 187 471
rect 129 -459 141 459
rect 175 -459 187 459
rect 129 -471 187 -459
rect 287 459 345 471
rect 287 -459 299 459
rect 333 -459 345 459
rect 287 -471 345 -459
<< mvndiffc >>
rect -333 -459 -299 459
rect -175 -459 -141 459
rect -17 -459 17 459
rect 141 -459 175 459
rect 299 -459 333 459
<< mvpsubdiff >>
rect -479 681 479 693
rect -479 647 -371 681
rect 371 647 479 681
rect -479 635 479 647
rect -479 585 -421 635
rect -479 -585 -467 585
rect -433 -585 -421 585
rect 421 585 479 635
rect -479 -635 -421 -585
rect 421 -585 433 585
rect 467 -585 479 585
rect 421 -635 479 -585
rect -479 -647 479 -635
rect -479 -681 -371 -647
rect 371 -681 479 -647
rect -479 -693 479 -681
<< mvpsubdiffcont >>
rect -371 647 371 681
rect -467 -585 -433 585
rect 433 -585 467 585
rect -371 -681 371 -647
<< poly >>
rect -287 543 -187 559
rect -287 509 -271 543
rect -203 509 -187 543
rect -287 471 -187 509
rect -129 543 -29 559
rect -129 509 -113 543
rect -45 509 -29 543
rect -129 471 -29 509
rect 29 543 129 559
rect 29 509 45 543
rect 113 509 129 543
rect 29 471 129 509
rect 187 543 287 559
rect 187 509 203 543
rect 271 509 287 543
rect 187 471 287 509
rect -287 -509 -187 -471
rect -287 -543 -271 -509
rect -203 -543 -187 -509
rect -287 -559 -187 -543
rect -129 -509 -29 -471
rect -129 -543 -113 -509
rect -45 -543 -29 -509
rect -129 -559 -29 -543
rect 29 -509 129 -471
rect 29 -543 45 -509
rect 113 -543 129 -509
rect 29 -559 129 -543
rect 187 -509 287 -471
rect 187 -543 203 -509
rect 271 -543 287 -509
rect 187 -559 287 -543
<< polycont >>
rect -271 509 -203 543
rect -113 509 -45 543
rect 45 509 113 543
rect 203 509 271 543
rect -271 -543 -203 -509
rect -113 -543 -45 -509
rect 45 -543 113 -509
rect 203 -543 271 -509
<< locali >>
rect -467 647 -371 681
rect 371 647 467 681
rect -467 585 -433 647
rect 433 585 467 647
rect -287 509 -271 543
rect -203 509 -187 543
rect -129 509 -113 543
rect -45 509 -29 543
rect 29 509 45 543
rect 113 509 129 543
rect 187 509 203 543
rect 271 509 287 543
rect -333 459 -299 475
rect -333 -475 -299 -459
rect -175 459 -141 475
rect -175 -475 -141 -459
rect -17 459 17 475
rect -17 -475 17 -459
rect 141 459 175 475
rect 141 -475 175 -459
rect 299 459 333 475
rect 299 -475 333 -459
rect -287 -543 -271 -509
rect -203 -543 -187 -509
rect -129 -543 -113 -509
rect -45 -543 -29 -509
rect 29 -543 45 -509
rect 113 -543 129 -509
rect 187 -543 203 -509
rect 271 -543 287 -509
rect -467 -647 -433 -585
rect 433 -647 467 -585
rect -467 -681 -371 -647
rect 371 -681 467 -647
<< viali >>
rect -271 509 -203 543
rect -113 509 -45 543
rect 45 509 113 543
rect 203 509 271 543
rect -333 -459 -299 459
rect -175 -459 -141 459
rect -17 -459 17 459
rect 141 -459 175 459
rect 299 -459 333 459
rect -271 -543 -203 -509
rect -113 -543 -45 -509
rect 45 -543 113 -509
rect 203 -543 271 -509
<< metal1 >>
rect -283 543 -191 549
rect -283 509 -271 543
rect -203 509 -191 543
rect -283 503 -191 509
rect -125 543 -33 549
rect -125 509 -113 543
rect -45 509 -33 543
rect -125 503 -33 509
rect 33 543 125 549
rect 33 509 45 543
rect 113 509 125 543
rect 33 503 125 509
rect 191 543 283 549
rect 191 509 203 543
rect 271 509 283 543
rect 191 503 283 509
rect -339 459 -293 471
rect -339 -459 -333 459
rect -299 -459 -293 459
rect -339 -471 -293 -459
rect -181 459 -135 471
rect -181 -459 -175 459
rect -141 -459 -135 459
rect -181 -471 -135 -459
rect -23 459 23 471
rect -23 -459 -17 459
rect 17 -459 23 459
rect -23 -471 23 -459
rect 135 459 181 471
rect 135 -459 141 459
rect 175 -459 181 459
rect 135 -471 181 -459
rect 293 459 339 471
rect 293 -459 299 459
rect 333 -459 339 459
rect 293 -471 339 -459
rect -283 -509 -191 -503
rect -283 -543 -271 -509
rect -203 -543 -191 -509
rect -283 -549 -191 -543
rect -125 -509 -33 -503
rect -125 -543 -113 -509
rect -45 -543 -33 -509
rect -125 -549 -33 -543
rect 33 -509 125 -503
rect 33 -543 45 -509
rect 113 -543 125 -509
rect 33 -549 125 -543
rect 191 -509 283 -503
rect 191 -543 203 -509
rect 271 -543 283 -509
rect 191 -549 283 -543
<< properties >>
string FIXED_BBOX -450 -664 450 664
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.7125 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
