magic
tech sky130A
magscale 1 2
timestamp 1769436194
<< mvnmos >>
rect -17703 -2031 -17603 1969
rect -17425 -2031 -17325 1969
rect -17147 -2031 -17047 1969
rect -16869 -2031 -16769 1969
rect -16591 -2031 -16491 1969
rect -16313 -2031 -16213 1969
rect -16035 -2031 -15935 1969
rect -15757 -2031 -15657 1969
rect -15479 -2031 -15379 1969
rect -15201 -2031 -15101 1969
rect -14923 -2031 -14823 1969
rect -14645 -2031 -14545 1969
rect -14367 -2031 -14267 1969
rect -14089 -2031 -13989 1969
rect -13811 -2031 -13711 1969
rect -13533 -2031 -13433 1969
rect -13255 -2031 -13155 1969
rect -12977 -2031 -12877 1969
rect -12699 -2031 -12599 1969
rect -12421 -2031 -12321 1969
rect -12143 -2031 -12043 1969
rect -11865 -2031 -11765 1969
rect -11587 -2031 -11487 1969
rect -11309 -2031 -11209 1969
rect -11031 -2031 -10931 1969
rect -10753 -2031 -10653 1969
rect -10475 -2031 -10375 1969
rect -10197 -2031 -10097 1969
rect -9919 -2031 -9819 1969
rect -9641 -2031 -9541 1969
rect -9363 -2031 -9263 1969
rect -9085 -2031 -8985 1969
rect -8807 -2031 -8707 1969
rect -8529 -2031 -8429 1969
rect -8251 -2031 -8151 1969
rect -7973 -2031 -7873 1969
rect -7695 -2031 -7595 1969
rect -7417 -2031 -7317 1969
rect -7139 -2031 -7039 1969
rect -6861 -2031 -6761 1969
rect -6583 -2031 -6483 1969
rect -6305 -2031 -6205 1969
rect -6027 -2031 -5927 1969
rect -5749 -2031 -5649 1969
rect -5471 -2031 -5371 1969
rect -5193 -2031 -5093 1969
rect -4915 -2031 -4815 1969
rect -4637 -2031 -4537 1969
rect -4359 -2031 -4259 1969
rect -4081 -2031 -3981 1969
rect -3803 -2031 -3703 1969
rect -3525 -2031 -3425 1969
rect -3247 -2031 -3147 1969
rect -2969 -2031 -2869 1969
rect -2691 -2031 -2591 1969
rect -2413 -2031 -2313 1969
rect -2135 -2031 -2035 1969
rect -1857 -2031 -1757 1969
rect -1579 -2031 -1479 1969
rect -1301 -2031 -1201 1969
rect -1023 -2031 -923 1969
rect -745 -2031 -645 1969
rect -467 -2031 -367 1969
rect -189 -2031 -89 1969
rect 89 -2031 189 1969
rect 367 -2031 467 1969
rect 645 -2031 745 1969
rect 923 -2031 1023 1969
rect 1201 -2031 1301 1969
rect 1479 -2031 1579 1969
rect 1757 -2031 1857 1969
rect 2035 -2031 2135 1969
rect 2313 -2031 2413 1969
rect 2591 -2031 2691 1969
rect 2869 -2031 2969 1969
rect 3147 -2031 3247 1969
rect 3425 -2031 3525 1969
rect 3703 -2031 3803 1969
rect 3981 -2031 4081 1969
rect 4259 -2031 4359 1969
rect 4537 -2031 4637 1969
rect 4815 -2031 4915 1969
rect 5093 -2031 5193 1969
rect 5371 -2031 5471 1969
rect 5649 -2031 5749 1969
rect 5927 -2031 6027 1969
rect 6205 -2031 6305 1969
rect 6483 -2031 6583 1969
rect 6761 -2031 6861 1969
rect 7039 -2031 7139 1969
rect 7317 -2031 7417 1969
rect 7595 -2031 7695 1969
rect 7873 -2031 7973 1969
rect 8151 -2031 8251 1969
rect 8429 -2031 8529 1969
rect 8707 -2031 8807 1969
rect 8985 -2031 9085 1969
rect 9263 -2031 9363 1969
rect 9541 -2031 9641 1969
rect 9819 -2031 9919 1969
rect 10097 -2031 10197 1969
rect 10375 -2031 10475 1969
rect 10653 -2031 10753 1969
rect 10931 -2031 11031 1969
rect 11209 -2031 11309 1969
rect 11487 -2031 11587 1969
rect 11765 -2031 11865 1969
rect 12043 -2031 12143 1969
rect 12321 -2031 12421 1969
rect 12599 -2031 12699 1969
rect 12877 -2031 12977 1969
rect 13155 -2031 13255 1969
rect 13433 -2031 13533 1969
rect 13711 -2031 13811 1969
rect 13989 -2031 14089 1969
rect 14267 -2031 14367 1969
rect 14545 -2031 14645 1969
rect 14823 -2031 14923 1969
rect 15101 -2031 15201 1969
rect 15379 -2031 15479 1969
rect 15657 -2031 15757 1969
rect 15935 -2031 16035 1969
rect 16213 -2031 16313 1969
rect 16491 -2031 16591 1969
rect 16769 -2031 16869 1969
rect 17047 -2031 17147 1969
rect 17325 -2031 17425 1969
rect 17603 -2031 17703 1969
<< mvndiff >>
rect -17761 1957 -17703 1969
rect -17761 -2019 -17749 1957
rect -17715 -2019 -17703 1957
rect -17761 -2031 -17703 -2019
rect -17603 1957 -17545 1969
rect -17603 -2019 -17591 1957
rect -17557 -2019 -17545 1957
rect -17603 -2031 -17545 -2019
rect -17483 1957 -17425 1969
rect -17483 -2019 -17471 1957
rect -17437 -2019 -17425 1957
rect -17483 -2031 -17425 -2019
rect -17325 1957 -17267 1969
rect -17325 -2019 -17313 1957
rect -17279 -2019 -17267 1957
rect -17325 -2031 -17267 -2019
rect -17205 1957 -17147 1969
rect -17205 -2019 -17193 1957
rect -17159 -2019 -17147 1957
rect -17205 -2031 -17147 -2019
rect -17047 1957 -16989 1969
rect -17047 -2019 -17035 1957
rect -17001 -2019 -16989 1957
rect -17047 -2031 -16989 -2019
rect -16927 1957 -16869 1969
rect -16927 -2019 -16915 1957
rect -16881 -2019 -16869 1957
rect -16927 -2031 -16869 -2019
rect -16769 1957 -16711 1969
rect -16769 -2019 -16757 1957
rect -16723 -2019 -16711 1957
rect -16769 -2031 -16711 -2019
rect -16649 1957 -16591 1969
rect -16649 -2019 -16637 1957
rect -16603 -2019 -16591 1957
rect -16649 -2031 -16591 -2019
rect -16491 1957 -16433 1969
rect -16491 -2019 -16479 1957
rect -16445 -2019 -16433 1957
rect -16491 -2031 -16433 -2019
rect -16371 1957 -16313 1969
rect -16371 -2019 -16359 1957
rect -16325 -2019 -16313 1957
rect -16371 -2031 -16313 -2019
rect -16213 1957 -16155 1969
rect -16213 -2019 -16201 1957
rect -16167 -2019 -16155 1957
rect -16213 -2031 -16155 -2019
rect -16093 1957 -16035 1969
rect -16093 -2019 -16081 1957
rect -16047 -2019 -16035 1957
rect -16093 -2031 -16035 -2019
rect -15935 1957 -15877 1969
rect -15935 -2019 -15923 1957
rect -15889 -2019 -15877 1957
rect -15935 -2031 -15877 -2019
rect -15815 1957 -15757 1969
rect -15815 -2019 -15803 1957
rect -15769 -2019 -15757 1957
rect -15815 -2031 -15757 -2019
rect -15657 1957 -15599 1969
rect -15657 -2019 -15645 1957
rect -15611 -2019 -15599 1957
rect -15657 -2031 -15599 -2019
rect -15537 1957 -15479 1969
rect -15537 -2019 -15525 1957
rect -15491 -2019 -15479 1957
rect -15537 -2031 -15479 -2019
rect -15379 1957 -15321 1969
rect -15379 -2019 -15367 1957
rect -15333 -2019 -15321 1957
rect -15379 -2031 -15321 -2019
rect -15259 1957 -15201 1969
rect -15259 -2019 -15247 1957
rect -15213 -2019 -15201 1957
rect -15259 -2031 -15201 -2019
rect -15101 1957 -15043 1969
rect -15101 -2019 -15089 1957
rect -15055 -2019 -15043 1957
rect -15101 -2031 -15043 -2019
rect -14981 1957 -14923 1969
rect -14981 -2019 -14969 1957
rect -14935 -2019 -14923 1957
rect -14981 -2031 -14923 -2019
rect -14823 1957 -14765 1969
rect -14823 -2019 -14811 1957
rect -14777 -2019 -14765 1957
rect -14823 -2031 -14765 -2019
rect -14703 1957 -14645 1969
rect -14703 -2019 -14691 1957
rect -14657 -2019 -14645 1957
rect -14703 -2031 -14645 -2019
rect -14545 1957 -14487 1969
rect -14545 -2019 -14533 1957
rect -14499 -2019 -14487 1957
rect -14545 -2031 -14487 -2019
rect -14425 1957 -14367 1969
rect -14425 -2019 -14413 1957
rect -14379 -2019 -14367 1957
rect -14425 -2031 -14367 -2019
rect -14267 1957 -14209 1969
rect -14267 -2019 -14255 1957
rect -14221 -2019 -14209 1957
rect -14267 -2031 -14209 -2019
rect -14147 1957 -14089 1969
rect -14147 -2019 -14135 1957
rect -14101 -2019 -14089 1957
rect -14147 -2031 -14089 -2019
rect -13989 1957 -13931 1969
rect -13989 -2019 -13977 1957
rect -13943 -2019 -13931 1957
rect -13989 -2031 -13931 -2019
rect -13869 1957 -13811 1969
rect -13869 -2019 -13857 1957
rect -13823 -2019 -13811 1957
rect -13869 -2031 -13811 -2019
rect -13711 1957 -13653 1969
rect -13711 -2019 -13699 1957
rect -13665 -2019 -13653 1957
rect -13711 -2031 -13653 -2019
rect -13591 1957 -13533 1969
rect -13591 -2019 -13579 1957
rect -13545 -2019 -13533 1957
rect -13591 -2031 -13533 -2019
rect -13433 1957 -13375 1969
rect -13433 -2019 -13421 1957
rect -13387 -2019 -13375 1957
rect -13433 -2031 -13375 -2019
rect -13313 1957 -13255 1969
rect -13313 -2019 -13301 1957
rect -13267 -2019 -13255 1957
rect -13313 -2031 -13255 -2019
rect -13155 1957 -13097 1969
rect -13155 -2019 -13143 1957
rect -13109 -2019 -13097 1957
rect -13155 -2031 -13097 -2019
rect -13035 1957 -12977 1969
rect -13035 -2019 -13023 1957
rect -12989 -2019 -12977 1957
rect -13035 -2031 -12977 -2019
rect -12877 1957 -12819 1969
rect -12877 -2019 -12865 1957
rect -12831 -2019 -12819 1957
rect -12877 -2031 -12819 -2019
rect -12757 1957 -12699 1969
rect -12757 -2019 -12745 1957
rect -12711 -2019 -12699 1957
rect -12757 -2031 -12699 -2019
rect -12599 1957 -12541 1969
rect -12599 -2019 -12587 1957
rect -12553 -2019 -12541 1957
rect -12599 -2031 -12541 -2019
rect -12479 1957 -12421 1969
rect -12479 -2019 -12467 1957
rect -12433 -2019 -12421 1957
rect -12479 -2031 -12421 -2019
rect -12321 1957 -12263 1969
rect -12321 -2019 -12309 1957
rect -12275 -2019 -12263 1957
rect -12321 -2031 -12263 -2019
rect -12201 1957 -12143 1969
rect -12201 -2019 -12189 1957
rect -12155 -2019 -12143 1957
rect -12201 -2031 -12143 -2019
rect -12043 1957 -11985 1969
rect -12043 -2019 -12031 1957
rect -11997 -2019 -11985 1957
rect -12043 -2031 -11985 -2019
rect -11923 1957 -11865 1969
rect -11923 -2019 -11911 1957
rect -11877 -2019 -11865 1957
rect -11923 -2031 -11865 -2019
rect -11765 1957 -11707 1969
rect -11765 -2019 -11753 1957
rect -11719 -2019 -11707 1957
rect -11765 -2031 -11707 -2019
rect -11645 1957 -11587 1969
rect -11645 -2019 -11633 1957
rect -11599 -2019 -11587 1957
rect -11645 -2031 -11587 -2019
rect -11487 1957 -11429 1969
rect -11487 -2019 -11475 1957
rect -11441 -2019 -11429 1957
rect -11487 -2031 -11429 -2019
rect -11367 1957 -11309 1969
rect -11367 -2019 -11355 1957
rect -11321 -2019 -11309 1957
rect -11367 -2031 -11309 -2019
rect -11209 1957 -11151 1969
rect -11209 -2019 -11197 1957
rect -11163 -2019 -11151 1957
rect -11209 -2031 -11151 -2019
rect -11089 1957 -11031 1969
rect -11089 -2019 -11077 1957
rect -11043 -2019 -11031 1957
rect -11089 -2031 -11031 -2019
rect -10931 1957 -10873 1969
rect -10931 -2019 -10919 1957
rect -10885 -2019 -10873 1957
rect -10931 -2031 -10873 -2019
rect -10811 1957 -10753 1969
rect -10811 -2019 -10799 1957
rect -10765 -2019 -10753 1957
rect -10811 -2031 -10753 -2019
rect -10653 1957 -10595 1969
rect -10653 -2019 -10641 1957
rect -10607 -2019 -10595 1957
rect -10653 -2031 -10595 -2019
rect -10533 1957 -10475 1969
rect -10533 -2019 -10521 1957
rect -10487 -2019 -10475 1957
rect -10533 -2031 -10475 -2019
rect -10375 1957 -10317 1969
rect -10375 -2019 -10363 1957
rect -10329 -2019 -10317 1957
rect -10375 -2031 -10317 -2019
rect -10255 1957 -10197 1969
rect -10255 -2019 -10243 1957
rect -10209 -2019 -10197 1957
rect -10255 -2031 -10197 -2019
rect -10097 1957 -10039 1969
rect -10097 -2019 -10085 1957
rect -10051 -2019 -10039 1957
rect -10097 -2031 -10039 -2019
rect -9977 1957 -9919 1969
rect -9977 -2019 -9965 1957
rect -9931 -2019 -9919 1957
rect -9977 -2031 -9919 -2019
rect -9819 1957 -9761 1969
rect -9819 -2019 -9807 1957
rect -9773 -2019 -9761 1957
rect -9819 -2031 -9761 -2019
rect -9699 1957 -9641 1969
rect -9699 -2019 -9687 1957
rect -9653 -2019 -9641 1957
rect -9699 -2031 -9641 -2019
rect -9541 1957 -9483 1969
rect -9541 -2019 -9529 1957
rect -9495 -2019 -9483 1957
rect -9541 -2031 -9483 -2019
rect -9421 1957 -9363 1969
rect -9421 -2019 -9409 1957
rect -9375 -2019 -9363 1957
rect -9421 -2031 -9363 -2019
rect -9263 1957 -9205 1969
rect -9263 -2019 -9251 1957
rect -9217 -2019 -9205 1957
rect -9263 -2031 -9205 -2019
rect -9143 1957 -9085 1969
rect -9143 -2019 -9131 1957
rect -9097 -2019 -9085 1957
rect -9143 -2031 -9085 -2019
rect -8985 1957 -8927 1969
rect -8985 -2019 -8973 1957
rect -8939 -2019 -8927 1957
rect -8985 -2031 -8927 -2019
rect -8865 1957 -8807 1969
rect -8865 -2019 -8853 1957
rect -8819 -2019 -8807 1957
rect -8865 -2031 -8807 -2019
rect -8707 1957 -8649 1969
rect -8707 -2019 -8695 1957
rect -8661 -2019 -8649 1957
rect -8707 -2031 -8649 -2019
rect -8587 1957 -8529 1969
rect -8587 -2019 -8575 1957
rect -8541 -2019 -8529 1957
rect -8587 -2031 -8529 -2019
rect -8429 1957 -8371 1969
rect -8429 -2019 -8417 1957
rect -8383 -2019 -8371 1957
rect -8429 -2031 -8371 -2019
rect -8309 1957 -8251 1969
rect -8309 -2019 -8297 1957
rect -8263 -2019 -8251 1957
rect -8309 -2031 -8251 -2019
rect -8151 1957 -8093 1969
rect -8151 -2019 -8139 1957
rect -8105 -2019 -8093 1957
rect -8151 -2031 -8093 -2019
rect -8031 1957 -7973 1969
rect -8031 -2019 -8019 1957
rect -7985 -2019 -7973 1957
rect -8031 -2031 -7973 -2019
rect -7873 1957 -7815 1969
rect -7873 -2019 -7861 1957
rect -7827 -2019 -7815 1957
rect -7873 -2031 -7815 -2019
rect -7753 1957 -7695 1969
rect -7753 -2019 -7741 1957
rect -7707 -2019 -7695 1957
rect -7753 -2031 -7695 -2019
rect -7595 1957 -7537 1969
rect -7595 -2019 -7583 1957
rect -7549 -2019 -7537 1957
rect -7595 -2031 -7537 -2019
rect -7475 1957 -7417 1969
rect -7475 -2019 -7463 1957
rect -7429 -2019 -7417 1957
rect -7475 -2031 -7417 -2019
rect -7317 1957 -7259 1969
rect -7317 -2019 -7305 1957
rect -7271 -2019 -7259 1957
rect -7317 -2031 -7259 -2019
rect -7197 1957 -7139 1969
rect -7197 -2019 -7185 1957
rect -7151 -2019 -7139 1957
rect -7197 -2031 -7139 -2019
rect -7039 1957 -6981 1969
rect -7039 -2019 -7027 1957
rect -6993 -2019 -6981 1957
rect -7039 -2031 -6981 -2019
rect -6919 1957 -6861 1969
rect -6919 -2019 -6907 1957
rect -6873 -2019 -6861 1957
rect -6919 -2031 -6861 -2019
rect -6761 1957 -6703 1969
rect -6761 -2019 -6749 1957
rect -6715 -2019 -6703 1957
rect -6761 -2031 -6703 -2019
rect -6641 1957 -6583 1969
rect -6641 -2019 -6629 1957
rect -6595 -2019 -6583 1957
rect -6641 -2031 -6583 -2019
rect -6483 1957 -6425 1969
rect -6483 -2019 -6471 1957
rect -6437 -2019 -6425 1957
rect -6483 -2031 -6425 -2019
rect -6363 1957 -6305 1969
rect -6363 -2019 -6351 1957
rect -6317 -2019 -6305 1957
rect -6363 -2031 -6305 -2019
rect -6205 1957 -6147 1969
rect -6205 -2019 -6193 1957
rect -6159 -2019 -6147 1957
rect -6205 -2031 -6147 -2019
rect -6085 1957 -6027 1969
rect -6085 -2019 -6073 1957
rect -6039 -2019 -6027 1957
rect -6085 -2031 -6027 -2019
rect -5927 1957 -5869 1969
rect -5927 -2019 -5915 1957
rect -5881 -2019 -5869 1957
rect -5927 -2031 -5869 -2019
rect -5807 1957 -5749 1969
rect -5807 -2019 -5795 1957
rect -5761 -2019 -5749 1957
rect -5807 -2031 -5749 -2019
rect -5649 1957 -5591 1969
rect -5649 -2019 -5637 1957
rect -5603 -2019 -5591 1957
rect -5649 -2031 -5591 -2019
rect -5529 1957 -5471 1969
rect -5529 -2019 -5517 1957
rect -5483 -2019 -5471 1957
rect -5529 -2031 -5471 -2019
rect -5371 1957 -5313 1969
rect -5371 -2019 -5359 1957
rect -5325 -2019 -5313 1957
rect -5371 -2031 -5313 -2019
rect -5251 1957 -5193 1969
rect -5251 -2019 -5239 1957
rect -5205 -2019 -5193 1957
rect -5251 -2031 -5193 -2019
rect -5093 1957 -5035 1969
rect -5093 -2019 -5081 1957
rect -5047 -2019 -5035 1957
rect -5093 -2031 -5035 -2019
rect -4973 1957 -4915 1969
rect -4973 -2019 -4961 1957
rect -4927 -2019 -4915 1957
rect -4973 -2031 -4915 -2019
rect -4815 1957 -4757 1969
rect -4815 -2019 -4803 1957
rect -4769 -2019 -4757 1957
rect -4815 -2031 -4757 -2019
rect -4695 1957 -4637 1969
rect -4695 -2019 -4683 1957
rect -4649 -2019 -4637 1957
rect -4695 -2031 -4637 -2019
rect -4537 1957 -4479 1969
rect -4537 -2019 -4525 1957
rect -4491 -2019 -4479 1957
rect -4537 -2031 -4479 -2019
rect -4417 1957 -4359 1969
rect -4417 -2019 -4405 1957
rect -4371 -2019 -4359 1957
rect -4417 -2031 -4359 -2019
rect -4259 1957 -4201 1969
rect -4259 -2019 -4247 1957
rect -4213 -2019 -4201 1957
rect -4259 -2031 -4201 -2019
rect -4139 1957 -4081 1969
rect -4139 -2019 -4127 1957
rect -4093 -2019 -4081 1957
rect -4139 -2031 -4081 -2019
rect -3981 1957 -3923 1969
rect -3981 -2019 -3969 1957
rect -3935 -2019 -3923 1957
rect -3981 -2031 -3923 -2019
rect -3861 1957 -3803 1969
rect -3861 -2019 -3849 1957
rect -3815 -2019 -3803 1957
rect -3861 -2031 -3803 -2019
rect -3703 1957 -3645 1969
rect -3703 -2019 -3691 1957
rect -3657 -2019 -3645 1957
rect -3703 -2031 -3645 -2019
rect -3583 1957 -3525 1969
rect -3583 -2019 -3571 1957
rect -3537 -2019 -3525 1957
rect -3583 -2031 -3525 -2019
rect -3425 1957 -3367 1969
rect -3425 -2019 -3413 1957
rect -3379 -2019 -3367 1957
rect -3425 -2031 -3367 -2019
rect -3305 1957 -3247 1969
rect -3305 -2019 -3293 1957
rect -3259 -2019 -3247 1957
rect -3305 -2031 -3247 -2019
rect -3147 1957 -3089 1969
rect -3147 -2019 -3135 1957
rect -3101 -2019 -3089 1957
rect -3147 -2031 -3089 -2019
rect -3027 1957 -2969 1969
rect -3027 -2019 -3015 1957
rect -2981 -2019 -2969 1957
rect -3027 -2031 -2969 -2019
rect -2869 1957 -2811 1969
rect -2869 -2019 -2857 1957
rect -2823 -2019 -2811 1957
rect -2869 -2031 -2811 -2019
rect -2749 1957 -2691 1969
rect -2749 -2019 -2737 1957
rect -2703 -2019 -2691 1957
rect -2749 -2031 -2691 -2019
rect -2591 1957 -2533 1969
rect -2591 -2019 -2579 1957
rect -2545 -2019 -2533 1957
rect -2591 -2031 -2533 -2019
rect -2471 1957 -2413 1969
rect -2471 -2019 -2459 1957
rect -2425 -2019 -2413 1957
rect -2471 -2031 -2413 -2019
rect -2313 1957 -2255 1969
rect -2313 -2019 -2301 1957
rect -2267 -2019 -2255 1957
rect -2313 -2031 -2255 -2019
rect -2193 1957 -2135 1969
rect -2193 -2019 -2181 1957
rect -2147 -2019 -2135 1957
rect -2193 -2031 -2135 -2019
rect -2035 1957 -1977 1969
rect -2035 -2019 -2023 1957
rect -1989 -2019 -1977 1957
rect -2035 -2031 -1977 -2019
rect -1915 1957 -1857 1969
rect -1915 -2019 -1903 1957
rect -1869 -2019 -1857 1957
rect -1915 -2031 -1857 -2019
rect -1757 1957 -1699 1969
rect -1757 -2019 -1745 1957
rect -1711 -2019 -1699 1957
rect -1757 -2031 -1699 -2019
rect -1637 1957 -1579 1969
rect -1637 -2019 -1625 1957
rect -1591 -2019 -1579 1957
rect -1637 -2031 -1579 -2019
rect -1479 1957 -1421 1969
rect -1479 -2019 -1467 1957
rect -1433 -2019 -1421 1957
rect -1479 -2031 -1421 -2019
rect -1359 1957 -1301 1969
rect -1359 -2019 -1347 1957
rect -1313 -2019 -1301 1957
rect -1359 -2031 -1301 -2019
rect -1201 1957 -1143 1969
rect -1201 -2019 -1189 1957
rect -1155 -2019 -1143 1957
rect -1201 -2031 -1143 -2019
rect -1081 1957 -1023 1969
rect -1081 -2019 -1069 1957
rect -1035 -2019 -1023 1957
rect -1081 -2031 -1023 -2019
rect -923 1957 -865 1969
rect -923 -2019 -911 1957
rect -877 -2019 -865 1957
rect -923 -2031 -865 -2019
rect -803 1957 -745 1969
rect -803 -2019 -791 1957
rect -757 -2019 -745 1957
rect -803 -2031 -745 -2019
rect -645 1957 -587 1969
rect -645 -2019 -633 1957
rect -599 -2019 -587 1957
rect -645 -2031 -587 -2019
rect -525 1957 -467 1969
rect -525 -2019 -513 1957
rect -479 -2019 -467 1957
rect -525 -2031 -467 -2019
rect -367 1957 -309 1969
rect -367 -2019 -355 1957
rect -321 -2019 -309 1957
rect -367 -2031 -309 -2019
rect -247 1957 -189 1969
rect -247 -2019 -235 1957
rect -201 -2019 -189 1957
rect -247 -2031 -189 -2019
rect -89 1957 -31 1969
rect -89 -2019 -77 1957
rect -43 -2019 -31 1957
rect -89 -2031 -31 -2019
rect 31 1957 89 1969
rect 31 -2019 43 1957
rect 77 -2019 89 1957
rect 31 -2031 89 -2019
rect 189 1957 247 1969
rect 189 -2019 201 1957
rect 235 -2019 247 1957
rect 189 -2031 247 -2019
rect 309 1957 367 1969
rect 309 -2019 321 1957
rect 355 -2019 367 1957
rect 309 -2031 367 -2019
rect 467 1957 525 1969
rect 467 -2019 479 1957
rect 513 -2019 525 1957
rect 467 -2031 525 -2019
rect 587 1957 645 1969
rect 587 -2019 599 1957
rect 633 -2019 645 1957
rect 587 -2031 645 -2019
rect 745 1957 803 1969
rect 745 -2019 757 1957
rect 791 -2019 803 1957
rect 745 -2031 803 -2019
rect 865 1957 923 1969
rect 865 -2019 877 1957
rect 911 -2019 923 1957
rect 865 -2031 923 -2019
rect 1023 1957 1081 1969
rect 1023 -2019 1035 1957
rect 1069 -2019 1081 1957
rect 1023 -2031 1081 -2019
rect 1143 1957 1201 1969
rect 1143 -2019 1155 1957
rect 1189 -2019 1201 1957
rect 1143 -2031 1201 -2019
rect 1301 1957 1359 1969
rect 1301 -2019 1313 1957
rect 1347 -2019 1359 1957
rect 1301 -2031 1359 -2019
rect 1421 1957 1479 1969
rect 1421 -2019 1433 1957
rect 1467 -2019 1479 1957
rect 1421 -2031 1479 -2019
rect 1579 1957 1637 1969
rect 1579 -2019 1591 1957
rect 1625 -2019 1637 1957
rect 1579 -2031 1637 -2019
rect 1699 1957 1757 1969
rect 1699 -2019 1711 1957
rect 1745 -2019 1757 1957
rect 1699 -2031 1757 -2019
rect 1857 1957 1915 1969
rect 1857 -2019 1869 1957
rect 1903 -2019 1915 1957
rect 1857 -2031 1915 -2019
rect 1977 1957 2035 1969
rect 1977 -2019 1989 1957
rect 2023 -2019 2035 1957
rect 1977 -2031 2035 -2019
rect 2135 1957 2193 1969
rect 2135 -2019 2147 1957
rect 2181 -2019 2193 1957
rect 2135 -2031 2193 -2019
rect 2255 1957 2313 1969
rect 2255 -2019 2267 1957
rect 2301 -2019 2313 1957
rect 2255 -2031 2313 -2019
rect 2413 1957 2471 1969
rect 2413 -2019 2425 1957
rect 2459 -2019 2471 1957
rect 2413 -2031 2471 -2019
rect 2533 1957 2591 1969
rect 2533 -2019 2545 1957
rect 2579 -2019 2591 1957
rect 2533 -2031 2591 -2019
rect 2691 1957 2749 1969
rect 2691 -2019 2703 1957
rect 2737 -2019 2749 1957
rect 2691 -2031 2749 -2019
rect 2811 1957 2869 1969
rect 2811 -2019 2823 1957
rect 2857 -2019 2869 1957
rect 2811 -2031 2869 -2019
rect 2969 1957 3027 1969
rect 2969 -2019 2981 1957
rect 3015 -2019 3027 1957
rect 2969 -2031 3027 -2019
rect 3089 1957 3147 1969
rect 3089 -2019 3101 1957
rect 3135 -2019 3147 1957
rect 3089 -2031 3147 -2019
rect 3247 1957 3305 1969
rect 3247 -2019 3259 1957
rect 3293 -2019 3305 1957
rect 3247 -2031 3305 -2019
rect 3367 1957 3425 1969
rect 3367 -2019 3379 1957
rect 3413 -2019 3425 1957
rect 3367 -2031 3425 -2019
rect 3525 1957 3583 1969
rect 3525 -2019 3537 1957
rect 3571 -2019 3583 1957
rect 3525 -2031 3583 -2019
rect 3645 1957 3703 1969
rect 3645 -2019 3657 1957
rect 3691 -2019 3703 1957
rect 3645 -2031 3703 -2019
rect 3803 1957 3861 1969
rect 3803 -2019 3815 1957
rect 3849 -2019 3861 1957
rect 3803 -2031 3861 -2019
rect 3923 1957 3981 1969
rect 3923 -2019 3935 1957
rect 3969 -2019 3981 1957
rect 3923 -2031 3981 -2019
rect 4081 1957 4139 1969
rect 4081 -2019 4093 1957
rect 4127 -2019 4139 1957
rect 4081 -2031 4139 -2019
rect 4201 1957 4259 1969
rect 4201 -2019 4213 1957
rect 4247 -2019 4259 1957
rect 4201 -2031 4259 -2019
rect 4359 1957 4417 1969
rect 4359 -2019 4371 1957
rect 4405 -2019 4417 1957
rect 4359 -2031 4417 -2019
rect 4479 1957 4537 1969
rect 4479 -2019 4491 1957
rect 4525 -2019 4537 1957
rect 4479 -2031 4537 -2019
rect 4637 1957 4695 1969
rect 4637 -2019 4649 1957
rect 4683 -2019 4695 1957
rect 4637 -2031 4695 -2019
rect 4757 1957 4815 1969
rect 4757 -2019 4769 1957
rect 4803 -2019 4815 1957
rect 4757 -2031 4815 -2019
rect 4915 1957 4973 1969
rect 4915 -2019 4927 1957
rect 4961 -2019 4973 1957
rect 4915 -2031 4973 -2019
rect 5035 1957 5093 1969
rect 5035 -2019 5047 1957
rect 5081 -2019 5093 1957
rect 5035 -2031 5093 -2019
rect 5193 1957 5251 1969
rect 5193 -2019 5205 1957
rect 5239 -2019 5251 1957
rect 5193 -2031 5251 -2019
rect 5313 1957 5371 1969
rect 5313 -2019 5325 1957
rect 5359 -2019 5371 1957
rect 5313 -2031 5371 -2019
rect 5471 1957 5529 1969
rect 5471 -2019 5483 1957
rect 5517 -2019 5529 1957
rect 5471 -2031 5529 -2019
rect 5591 1957 5649 1969
rect 5591 -2019 5603 1957
rect 5637 -2019 5649 1957
rect 5591 -2031 5649 -2019
rect 5749 1957 5807 1969
rect 5749 -2019 5761 1957
rect 5795 -2019 5807 1957
rect 5749 -2031 5807 -2019
rect 5869 1957 5927 1969
rect 5869 -2019 5881 1957
rect 5915 -2019 5927 1957
rect 5869 -2031 5927 -2019
rect 6027 1957 6085 1969
rect 6027 -2019 6039 1957
rect 6073 -2019 6085 1957
rect 6027 -2031 6085 -2019
rect 6147 1957 6205 1969
rect 6147 -2019 6159 1957
rect 6193 -2019 6205 1957
rect 6147 -2031 6205 -2019
rect 6305 1957 6363 1969
rect 6305 -2019 6317 1957
rect 6351 -2019 6363 1957
rect 6305 -2031 6363 -2019
rect 6425 1957 6483 1969
rect 6425 -2019 6437 1957
rect 6471 -2019 6483 1957
rect 6425 -2031 6483 -2019
rect 6583 1957 6641 1969
rect 6583 -2019 6595 1957
rect 6629 -2019 6641 1957
rect 6583 -2031 6641 -2019
rect 6703 1957 6761 1969
rect 6703 -2019 6715 1957
rect 6749 -2019 6761 1957
rect 6703 -2031 6761 -2019
rect 6861 1957 6919 1969
rect 6861 -2019 6873 1957
rect 6907 -2019 6919 1957
rect 6861 -2031 6919 -2019
rect 6981 1957 7039 1969
rect 6981 -2019 6993 1957
rect 7027 -2019 7039 1957
rect 6981 -2031 7039 -2019
rect 7139 1957 7197 1969
rect 7139 -2019 7151 1957
rect 7185 -2019 7197 1957
rect 7139 -2031 7197 -2019
rect 7259 1957 7317 1969
rect 7259 -2019 7271 1957
rect 7305 -2019 7317 1957
rect 7259 -2031 7317 -2019
rect 7417 1957 7475 1969
rect 7417 -2019 7429 1957
rect 7463 -2019 7475 1957
rect 7417 -2031 7475 -2019
rect 7537 1957 7595 1969
rect 7537 -2019 7549 1957
rect 7583 -2019 7595 1957
rect 7537 -2031 7595 -2019
rect 7695 1957 7753 1969
rect 7695 -2019 7707 1957
rect 7741 -2019 7753 1957
rect 7695 -2031 7753 -2019
rect 7815 1957 7873 1969
rect 7815 -2019 7827 1957
rect 7861 -2019 7873 1957
rect 7815 -2031 7873 -2019
rect 7973 1957 8031 1969
rect 7973 -2019 7985 1957
rect 8019 -2019 8031 1957
rect 7973 -2031 8031 -2019
rect 8093 1957 8151 1969
rect 8093 -2019 8105 1957
rect 8139 -2019 8151 1957
rect 8093 -2031 8151 -2019
rect 8251 1957 8309 1969
rect 8251 -2019 8263 1957
rect 8297 -2019 8309 1957
rect 8251 -2031 8309 -2019
rect 8371 1957 8429 1969
rect 8371 -2019 8383 1957
rect 8417 -2019 8429 1957
rect 8371 -2031 8429 -2019
rect 8529 1957 8587 1969
rect 8529 -2019 8541 1957
rect 8575 -2019 8587 1957
rect 8529 -2031 8587 -2019
rect 8649 1957 8707 1969
rect 8649 -2019 8661 1957
rect 8695 -2019 8707 1957
rect 8649 -2031 8707 -2019
rect 8807 1957 8865 1969
rect 8807 -2019 8819 1957
rect 8853 -2019 8865 1957
rect 8807 -2031 8865 -2019
rect 8927 1957 8985 1969
rect 8927 -2019 8939 1957
rect 8973 -2019 8985 1957
rect 8927 -2031 8985 -2019
rect 9085 1957 9143 1969
rect 9085 -2019 9097 1957
rect 9131 -2019 9143 1957
rect 9085 -2031 9143 -2019
rect 9205 1957 9263 1969
rect 9205 -2019 9217 1957
rect 9251 -2019 9263 1957
rect 9205 -2031 9263 -2019
rect 9363 1957 9421 1969
rect 9363 -2019 9375 1957
rect 9409 -2019 9421 1957
rect 9363 -2031 9421 -2019
rect 9483 1957 9541 1969
rect 9483 -2019 9495 1957
rect 9529 -2019 9541 1957
rect 9483 -2031 9541 -2019
rect 9641 1957 9699 1969
rect 9641 -2019 9653 1957
rect 9687 -2019 9699 1957
rect 9641 -2031 9699 -2019
rect 9761 1957 9819 1969
rect 9761 -2019 9773 1957
rect 9807 -2019 9819 1957
rect 9761 -2031 9819 -2019
rect 9919 1957 9977 1969
rect 9919 -2019 9931 1957
rect 9965 -2019 9977 1957
rect 9919 -2031 9977 -2019
rect 10039 1957 10097 1969
rect 10039 -2019 10051 1957
rect 10085 -2019 10097 1957
rect 10039 -2031 10097 -2019
rect 10197 1957 10255 1969
rect 10197 -2019 10209 1957
rect 10243 -2019 10255 1957
rect 10197 -2031 10255 -2019
rect 10317 1957 10375 1969
rect 10317 -2019 10329 1957
rect 10363 -2019 10375 1957
rect 10317 -2031 10375 -2019
rect 10475 1957 10533 1969
rect 10475 -2019 10487 1957
rect 10521 -2019 10533 1957
rect 10475 -2031 10533 -2019
rect 10595 1957 10653 1969
rect 10595 -2019 10607 1957
rect 10641 -2019 10653 1957
rect 10595 -2031 10653 -2019
rect 10753 1957 10811 1969
rect 10753 -2019 10765 1957
rect 10799 -2019 10811 1957
rect 10753 -2031 10811 -2019
rect 10873 1957 10931 1969
rect 10873 -2019 10885 1957
rect 10919 -2019 10931 1957
rect 10873 -2031 10931 -2019
rect 11031 1957 11089 1969
rect 11031 -2019 11043 1957
rect 11077 -2019 11089 1957
rect 11031 -2031 11089 -2019
rect 11151 1957 11209 1969
rect 11151 -2019 11163 1957
rect 11197 -2019 11209 1957
rect 11151 -2031 11209 -2019
rect 11309 1957 11367 1969
rect 11309 -2019 11321 1957
rect 11355 -2019 11367 1957
rect 11309 -2031 11367 -2019
rect 11429 1957 11487 1969
rect 11429 -2019 11441 1957
rect 11475 -2019 11487 1957
rect 11429 -2031 11487 -2019
rect 11587 1957 11645 1969
rect 11587 -2019 11599 1957
rect 11633 -2019 11645 1957
rect 11587 -2031 11645 -2019
rect 11707 1957 11765 1969
rect 11707 -2019 11719 1957
rect 11753 -2019 11765 1957
rect 11707 -2031 11765 -2019
rect 11865 1957 11923 1969
rect 11865 -2019 11877 1957
rect 11911 -2019 11923 1957
rect 11865 -2031 11923 -2019
rect 11985 1957 12043 1969
rect 11985 -2019 11997 1957
rect 12031 -2019 12043 1957
rect 11985 -2031 12043 -2019
rect 12143 1957 12201 1969
rect 12143 -2019 12155 1957
rect 12189 -2019 12201 1957
rect 12143 -2031 12201 -2019
rect 12263 1957 12321 1969
rect 12263 -2019 12275 1957
rect 12309 -2019 12321 1957
rect 12263 -2031 12321 -2019
rect 12421 1957 12479 1969
rect 12421 -2019 12433 1957
rect 12467 -2019 12479 1957
rect 12421 -2031 12479 -2019
rect 12541 1957 12599 1969
rect 12541 -2019 12553 1957
rect 12587 -2019 12599 1957
rect 12541 -2031 12599 -2019
rect 12699 1957 12757 1969
rect 12699 -2019 12711 1957
rect 12745 -2019 12757 1957
rect 12699 -2031 12757 -2019
rect 12819 1957 12877 1969
rect 12819 -2019 12831 1957
rect 12865 -2019 12877 1957
rect 12819 -2031 12877 -2019
rect 12977 1957 13035 1969
rect 12977 -2019 12989 1957
rect 13023 -2019 13035 1957
rect 12977 -2031 13035 -2019
rect 13097 1957 13155 1969
rect 13097 -2019 13109 1957
rect 13143 -2019 13155 1957
rect 13097 -2031 13155 -2019
rect 13255 1957 13313 1969
rect 13255 -2019 13267 1957
rect 13301 -2019 13313 1957
rect 13255 -2031 13313 -2019
rect 13375 1957 13433 1969
rect 13375 -2019 13387 1957
rect 13421 -2019 13433 1957
rect 13375 -2031 13433 -2019
rect 13533 1957 13591 1969
rect 13533 -2019 13545 1957
rect 13579 -2019 13591 1957
rect 13533 -2031 13591 -2019
rect 13653 1957 13711 1969
rect 13653 -2019 13665 1957
rect 13699 -2019 13711 1957
rect 13653 -2031 13711 -2019
rect 13811 1957 13869 1969
rect 13811 -2019 13823 1957
rect 13857 -2019 13869 1957
rect 13811 -2031 13869 -2019
rect 13931 1957 13989 1969
rect 13931 -2019 13943 1957
rect 13977 -2019 13989 1957
rect 13931 -2031 13989 -2019
rect 14089 1957 14147 1969
rect 14089 -2019 14101 1957
rect 14135 -2019 14147 1957
rect 14089 -2031 14147 -2019
rect 14209 1957 14267 1969
rect 14209 -2019 14221 1957
rect 14255 -2019 14267 1957
rect 14209 -2031 14267 -2019
rect 14367 1957 14425 1969
rect 14367 -2019 14379 1957
rect 14413 -2019 14425 1957
rect 14367 -2031 14425 -2019
rect 14487 1957 14545 1969
rect 14487 -2019 14499 1957
rect 14533 -2019 14545 1957
rect 14487 -2031 14545 -2019
rect 14645 1957 14703 1969
rect 14645 -2019 14657 1957
rect 14691 -2019 14703 1957
rect 14645 -2031 14703 -2019
rect 14765 1957 14823 1969
rect 14765 -2019 14777 1957
rect 14811 -2019 14823 1957
rect 14765 -2031 14823 -2019
rect 14923 1957 14981 1969
rect 14923 -2019 14935 1957
rect 14969 -2019 14981 1957
rect 14923 -2031 14981 -2019
rect 15043 1957 15101 1969
rect 15043 -2019 15055 1957
rect 15089 -2019 15101 1957
rect 15043 -2031 15101 -2019
rect 15201 1957 15259 1969
rect 15201 -2019 15213 1957
rect 15247 -2019 15259 1957
rect 15201 -2031 15259 -2019
rect 15321 1957 15379 1969
rect 15321 -2019 15333 1957
rect 15367 -2019 15379 1957
rect 15321 -2031 15379 -2019
rect 15479 1957 15537 1969
rect 15479 -2019 15491 1957
rect 15525 -2019 15537 1957
rect 15479 -2031 15537 -2019
rect 15599 1957 15657 1969
rect 15599 -2019 15611 1957
rect 15645 -2019 15657 1957
rect 15599 -2031 15657 -2019
rect 15757 1957 15815 1969
rect 15757 -2019 15769 1957
rect 15803 -2019 15815 1957
rect 15757 -2031 15815 -2019
rect 15877 1957 15935 1969
rect 15877 -2019 15889 1957
rect 15923 -2019 15935 1957
rect 15877 -2031 15935 -2019
rect 16035 1957 16093 1969
rect 16035 -2019 16047 1957
rect 16081 -2019 16093 1957
rect 16035 -2031 16093 -2019
rect 16155 1957 16213 1969
rect 16155 -2019 16167 1957
rect 16201 -2019 16213 1957
rect 16155 -2031 16213 -2019
rect 16313 1957 16371 1969
rect 16313 -2019 16325 1957
rect 16359 -2019 16371 1957
rect 16313 -2031 16371 -2019
rect 16433 1957 16491 1969
rect 16433 -2019 16445 1957
rect 16479 -2019 16491 1957
rect 16433 -2031 16491 -2019
rect 16591 1957 16649 1969
rect 16591 -2019 16603 1957
rect 16637 -2019 16649 1957
rect 16591 -2031 16649 -2019
rect 16711 1957 16769 1969
rect 16711 -2019 16723 1957
rect 16757 -2019 16769 1957
rect 16711 -2031 16769 -2019
rect 16869 1957 16927 1969
rect 16869 -2019 16881 1957
rect 16915 -2019 16927 1957
rect 16869 -2031 16927 -2019
rect 16989 1957 17047 1969
rect 16989 -2019 17001 1957
rect 17035 -2019 17047 1957
rect 16989 -2031 17047 -2019
rect 17147 1957 17205 1969
rect 17147 -2019 17159 1957
rect 17193 -2019 17205 1957
rect 17147 -2031 17205 -2019
rect 17267 1957 17325 1969
rect 17267 -2019 17279 1957
rect 17313 -2019 17325 1957
rect 17267 -2031 17325 -2019
rect 17425 1957 17483 1969
rect 17425 -2019 17437 1957
rect 17471 -2019 17483 1957
rect 17425 -2031 17483 -2019
rect 17545 1957 17603 1969
rect 17545 -2019 17557 1957
rect 17591 -2019 17603 1957
rect 17545 -2031 17603 -2019
rect 17703 1957 17761 1969
rect 17703 -2019 17715 1957
rect 17749 -2019 17761 1957
rect 17703 -2031 17761 -2019
<< mvndiffc >>
rect -17749 -2019 -17715 1957
rect -17591 -2019 -17557 1957
rect -17471 -2019 -17437 1957
rect -17313 -2019 -17279 1957
rect -17193 -2019 -17159 1957
rect -17035 -2019 -17001 1957
rect -16915 -2019 -16881 1957
rect -16757 -2019 -16723 1957
rect -16637 -2019 -16603 1957
rect -16479 -2019 -16445 1957
rect -16359 -2019 -16325 1957
rect -16201 -2019 -16167 1957
rect -16081 -2019 -16047 1957
rect -15923 -2019 -15889 1957
rect -15803 -2019 -15769 1957
rect -15645 -2019 -15611 1957
rect -15525 -2019 -15491 1957
rect -15367 -2019 -15333 1957
rect -15247 -2019 -15213 1957
rect -15089 -2019 -15055 1957
rect -14969 -2019 -14935 1957
rect -14811 -2019 -14777 1957
rect -14691 -2019 -14657 1957
rect -14533 -2019 -14499 1957
rect -14413 -2019 -14379 1957
rect -14255 -2019 -14221 1957
rect -14135 -2019 -14101 1957
rect -13977 -2019 -13943 1957
rect -13857 -2019 -13823 1957
rect -13699 -2019 -13665 1957
rect -13579 -2019 -13545 1957
rect -13421 -2019 -13387 1957
rect -13301 -2019 -13267 1957
rect -13143 -2019 -13109 1957
rect -13023 -2019 -12989 1957
rect -12865 -2019 -12831 1957
rect -12745 -2019 -12711 1957
rect -12587 -2019 -12553 1957
rect -12467 -2019 -12433 1957
rect -12309 -2019 -12275 1957
rect -12189 -2019 -12155 1957
rect -12031 -2019 -11997 1957
rect -11911 -2019 -11877 1957
rect -11753 -2019 -11719 1957
rect -11633 -2019 -11599 1957
rect -11475 -2019 -11441 1957
rect -11355 -2019 -11321 1957
rect -11197 -2019 -11163 1957
rect -11077 -2019 -11043 1957
rect -10919 -2019 -10885 1957
rect -10799 -2019 -10765 1957
rect -10641 -2019 -10607 1957
rect -10521 -2019 -10487 1957
rect -10363 -2019 -10329 1957
rect -10243 -2019 -10209 1957
rect -10085 -2019 -10051 1957
rect -9965 -2019 -9931 1957
rect -9807 -2019 -9773 1957
rect -9687 -2019 -9653 1957
rect -9529 -2019 -9495 1957
rect -9409 -2019 -9375 1957
rect -9251 -2019 -9217 1957
rect -9131 -2019 -9097 1957
rect -8973 -2019 -8939 1957
rect -8853 -2019 -8819 1957
rect -8695 -2019 -8661 1957
rect -8575 -2019 -8541 1957
rect -8417 -2019 -8383 1957
rect -8297 -2019 -8263 1957
rect -8139 -2019 -8105 1957
rect -8019 -2019 -7985 1957
rect -7861 -2019 -7827 1957
rect -7741 -2019 -7707 1957
rect -7583 -2019 -7549 1957
rect -7463 -2019 -7429 1957
rect -7305 -2019 -7271 1957
rect -7185 -2019 -7151 1957
rect -7027 -2019 -6993 1957
rect -6907 -2019 -6873 1957
rect -6749 -2019 -6715 1957
rect -6629 -2019 -6595 1957
rect -6471 -2019 -6437 1957
rect -6351 -2019 -6317 1957
rect -6193 -2019 -6159 1957
rect -6073 -2019 -6039 1957
rect -5915 -2019 -5881 1957
rect -5795 -2019 -5761 1957
rect -5637 -2019 -5603 1957
rect -5517 -2019 -5483 1957
rect -5359 -2019 -5325 1957
rect -5239 -2019 -5205 1957
rect -5081 -2019 -5047 1957
rect -4961 -2019 -4927 1957
rect -4803 -2019 -4769 1957
rect -4683 -2019 -4649 1957
rect -4525 -2019 -4491 1957
rect -4405 -2019 -4371 1957
rect -4247 -2019 -4213 1957
rect -4127 -2019 -4093 1957
rect -3969 -2019 -3935 1957
rect -3849 -2019 -3815 1957
rect -3691 -2019 -3657 1957
rect -3571 -2019 -3537 1957
rect -3413 -2019 -3379 1957
rect -3293 -2019 -3259 1957
rect -3135 -2019 -3101 1957
rect -3015 -2019 -2981 1957
rect -2857 -2019 -2823 1957
rect -2737 -2019 -2703 1957
rect -2579 -2019 -2545 1957
rect -2459 -2019 -2425 1957
rect -2301 -2019 -2267 1957
rect -2181 -2019 -2147 1957
rect -2023 -2019 -1989 1957
rect -1903 -2019 -1869 1957
rect -1745 -2019 -1711 1957
rect -1625 -2019 -1591 1957
rect -1467 -2019 -1433 1957
rect -1347 -2019 -1313 1957
rect -1189 -2019 -1155 1957
rect -1069 -2019 -1035 1957
rect -911 -2019 -877 1957
rect -791 -2019 -757 1957
rect -633 -2019 -599 1957
rect -513 -2019 -479 1957
rect -355 -2019 -321 1957
rect -235 -2019 -201 1957
rect -77 -2019 -43 1957
rect 43 -2019 77 1957
rect 201 -2019 235 1957
rect 321 -2019 355 1957
rect 479 -2019 513 1957
rect 599 -2019 633 1957
rect 757 -2019 791 1957
rect 877 -2019 911 1957
rect 1035 -2019 1069 1957
rect 1155 -2019 1189 1957
rect 1313 -2019 1347 1957
rect 1433 -2019 1467 1957
rect 1591 -2019 1625 1957
rect 1711 -2019 1745 1957
rect 1869 -2019 1903 1957
rect 1989 -2019 2023 1957
rect 2147 -2019 2181 1957
rect 2267 -2019 2301 1957
rect 2425 -2019 2459 1957
rect 2545 -2019 2579 1957
rect 2703 -2019 2737 1957
rect 2823 -2019 2857 1957
rect 2981 -2019 3015 1957
rect 3101 -2019 3135 1957
rect 3259 -2019 3293 1957
rect 3379 -2019 3413 1957
rect 3537 -2019 3571 1957
rect 3657 -2019 3691 1957
rect 3815 -2019 3849 1957
rect 3935 -2019 3969 1957
rect 4093 -2019 4127 1957
rect 4213 -2019 4247 1957
rect 4371 -2019 4405 1957
rect 4491 -2019 4525 1957
rect 4649 -2019 4683 1957
rect 4769 -2019 4803 1957
rect 4927 -2019 4961 1957
rect 5047 -2019 5081 1957
rect 5205 -2019 5239 1957
rect 5325 -2019 5359 1957
rect 5483 -2019 5517 1957
rect 5603 -2019 5637 1957
rect 5761 -2019 5795 1957
rect 5881 -2019 5915 1957
rect 6039 -2019 6073 1957
rect 6159 -2019 6193 1957
rect 6317 -2019 6351 1957
rect 6437 -2019 6471 1957
rect 6595 -2019 6629 1957
rect 6715 -2019 6749 1957
rect 6873 -2019 6907 1957
rect 6993 -2019 7027 1957
rect 7151 -2019 7185 1957
rect 7271 -2019 7305 1957
rect 7429 -2019 7463 1957
rect 7549 -2019 7583 1957
rect 7707 -2019 7741 1957
rect 7827 -2019 7861 1957
rect 7985 -2019 8019 1957
rect 8105 -2019 8139 1957
rect 8263 -2019 8297 1957
rect 8383 -2019 8417 1957
rect 8541 -2019 8575 1957
rect 8661 -2019 8695 1957
rect 8819 -2019 8853 1957
rect 8939 -2019 8973 1957
rect 9097 -2019 9131 1957
rect 9217 -2019 9251 1957
rect 9375 -2019 9409 1957
rect 9495 -2019 9529 1957
rect 9653 -2019 9687 1957
rect 9773 -2019 9807 1957
rect 9931 -2019 9965 1957
rect 10051 -2019 10085 1957
rect 10209 -2019 10243 1957
rect 10329 -2019 10363 1957
rect 10487 -2019 10521 1957
rect 10607 -2019 10641 1957
rect 10765 -2019 10799 1957
rect 10885 -2019 10919 1957
rect 11043 -2019 11077 1957
rect 11163 -2019 11197 1957
rect 11321 -2019 11355 1957
rect 11441 -2019 11475 1957
rect 11599 -2019 11633 1957
rect 11719 -2019 11753 1957
rect 11877 -2019 11911 1957
rect 11997 -2019 12031 1957
rect 12155 -2019 12189 1957
rect 12275 -2019 12309 1957
rect 12433 -2019 12467 1957
rect 12553 -2019 12587 1957
rect 12711 -2019 12745 1957
rect 12831 -2019 12865 1957
rect 12989 -2019 13023 1957
rect 13109 -2019 13143 1957
rect 13267 -2019 13301 1957
rect 13387 -2019 13421 1957
rect 13545 -2019 13579 1957
rect 13665 -2019 13699 1957
rect 13823 -2019 13857 1957
rect 13943 -2019 13977 1957
rect 14101 -2019 14135 1957
rect 14221 -2019 14255 1957
rect 14379 -2019 14413 1957
rect 14499 -2019 14533 1957
rect 14657 -2019 14691 1957
rect 14777 -2019 14811 1957
rect 14935 -2019 14969 1957
rect 15055 -2019 15089 1957
rect 15213 -2019 15247 1957
rect 15333 -2019 15367 1957
rect 15491 -2019 15525 1957
rect 15611 -2019 15645 1957
rect 15769 -2019 15803 1957
rect 15889 -2019 15923 1957
rect 16047 -2019 16081 1957
rect 16167 -2019 16201 1957
rect 16325 -2019 16359 1957
rect 16445 -2019 16479 1957
rect 16603 -2019 16637 1957
rect 16723 -2019 16757 1957
rect 16881 -2019 16915 1957
rect 17001 -2019 17035 1957
rect 17159 -2019 17193 1957
rect 17279 -2019 17313 1957
rect 17437 -2019 17471 1957
rect 17557 -2019 17591 1957
rect 17715 -2019 17749 1957
<< poly >>
rect -17703 2041 -17603 2057
rect -17703 2007 -17687 2041
rect -17619 2007 -17603 2041
rect -17703 1969 -17603 2007
rect -17425 2041 -17325 2057
rect -17425 2007 -17409 2041
rect -17341 2007 -17325 2041
rect -17425 1969 -17325 2007
rect -17147 2041 -17047 2057
rect -17147 2007 -17131 2041
rect -17063 2007 -17047 2041
rect -17147 1969 -17047 2007
rect -16869 2041 -16769 2057
rect -16869 2007 -16853 2041
rect -16785 2007 -16769 2041
rect -16869 1969 -16769 2007
rect -16591 2041 -16491 2057
rect -16591 2007 -16575 2041
rect -16507 2007 -16491 2041
rect -16591 1969 -16491 2007
rect -16313 2041 -16213 2057
rect -16313 2007 -16297 2041
rect -16229 2007 -16213 2041
rect -16313 1969 -16213 2007
rect -16035 2041 -15935 2057
rect -16035 2007 -16019 2041
rect -15951 2007 -15935 2041
rect -16035 1969 -15935 2007
rect -15757 2041 -15657 2057
rect -15757 2007 -15741 2041
rect -15673 2007 -15657 2041
rect -15757 1969 -15657 2007
rect -15479 2041 -15379 2057
rect -15479 2007 -15463 2041
rect -15395 2007 -15379 2041
rect -15479 1969 -15379 2007
rect -15201 2041 -15101 2057
rect -15201 2007 -15185 2041
rect -15117 2007 -15101 2041
rect -15201 1969 -15101 2007
rect -14923 2041 -14823 2057
rect -14923 2007 -14907 2041
rect -14839 2007 -14823 2041
rect -14923 1969 -14823 2007
rect -14645 2041 -14545 2057
rect -14645 2007 -14629 2041
rect -14561 2007 -14545 2041
rect -14645 1969 -14545 2007
rect -14367 2041 -14267 2057
rect -14367 2007 -14351 2041
rect -14283 2007 -14267 2041
rect -14367 1969 -14267 2007
rect -14089 2041 -13989 2057
rect -14089 2007 -14073 2041
rect -14005 2007 -13989 2041
rect -14089 1969 -13989 2007
rect -13811 2041 -13711 2057
rect -13811 2007 -13795 2041
rect -13727 2007 -13711 2041
rect -13811 1969 -13711 2007
rect -13533 2041 -13433 2057
rect -13533 2007 -13517 2041
rect -13449 2007 -13433 2041
rect -13533 1969 -13433 2007
rect -13255 2041 -13155 2057
rect -13255 2007 -13239 2041
rect -13171 2007 -13155 2041
rect -13255 1969 -13155 2007
rect -12977 2041 -12877 2057
rect -12977 2007 -12961 2041
rect -12893 2007 -12877 2041
rect -12977 1969 -12877 2007
rect -12699 2041 -12599 2057
rect -12699 2007 -12683 2041
rect -12615 2007 -12599 2041
rect -12699 1969 -12599 2007
rect -12421 2041 -12321 2057
rect -12421 2007 -12405 2041
rect -12337 2007 -12321 2041
rect -12421 1969 -12321 2007
rect -12143 2041 -12043 2057
rect -12143 2007 -12127 2041
rect -12059 2007 -12043 2041
rect -12143 1969 -12043 2007
rect -11865 2041 -11765 2057
rect -11865 2007 -11849 2041
rect -11781 2007 -11765 2041
rect -11865 1969 -11765 2007
rect -11587 2041 -11487 2057
rect -11587 2007 -11571 2041
rect -11503 2007 -11487 2041
rect -11587 1969 -11487 2007
rect -11309 2041 -11209 2057
rect -11309 2007 -11293 2041
rect -11225 2007 -11209 2041
rect -11309 1969 -11209 2007
rect -11031 2041 -10931 2057
rect -11031 2007 -11015 2041
rect -10947 2007 -10931 2041
rect -11031 1969 -10931 2007
rect -10753 2041 -10653 2057
rect -10753 2007 -10737 2041
rect -10669 2007 -10653 2041
rect -10753 1969 -10653 2007
rect -10475 2041 -10375 2057
rect -10475 2007 -10459 2041
rect -10391 2007 -10375 2041
rect -10475 1969 -10375 2007
rect -10197 2041 -10097 2057
rect -10197 2007 -10181 2041
rect -10113 2007 -10097 2041
rect -10197 1969 -10097 2007
rect -9919 2041 -9819 2057
rect -9919 2007 -9903 2041
rect -9835 2007 -9819 2041
rect -9919 1969 -9819 2007
rect -9641 2041 -9541 2057
rect -9641 2007 -9625 2041
rect -9557 2007 -9541 2041
rect -9641 1969 -9541 2007
rect -9363 2041 -9263 2057
rect -9363 2007 -9347 2041
rect -9279 2007 -9263 2041
rect -9363 1969 -9263 2007
rect -9085 2041 -8985 2057
rect -9085 2007 -9069 2041
rect -9001 2007 -8985 2041
rect -9085 1969 -8985 2007
rect -8807 2041 -8707 2057
rect -8807 2007 -8791 2041
rect -8723 2007 -8707 2041
rect -8807 1969 -8707 2007
rect -8529 2041 -8429 2057
rect -8529 2007 -8513 2041
rect -8445 2007 -8429 2041
rect -8529 1969 -8429 2007
rect -8251 2041 -8151 2057
rect -8251 2007 -8235 2041
rect -8167 2007 -8151 2041
rect -8251 1969 -8151 2007
rect -7973 2041 -7873 2057
rect -7973 2007 -7957 2041
rect -7889 2007 -7873 2041
rect -7973 1969 -7873 2007
rect -7695 2041 -7595 2057
rect -7695 2007 -7679 2041
rect -7611 2007 -7595 2041
rect -7695 1969 -7595 2007
rect -7417 2041 -7317 2057
rect -7417 2007 -7401 2041
rect -7333 2007 -7317 2041
rect -7417 1969 -7317 2007
rect -7139 2041 -7039 2057
rect -7139 2007 -7123 2041
rect -7055 2007 -7039 2041
rect -7139 1969 -7039 2007
rect -6861 2041 -6761 2057
rect -6861 2007 -6845 2041
rect -6777 2007 -6761 2041
rect -6861 1969 -6761 2007
rect -6583 2041 -6483 2057
rect -6583 2007 -6567 2041
rect -6499 2007 -6483 2041
rect -6583 1969 -6483 2007
rect -6305 2041 -6205 2057
rect -6305 2007 -6289 2041
rect -6221 2007 -6205 2041
rect -6305 1969 -6205 2007
rect -6027 2041 -5927 2057
rect -6027 2007 -6011 2041
rect -5943 2007 -5927 2041
rect -6027 1969 -5927 2007
rect -5749 2041 -5649 2057
rect -5749 2007 -5733 2041
rect -5665 2007 -5649 2041
rect -5749 1969 -5649 2007
rect -5471 2041 -5371 2057
rect -5471 2007 -5455 2041
rect -5387 2007 -5371 2041
rect -5471 1969 -5371 2007
rect -5193 2041 -5093 2057
rect -5193 2007 -5177 2041
rect -5109 2007 -5093 2041
rect -5193 1969 -5093 2007
rect -4915 2041 -4815 2057
rect -4915 2007 -4899 2041
rect -4831 2007 -4815 2041
rect -4915 1969 -4815 2007
rect -4637 2041 -4537 2057
rect -4637 2007 -4621 2041
rect -4553 2007 -4537 2041
rect -4637 1969 -4537 2007
rect -4359 2041 -4259 2057
rect -4359 2007 -4343 2041
rect -4275 2007 -4259 2041
rect -4359 1969 -4259 2007
rect -4081 2041 -3981 2057
rect -4081 2007 -4065 2041
rect -3997 2007 -3981 2041
rect -4081 1969 -3981 2007
rect -3803 2041 -3703 2057
rect -3803 2007 -3787 2041
rect -3719 2007 -3703 2041
rect -3803 1969 -3703 2007
rect -3525 2041 -3425 2057
rect -3525 2007 -3509 2041
rect -3441 2007 -3425 2041
rect -3525 1969 -3425 2007
rect -3247 2041 -3147 2057
rect -3247 2007 -3231 2041
rect -3163 2007 -3147 2041
rect -3247 1969 -3147 2007
rect -2969 2041 -2869 2057
rect -2969 2007 -2953 2041
rect -2885 2007 -2869 2041
rect -2969 1969 -2869 2007
rect -2691 2041 -2591 2057
rect -2691 2007 -2675 2041
rect -2607 2007 -2591 2041
rect -2691 1969 -2591 2007
rect -2413 2041 -2313 2057
rect -2413 2007 -2397 2041
rect -2329 2007 -2313 2041
rect -2413 1969 -2313 2007
rect -2135 2041 -2035 2057
rect -2135 2007 -2119 2041
rect -2051 2007 -2035 2041
rect -2135 1969 -2035 2007
rect -1857 2041 -1757 2057
rect -1857 2007 -1841 2041
rect -1773 2007 -1757 2041
rect -1857 1969 -1757 2007
rect -1579 2041 -1479 2057
rect -1579 2007 -1563 2041
rect -1495 2007 -1479 2041
rect -1579 1969 -1479 2007
rect -1301 2041 -1201 2057
rect -1301 2007 -1285 2041
rect -1217 2007 -1201 2041
rect -1301 1969 -1201 2007
rect -1023 2041 -923 2057
rect -1023 2007 -1007 2041
rect -939 2007 -923 2041
rect -1023 1969 -923 2007
rect -745 2041 -645 2057
rect -745 2007 -729 2041
rect -661 2007 -645 2041
rect -745 1969 -645 2007
rect -467 2041 -367 2057
rect -467 2007 -451 2041
rect -383 2007 -367 2041
rect -467 1969 -367 2007
rect -189 2041 -89 2057
rect -189 2007 -173 2041
rect -105 2007 -89 2041
rect -189 1969 -89 2007
rect 89 2041 189 2057
rect 89 2007 105 2041
rect 173 2007 189 2041
rect 89 1969 189 2007
rect 367 2041 467 2057
rect 367 2007 383 2041
rect 451 2007 467 2041
rect 367 1969 467 2007
rect 645 2041 745 2057
rect 645 2007 661 2041
rect 729 2007 745 2041
rect 645 1969 745 2007
rect 923 2041 1023 2057
rect 923 2007 939 2041
rect 1007 2007 1023 2041
rect 923 1969 1023 2007
rect 1201 2041 1301 2057
rect 1201 2007 1217 2041
rect 1285 2007 1301 2041
rect 1201 1969 1301 2007
rect 1479 2041 1579 2057
rect 1479 2007 1495 2041
rect 1563 2007 1579 2041
rect 1479 1969 1579 2007
rect 1757 2041 1857 2057
rect 1757 2007 1773 2041
rect 1841 2007 1857 2041
rect 1757 1969 1857 2007
rect 2035 2041 2135 2057
rect 2035 2007 2051 2041
rect 2119 2007 2135 2041
rect 2035 1969 2135 2007
rect 2313 2041 2413 2057
rect 2313 2007 2329 2041
rect 2397 2007 2413 2041
rect 2313 1969 2413 2007
rect 2591 2041 2691 2057
rect 2591 2007 2607 2041
rect 2675 2007 2691 2041
rect 2591 1969 2691 2007
rect 2869 2041 2969 2057
rect 2869 2007 2885 2041
rect 2953 2007 2969 2041
rect 2869 1969 2969 2007
rect 3147 2041 3247 2057
rect 3147 2007 3163 2041
rect 3231 2007 3247 2041
rect 3147 1969 3247 2007
rect 3425 2041 3525 2057
rect 3425 2007 3441 2041
rect 3509 2007 3525 2041
rect 3425 1969 3525 2007
rect 3703 2041 3803 2057
rect 3703 2007 3719 2041
rect 3787 2007 3803 2041
rect 3703 1969 3803 2007
rect 3981 2041 4081 2057
rect 3981 2007 3997 2041
rect 4065 2007 4081 2041
rect 3981 1969 4081 2007
rect 4259 2041 4359 2057
rect 4259 2007 4275 2041
rect 4343 2007 4359 2041
rect 4259 1969 4359 2007
rect 4537 2041 4637 2057
rect 4537 2007 4553 2041
rect 4621 2007 4637 2041
rect 4537 1969 4637 2007
rect 4815 2041 4915 2057
rect 4815 2007 4831 2041
rect 4899 2007 4915 2041
rect 4815 1969 4915 2007
rect 5093 2041 5193 2057
rect 5093 2007 5109 2041
rect 5177 2007 5193 2041
rect 5093 1969 5193 2007
rect 5371 2041 5471 2057
rect 5371 2007 5387 2041
rect 5455 2007 5471 2041
rect 5371 1969 5471 2007
rect 5649 2041 5749 2057
rect 5649 2007 5665 2041
rect 5733 2007 5749 2041
rect 5649 1969 5749 2007
rect 5927 2041 6027 2057
rect 5927 2007 5943 2041
rect 6011 2007 6027 2041
rect 5927 1969 6027 2007
rect 6205 2041 6305 2057
rect 6205 2007 6221 2041
rect 6289 2007 6305 2041
rect 6205 1969 6305 2007
rect 6483 2041 6583 2057
rect 6483 2007 6499 2041
rect 6567 2007 6583 2041
rect 6483 1969 6583 2007
rect 6761 2041 6861 2057
rect 6761 2007 6777 2041
rect 6845 2007 6861 2041
rect 6761 1969 6861 2007
rect 7039 2041 7139 2057
rect 7039 2007 7055 2041
rect 7123 2007 7139 2041
rect 7039 1969 7139 2007
rect 7317 2041 7417 2057
rect 7317 2007 7333 2041
rect 7401 2007 7417 2041
rect 7317 1969 7417 2007
rect 7595 2041 7695 2057
rect 7595 2007 7611 2041
rect 7679 2007 7695 2041
rect 7595 1969 7695 2007
rect 7873 2041 7973 2057
rect 7873 2007 7889 2041
rect 7957 2007 7973 2041
rect 7873 1969 7973 2007
rect 8151 2041 8251 2057
rect 8151 2007 8167 2041
rect 8235 2007 8251 2041
rect 8151 1969 8251 2007
rect 8429 2041 8529 2057
rect 8429 2007 8445 2041
rect 8513 2007 8529 2041
rect 8429 1969 8529 2007
rect 8707 2041 8807 2057
rect 8707 2007 8723 2041
rect 8791 2007 8807 2041
rect 8707 1969 8807 2007
rect 8985 2041 9085 2057
rect 8985 2007 9001 2041
rect 9069 2007 9085 2041
rect 8985 1969 9085 2007
rect 9263 2041 9363 2057
rect 9263 2007 9279 2041
rect 9347 2007 9363 2041
rect 9263 1969 9363 2007
rect 9541 2041 9641 2057
rect 9541 2007 9557 2041
rect 9625 2007 9641 2041
rect 9541 1969 9641 2007
rect 9819 2041 9919 2057
rect 9819 2007 9835 2041
rect 9903 2007 9919 2041
rect 9819 1969 9919 2007
rect 10097 2041 10197 2057
rect 10097 2007 10113 2041
rect 10181 2007 10197 2041
rect 10097 1969 10197 2007
rect 10375 2041 10475 2057
rect 10375 2007 10391 2041
rect 10459 2007 10475 2041
rect 10375 1969 10475 2007
rect 10653 2041 10753 2057
rect 10653 2007 10669 2041
rect 10737 2007 10753 2041
rect 10653 1969 10753 2007
rect 10931 2041 11031 2057
rect 10931 2007 10947 2041
rect 11015 2007 11031 2041
rect 10931 1969 11031 2007
rect 11209 2041 11309 2057
rect 11209 2007 11225 2041
rect 11293 2007 11309 2041
rect 11209 1969 11309 2007
rect 11487 2041 11587 2057
rect 11487 2007 11503 2041
rect 11571 2007 11587 2041
rect 11487 1969 11587 2007
rect 11765 2041 11865 2057
rect 11765 2007 11781 2041
rect 11849 2007 11865 2041
rect 11765 1969 11865 2007
rect 12043 2041 12143 2057
rect 12043 2007 12059 2041
rect 12127 2007 12143 2041
rect 12043 1969 12143 2007
rect 12321 2041 12421 2057
rect 12321 2007 12337 2041
rect 12405 2007 12421 2041
rect 12321 1969 12421 2007
rect 12599 2041 12699 2057
rect 12599 2007 12615 2041
rect 12683 2007 12699 2041
rect 12599 1969 12699 2007
rect 12877 2041 12977 2057
rect 12877 2007 12893 2041
rect 12961 2007 12977 2041
rect 12877 1969 12977 2007
rect 13155 2041 13255 2057
rect 13155 2007 13171 2041
rect 13239 2007 13255 2041
rect 13155 1969 13255 2007
rect 13433 2041 13533 2057
rect 13433 2007 13449 2041
rect 13517 2007 13533 2041
rect 13433 1969 13533 2007
rect 13711 2041 13811 2057
rect 13711 2007 13727 2041
rect 13795 2007 13811 2041
rect 13711 1969 13811 2007
rect 13989 2041 14089 2057
rect 13989 2007 14005 2041
rect 14073 2007 14089 2041
rect 13989 1969 14089 2007
rect 14267 2041 14367 2057
rect 14267 2007 14283 2041
rect 14351 2007 14367 2041
rect 14267 1969 14367 2007
rect 14545 2041 14645 2057
rect 14545 2007 14561 2041
rect 14629 2007 14645 2041
rect 14545 1969 14645 2007
rect 14823 2041 14923 2057
rect 14823 2007 14839 2041
rect 14907 2007 14923 2041
rect 14823 1969 14923 2007
rect 15101 2041 15201 2057
rect 15101 2007 15117 2041
rect 15185 2007 15201 2041
rect 15101 1969 15201 2007
rect 15379 2041 15479 2057
rect 15379 2007 15395 2041
rect 15463 2007 15479 2041
rect 15379 1969 15479 2007
rect 15657 2041 15757 2057
rect 15657 2007 15673 2041
rect 15741 2007 15757 2041
rect 15657 1969 15757 2007
rect 15935 2041 16035 2057
rect 15935 2007 15951 2041
rect 16019 2007 16035 2041
rect 15935 1969 16035 2007
rect 16213 2041 16313 2057
rect 16213 2007 16229 2041
rect 16297 2007 16313 2041
rect 16213 1969 16313 2007
rect 16491 2041 16591 2057
rect 16491 2007 16507 2041
rect 16575 2007 16591 2041
rect 16491 1969 16591 2007
rect 16769 2041 16869 2057
rect 16769 2007 16785 2041
rect 16853 2007 16869 2041
rect 16769 1969 16869 2007
rect 17047 2041 17147 2057
rect 17047 2007 17063 2041
rect 17131 2007 17147 2041
rect 17047 1969 17147 2007
rect 17325 2041 17425 2057
rect 17325 2007 17341 2041
rect 17409 2007 17425 2041
rect 17325 1969 17425 2007
rect 17603 2041 17703 2057
rect 17603 2007 17619 2041
rect 17687 2007 17703 2041
rect 17603 1969 17703 2007
rect -17703 -2057 -17603 -2031
rect -17425 -2057 -17325 -2031
rect -17147 -2057 -17047 -2031
rect -16869 -2057 -16769 -2031
rect -16591 -2057 -16491 -2031
rect -16313 -2057 -16213 -2031
rect -16035 -2057 -15935 -2031
rect -15757 -2057 -15657 -2031
rect -15479 -2057 -15379 -2031
rect -15201 -2057 -15101 -2031
rect -14923 -2057 -14823 -2031
rect -14645 -2057 -14545 -2031
rect -14367 -2057 -14267 -2031
rect -14089 -2057 -13989 -2031
rect -13811 -2057 -13711 -2031
rect -13533 -2057 -13433 -2031
rect -13255 -2057 -13155 -2031
rect -12977 -2057 -12877 -2031
rect -12699 -2057 -12599 -2031
rect -12421 -2057 -12321 -2031
rect -12143 -2057 -12043 -2031
rect -11865 -2057 -11765 -2031
rect -11587 -2057 -11487 -2031
rect -11309 -2057 -11209 -2031
rect -11031 -2057 -10931 -2031
rect -10753 -2057 -10653 -2031
rect -10475 -2057 -10375 -2031
rect -10197 -2057 -10097 -2031
rect -9919 -2057 -9819 -2031
rect -9641 -2057 -9541 -2031
rect -9363 -2057 -9263 -2031
rect -9085 -2057 -8985 -2031
rect -8807 -2057 -8707 -2031
rect -8529 -2057 -8429 -2031
rect -8251 -2057 -8151 -2031
rect -7973 -2057 -7873 -2031
rect -7695 -2057 -7595 -2031
rect -7417 -2057 -7317 -2031
rect -7139 -2057 -7039 -2031
rect -6861 -2057 -6761 -2031
rect -6583 -2057 -6483 -2031
rect -6305 -2057 -6205 -2031
rect -6027 -2057 -5927 -2031
rect -5749 -2057 -5649 -2031
rect -5471 -2057 -5371 -2031
rect -5193 -2057 -5093 -2031
rect -4915 -2057 -4815 -2031
rect -4637 -2057 -4537 -2031
rect -4359 -2057 -4259 -2031
rect -4081 -2057 -3981 -2031
rect -3803 -2057 -3703 -2031
rect -3525 -2057 -3425 -2031
rect -3247 -2057 -3147 -2031
rect -2969 -2057 -2869 -2031
rect -2691 -2057 -2591 -2031
rect -2413 -2057 -2313 -2031
rect -2135 -2057 -2035 -2031
rect -1857 -2057 -1757 -2031
rect -1579 -2057 -1479 -2031
rect -1301 -2057 -1201 -2031
rect -1023 -2057 -923 -2031
rect -745 -2057 -645 -2031
rect -467 -2057 -367 -2031
rect -189 -2057 -89 -2031
rect 89 -2057 189 -2031
rect 367 -2057 467 -2031
rect 645 -2057 745 -2031
rect 923 -2057 1023 -2031
rect 1201 -2057 1301 -2031
rect 1479 -2057 1579 -2031
rect 1757 -2057 1857 -2031
rect 2035 -2057 2135 -2031
rect 2313 -2057 2413 -2031
rect 2591 -2057 2691 -2031
rect 2869 -2057 2969 -2031
rect 3147 -2057 3247 -2031
rect 3425 -2057 3525 -2031
rect 3703 -2057 3803 -2031
rect 3981 -2057 4081 -2031
rect 4259 -2057 4359 -2031
rect 4537 -2057 4637 -2031
rect 4815 -2057 4915 -2031
rect 5093 -2057 5193 -2031
rect 5371 -2057 5471 -2031
rect 5649 -2057 5749 -2031
rect 5927 -2057 6027 -2031
rect 6205 -2057 6305 -2031
rect 6483 -2057 6583 -2031
rect 6761 -2057 6861 -2031
rect 7039 -2057 7139 -2031
rect 7317 -2057 7417 -2031
rect 7595 -2057 7695 -2031
rect 7873 -2057 7973 -2031
rect 8151 -2057 8251 -2031
rect 8429 -2057 8529 -2031
rect 8707 -2057 8807 -2031
rect 8985 -2057 9085 -2031
rect 9263 -2057 9363 -2031
rect 9541 -2057 9641 -2031
rect 9819 -2057 9919 -2031
rect 10097 -2057 10197 -2031
rect 10375 -2057 10475 -2031
rect 10653 -2057 10753 -2031
rect 10931 -2057 11031 -2031
rect 11209 -2057 11309 -2031
rect 11487 -2057 11587 -2031
rect 11765 -2057 11865 -2031
rect 12043 -2057 12143 -2031
rect 12321 -2057 12421 -2031
rect 12599 -2057 12699 -2031
rect 12877 -2057 12977 -2031
rect 13155 -2057 13255 -2031
rect 13433 -2057 13533 -2031
rect 13711 -2057 13811 -2031
rect 13989 -2057 14089 -2031
rect 14267 -2057 14367 -2031
rect 14545 -2057 14645 -2031
rect 14823 -2057 14923 -2031
rect 15101 -2057 15201 -2031
rect 15379 -2057 15479 -2031
rect 15657 -2057 15757 -2031
rect 15935 -2057 16035 -2031
rect 16213 -2057 16313 -2031
rect 16491 -2057 16591 -2031
rect 16769 -2057 16869 -2031
rect 17047 -2057 17147 -2031
rect 17325 -2057 17425 -2031
rect 17603 -2057 17703 -2031
<< polycont >>
rect -17687 2007 -17619 2041
rect -17409 2007 -17341 2041
rect -17131 2007 -17063 2041
rect -16853 2007 -16785 2041
rect -16575 2007 -16507 2041
rect -16297 2007 -16229 2041
rect -16019 2007 -15951 2041
rect -15741 2007 -15673 2041
rect -15463 2007 -15395 2041
rect -15185 2007 -15117 2041
rect -14907 2007 -14839 2041
rect -14629 2007 -14561 2041
rect -14351 2007 -14283 2041
rect -14073 2007 -14005 2041
rect -13795 2007 -13727 2041
rect -13517 2007 -13449 2041
rect -13239 2007 -13171 2041
rect -12961 2007 -12893 2041
rect -12683 2007 -12615 2041
rect -12405 2007 -12337 2041
rect -12127 2007 -12059 2041
rect -11849 2007 -11781 2041
rect -11571 2007 -11503 2041
rect -11293 2007 -11225 2041
rect -11015 2007 -10947 2041
rect -10737 2007 -10669 2041
rect -10459 2007 -10391 2041
rect -10181 2007 -10113 2041
rect -9903 2007 -9835 2041
rect -9625 2007 -9557 2041
rect -9347 2007 -9279 2041
rect -9069 2007 -9001 2041
rect -8791 2007 -8723 2041
rect -8513 2007 -8445 2041
rect -8235 2007 -8167 2041
rect -7957 2007 -7889 2041
rect -7679 2007 -7611 2041
rect -7401 2007 -7333 2041
rect -7123 2007 -7055 2041
rect -6845 2007 -6777 2041
rect -6567 2007 -6499 2041
rect -6289 2007 -6221 2041
rect -6011 2007 -5943 2041
rect -5733 2007 -5665 2041
rect -5455 2007 -5387 2041
rect -5177 2007 -5109 2041
rect -4899 2007 -4831 2041
rect -4621 2007 -4553 2041
rect -4343 2007 -4275 2041
rect -4065 2007 -3997 2041
rect -3787 2007 -3719 2041
rect -3509 2007 -3441 2041
rect -3231 2007 -3163 2041
rect -2953 2007 -2885 2041
rect -2675 2007 -2607 2041
rect -2397 2007 -2329 2041
rect -2119 2007 -2051 2041
rect -1841 2007 -1773 2041
rect -1563 2007 -1495 2041
rect -1285 2007 -1217 2041
rect -1007 2007 -939 2041
rect -729 2007 -661 2041
rect -451 2007 -383 2041
rect -173 2007 -105 2041
rect 105 2007 173 2041
rect 383 2007 451 2041
rect 661 2007 729 2041
rect 939 2007 1007 2041
rect 1217 2007 1285 2041
rect 1495 2007 1563 2041
rect 1773 2007 1841 2041
rect 2051 2007 2119 2041
rect 2329 2007 2397 2041
rect 2607 2007 2675 2041
rect 2885 2007 2953 2041
rect 3163 2007 3231 2041
rect 3441 2007 3509 2041
rect 3719 2007 3787 2041
rect 3997 2007 4065 2041
rect 4275 2007 4343 2041
rect 4553 2007 4621 2041
rect 4831 2007 4899 2041
rect 5109 2007 5177 2041
rect 5387 2007 5455 2041
rect 5665 2007 5733 2041
rect 5943 2007 6011 2041
rect 6221 2007 6289 2041
rect 6499 2007 6567 2041
rect 6777 2007 6845 2041
rect 7055 2007 7123 2041
rect 7333 2007 7401 2041
rect 7611 2007 7679 2041
rect 7889 2007 7957 2041
rect 8167 2007 8235 2041
rect 8445 2007 8513 2041
rect 8723 2007 8791 2041
rect 9001 2007 9069 2041
rect 9279 2007 9347 2041
rect 9557 2007 9625 2041
rect 9835 2007 9903 2041
rect 10113 2007 10181 2041
rect 10391 2007 10459 2041
rect 10669 2007 10737 2041
rect 10947 2007 11015 2041
rect 11225 2007 11293 2041
rect 11503 2007 11571 2041
rect 11781 2007 11849 2041
rect 12059 2007 12127 2041
rect 12337 2007 12405 2041
rect 12615 2007 12683 2041
rect 12893 2007 12961 2041
rect 13171 2007 13239 2041
rect 13449 2007 13517 2041
rect 13727 2007 13795 2041
rect 14005 2007 14073 2041
rect 14283 2007 14351 2041
rect 14561 2007 14629 2041
rect 14839 2007 14907 2041
rect 15117 2007 15185 2041
rect 15395 2007 15463 2041
rect 15673 2007 15741 2041
rect 15951 2007 16019 2041
rect 16229 2007 16297 2041
rect 16507 2007 16575 2041
rect 16785 2007 16853 2041
rect 17063 2007 17131 2041
rect 17341 2007 17409 2041
rect 17619 2007 17687 2041
<< locali >>
rect -17703 2007 -17687 2041
rect -17619 2007 -17603 2041
rect -17425 2007 -17409 2041
rect -17341 2007 -17325 2041
rect -17147 2007 -17131 2041
rect -17063 2007 -17047 2041
rect -16869 2007 -16853 2041
rect -16785 2007 -16769 2041
rect -16591 2007 -16575 2041
rect -16507 2007 -16491 2041
rect -16313 2007 -16297 2041
rect -16229 2007 -16213 2041
rect -16035 2007 -16019 2041
rect -15951 2007 -15935 2041
rect -15757 2007 -15741 2041
rect -15673 2007 -15657 2041
rect -15479 2007 -15463 2041
rect -15395 2007 -15379 2041
rect -15201 2007 -15185 2041
rect -15117 2007 -15101 2041
rect -14923 2007 -14907 2041
rect -14839 2007 -14823 2041
rect -14645 2007 -14629 2041
rect -14561 2007 -14545 2041
rect -14367 2007 -14351 2041
rect -14283 2007 -14267 2041
rect -14089 2007 -14073 2041
rect -14005 2007 -13989 2041
rect -13811 2007 -13795 2041
rect -13727 2007 -13711 2041
rect -13533 2007 -13517 2041
rect -13449 2007 -13433 2041
rect -13255 2007 -13239 2041
rect -13171 2007 -13155 2041
rect -12977 2007 -12961 2041
rect -12893 2007 -12877 2041
rect -12699 2007 -12683 2041
rect -12615 2007 -12599 2041
rect -12421 2007 -12405 2041
rect -12337 2007 -12321 2041
rect -12143 2007 -12127 2041
rect -12059 2007 -12043 2041
rect -11865 2007 -11849 2041
rect -11781 2007 -11765 2041
rect -11587 2007 -11571 2041
rect -11503 2007 -11487 2041
rect -11309 2007 -11293 2041
rect -11225 2007 -11209 2041
rect -11031 2007 -11015 2041
rect -10947 2007 -10931 2041
rect -10753 2007 -10737 2041
rect -10669 2007 -10653 2041
rect -10475 2007 -10459 2041
rect -10391 2007 -10375 2041
rect -10197 2007 -10181 2041
rect -10113 2007 -10097 2041
rect -9919 2007 -9903 2041
rect -9835 2007 -9819 2041
rect -9641 2007 -9625 2041
rect -9557 2007 -9541 2041
rect -9363 2007 -9347 2041
rect -9279 2007 -9263 2041
rect -9085 2007 -9069 2041
rect -9001 2007 -8985 2041
rect -8807 2007 -8791 2041
rect -8723 2007 -8707 2041
rect -8529 2007 -8513 2041
rect -8445 2007 -8429 2041
rect -8251 2007 -8235 2041
rect -8167 2007 -8151 2041
rect -7973 2007 -7957 2041
rect -7889 2007 -7873 2041
rect -7695 2007 -7679 2041
rect -7611 2007 -7595 2041
rect -7417 2007 -7401 2041
rect -7333 2007 -7317 2041
rect -7139 2007 -7123 2041
rect -7055 2007 -7039 2041
rect -6861 2007 -6845 2041
rect -6777 2007 -6761 2041
rect -6583 2007 -6567 2041
rect -6499 2007 -6483 2041
rect -6305 2007 -6289 2041
rect -6221 2007 -6205 2041
rect -6027 2007 -6011 2041
rect -5943 2007 -5927 2041
rect -5749 2007 -5733 2041
rect -5665 2007 -5649 2041
rect -5471 2007 -5455 2041
rect -5387 2007 -5371 2041
rect -5193 2007 -5177 2041
rect -5109 2007 -5093 2041
rect -4915 2007 -4899 2041
rect -4831 2007 -4815 2041
rect -4637 2007 -4621 2041
rect -4553 2007 -4537 2041
rect -4359 2007 -4343 2041
rect -4275 2007 -4259 2041
rect -4081 2007 -4065 2041
rect -3997 2007 -3981 2041
rect -3803 2007 -3787 2041
rect -3719 2007 -3703 2041
rect -3525 2007 -3509 2041
rect -3441 2007 -3425 2041
rect -3247 2007 -3231 2041
rect -3163 2007 -3147 2041
rect -2969 2007 -2953 2041
rect -2885 2007 -2869 2041
rect -2691 2007 -2675 2041
rect -2607 2007 -2591 2041
rect -2413 2007 -2397 2041
rect -2329 2007 -2313 2041
rect -2135 2007 -2119 2041
rect -2051 2007 -2035 2041
rect -1857 2007 -1841 2041
rect -1773 2007 -1757 2041
rect -1579 2007 -1563 2041
rect -1495 2007 -1479 2041
rect -1301 2007 -1285 2041
rect -1217 2007 -1201 2041
rect -1023 2007 -1007 2041
rect -939 2007 -923 2041
rect -745 2007 -729 2041
rect -661 2007 -645 2041
rect -467 2007 -451 2041
rect -383 2007 -367 2041
rect -189 2007 -173 2041
rect -105 2007 -89 2041
rect 89 2007 105 2041
rect 173 2007 189 2041
rect 367 2007 383 2041
rect 451 2007 467 2041
rect 645 2007 661 2041
rect 729 2007 745 2041
rect 923 2007 939 2041
rect 1007 2007 1023 2041
rect 1201 2007 1217 2041
rect 1285 2007 1301 2041
rect 1479 2007 1495 2041
rect 1563 2007 1579 2041
rect 1757 2007 1773 2041
rect 1841 2007 1857 2041
rect 2035 2007 2051 2041
rect 2119 2007 2135 2041
rect 2313 2007 2329 2041
rect 2397 2007 2413 2041
rect 2591 2007 2607 2041
rect 2675 2007 2691 2041
rect 2869 2007 2885 2041
rect 2953 2007 2969 2041
rect 3147 2007 3163 2041
rect 3231 2007 3247 2041
rect 3425 2007 3441 2041
rect 3509 2007 3525 2041
rect 3703 2007 3719 2041
rect 3787 2007 3803 2041
rect 3981 2007 3997 2041
rect 4065 2007 4081 2041
rect 4259 2007 4275 2041
rect 4343 2007 4359 2041
rect 4537 2007 4553 2041
rect 4621 2007 4637 2041
rect 4815 2007 4831 2041
rect 4899 2007 4915 2041
rect 5093 2007 5109 2041
rect 5177 2007 5193 2041
rect 5371 2007 5387 2041
rect 5455 2007 5471 2041
rect 5649 2007 5665 2041
rect 5733 2007 5749 2041
rect 5927 2007 5943 2041
rect 6011 2007 6027 2041
rect 6205 2007 6221 2041
rect 6289 2007 6305 2041
rect 6483 2007 6499 2041
rect 6567 2007 6583 2041
rect 6761 2007 6777 2041
rect 6845 2007 6861 2041
rect 7039 2007 7055 2041
rect 7123 2007 7139 2041
rect 7317 2007 7333 2041
rect 7401 2007 7417 2041
rect 7595 2007 7611 2041
rect 7679 2007 7695 2041
rect 7873 2007 7889 2041
rect 7957 2007 7973 2041
rect 8151 2007 8167 2041
rect 8235 2007 8251 2041
rect 8429 2007 8445 2041
rect 8513 2007 8529 2041
rect 8707 2007 8723 2041
rect 8791 2007 8807 2041
rect 8985 2007 9001 2041
rect 9069 2007 9085 2041
rect 9263 2007 9279 2041
rect 9347 2007 9363 2041
rect 9541 2007 9557 2041
rect 9625 2007 9641 2041
rect 9819 2007 9835 2041
rect 9903 2007 9919 2041
rect 10097 2007 10113 2041
rect 10181 2007 10197 2041
rect 10375 2007 10391 2041
rect 10459 2007 10475 2041
rect 10653 2007 10669 2041
rect 10737 2007 10753 2041
rect 10931 2007 10947 2041
rect 11015 2007 11031 2041
rect 11209 2007 11225 2041
rect 11293 2007 11309 2041
rect 11487 2007 11503 2041
rect 11571 2007 11587 2041
rect 11765 2007 11781 2041
rect 11849 2007 11865 2041
rect 12043 2007 12059 2041
rect 12127 2007 12143 2041
rect 12321 2007 12337 2041
rect 12405 2007 12421 2041
rect 12599 2007 12615 2041
rect 12683 2007 12699 2041
rect 12877 2007 12893 2041
rect 12961 2007 12977 2041
rect 13155 2007 13171 2041
rect 13239 2007 13255 2041
rect 13433 2007 13449 2041
rect 13517 2007 13533 2041
rect 13711 2007 13727 2041
rect 13795 2007 13811 2041
rect 13989 2007 14005 2041
rect 14073 2007 14089 2041
rect 14267 2007 14283 2041
rect 14351 2007 14367 2041
rect 14545 2007 14561 2041
rect 14629 2007 14645 2041
rect 14823 2007 14839 2041
rect 14907 2007 14923 2041
rect 15101 2007 15117 2041
rect 15185 2007 15201 2041
rect 15379 2007 15395 2041
rect 15463 2007 15479 2041
rect 15657 2007 15673 2041
rect 15741 2007 15757 2041
rect 15935 2007 15951 2041
rect 16019 2007 16035 2041
rect 16213 2007 16229 2041
rect 16297 2007 16313 2041
rect 16491 2007 16507 2041
rect 16575 2007 16591 2041
rect 16769 2007 16785 2041
rect 16853 2007 16869 2041
rect 17047 2007 17063 2041
rect 17131 2007 17147 2041
rect 17325 2007 17341 2041
rect 17409 2007 17425 2041
rect 17603 2007 17619 2041
rect 17687 2007 17703 2041
rect -17749 1957 -17715 1973
rect -17749 -2035 -17715 -2019
rect -17591 1957 -17557 1973
rect -17591 -2035 -17557 -2019
rect -17471 1957 -17437 1973
rect -17471 -2035 -17437 -2019
rect -17313 1957 -17279 1973
rect -17313 -2035 -17279 -2019
rect -17193 1957 -17159 1973
rect -17193 -2035 -17159 -2019
rect -17035 1957 -17001 1973
rect -17035 -2035 -17001 -2019
rect -16915 1957 -16881 1973
rect -16915 -2035 -16881 -2019
rect -16757 1957 -16723 1973
rect -16757 -2035 -16723 -2019
rect -16637 1957 -16603 1973
rect -16637 -2035 -16603 -2019
rect -16479 1957 -16445 1973
rect -16479 -2035 -16445 -2019
rect -16359 1957 -16325 1973
rect -16359 -2035 -16325 -2019
rect -16201 1957 -16167 1973
rect -16201 -2035 -16167 -2019
rect -16081 1957 -16047 1973
rect -16081 -2035 -16047 -2019
rect -15923 1957 -15889 1973
rect -15923 -2035 -15889 -2019
rect -15803 1957 -15769 1973
rect -15803 -2035 -15769 -2019
rect -15645 1957 -15611 1973
rect -15645 -2035 -15611 -2019
rect -15525 1957 -15491 1973
rect -15525 -2035 -15491 -2019
rect -15367 1957 -15333 1973
rect -15367 -2035 -15333 -2019
rect -15247 1957 -15213 1973
rect -15247 -2035 -15213 -2019
rect -15089 1957 -15055 1973
rect -15089 -2035 -15055 -2019
rect -14969 1957 -14935 1973
rect -14969 -2035 -14935 -2019
rect -14811 1957 -14777 1973
rect -14811 -2035 -14777 -2019
rect -14691 1957 -14657 1973
rect -14691 -2035 -14657 -2019
rect -14533 1957 -14499 1973
rect -14533 -2035 -14499 -2019
rect -14413 1957 -14379 1973
rect -14413 -2035 -14379 -2019
rect -14255 1957 -14221 1973
rect -14255 -2035 -14221 -2019
rect -14135 1957 -14101 1973
rect -14135 -2035 -14101 -2019
rect -13977 1957 -13943 1973
rect -13977 -2035 -13943 -2019
rect -13857 1957 -13823 1973
rect -13857 -2035 -13823 -2019
rect -13699 1957 -13665 1973
rect -13699 -2035 -13665 -2019
rect -13579 1957 -13545 1973
rect -13579 -2035 -13545 -2019
rect -13421 1957 -13387 1973
rect -13421 -2035 -13387 -2019
rect -13301 1957 -13267 1973
rect -13301 -2035 -13267 -2019
rect -13143 1957 -13109 1973
rect -13143 -2035 -13109 -2019
rect -13023 1957 -12989 1973
rect -13023 -2035 -12989 -2019
rect -12865 1957 -12831 1973
rect -12865 -2035 -12831 -2019
rect -12745 1957 -12711 1973
rect -12745 -2035 -12711 -2019
rect -12587 1957 -12553 1973
rect -12587 -2035 -12553 -2019
rect -12467 1957 -12433 1973
rect -12467 -2035 -12433 -2019
rect -12309 1957 -12275 1973
rect -12309 -2035 -12275 -2019
rect -12189 1957 -12155 1973
rect -12189 -2035 -12155 -2019
rect -12031 1957 -11997 1973
rect -12031 -2035 -11997 -2019
rect -11911 1957 -11877 1973
rect -11911 -2035 -11877 -2019
rect -11753 1957 -11719 1973
rect -11753 -2035 -11719 -2019
rect -11633 1957 -11599 1973
rect -11633 -2035 -11599 -2019
rect -11475 1957 -11441 1973
rect -11475 -2035 -11441 -2019
rect -11355 1957 -11321 1973
rect -11355 -2035 -11321 -2019
rect -11197 1957 -11163 1973
rect -11197 -2035 -11163 -2019
rect -11077 1957 -11043 1973
rect -11077 -2035 -11043 -2019
rect -10919 1957 -10885 1973
rect -10919 -2035 -10885 -2019
rect -10799 1957 -10765 1973
rect -10799 -2035 -10765 -2019
rect -10641 1957 -10607 1973
rect -10641 -2035 -10607 -2019
rect -10521 1957 -10487 1973
rect -10521 -2035 -10487 -2019
rect -10363 1957 -10329 1973
rect -10363 -2035 -10329 -2019
rect -10243 1957 -10209 1973
rect -10243 -2035 -10209 -2019
rect -10085 1957 -10051 1973
rect -10085 -2035 -10051 -2019
rect -9965 1957 -9931 1973
rect -9965 -2035 -9931 -2019
rect -9807 1957 -9773 1973
rect -9807 -2035 -9773 -2019
rect -9687 1957 -9653 1973
rect -9687 -2035 -9653 -2019
rect -9529 1957 -9495 1973
rect -9529 -2035 -9495 -2019
rect -9409 1957 -9375 1973
rect -9409 -2035 -9375 -2019
rect -9251 1957 -9217 1973
rect -9251 -2035 -9217 -2019
rect -9131 1957 -9097 1973
rect -9131 -2035 -9097 -2019
rect -8973 1957 -8939 1973
rect -8973 -2035 -8939 -2019
rect -8853 1957 -8819 1973
rect -8853 -2035 -8819 -2019
rect -8695 1957 -8661 1973
rect -8695 -2035 -8661 -2019
rect -8575 1957 -8541 1973
rect -8575 -2035 -8541 -2019
rect -8417 1957 -8383 1973
rect -8417 -2035 -8383 -2019
rect -8297 1957 -8263 1973
rect -8297 -2035 -8263 -2019
rect -8139 1957 -8105 1973
rect -8139 -2035 -8105 -2019
rect -8019 1957 -7985 1973
rect -8019 -2035 -7985 -2019
rect -7861 1957 -7827 1973
rect -7861 -2035 -7827 -2019
rect -7741 1957 -7707 1973
rect -7741 -2035 -7707 -2019
rect -7583 1957 -7549 1973
rect -7583 -2035 -7549 -2019
rect -7463 1957 -7429 1973
rect -7463 -2035 -7429 -2019
rect -7305 1957 -7271 1973
rect -7305 -2035 -7271 -2019
rect -7185 1957 -7151 1973
rect -7185 -2035 -7151 -2019
rect -7027 1957 -6993 1973
rect -7027 -2035 -6993 -2019
rect -6907 1957 -6873 1973
rect -6907 -2035 -6873 -2019
rect -6749 1957 -6715 1973
rect -6749 -2035 -6715 -2019
rect -6629 1957 -6595 1973
rect -6629 -2035 -6595 -2019
rect -6471 1957 -6437 1973
rect -6471 -2035 -6437 -2019
rect -6351 1957 -6317 1973
rect -6351 -2035 -6317 -2019
rect -6193 1957 -6159 1973
rect -6193 -2035 -6159 -2019
rect -6073 1957 -6039 1973
rect -6073 -2035 -6039 -2019
rect -5915 1957 -5881 1973
rect -5915 -2035 -5881 -2019
rect -5795 1957 -5761 1973
rect -5795 -2035 -5761 -2019
rect -5637 1957 -5603 1973
rect -5637 -2035 -5603 -2019
rect -5517 1957 -5483 1973
rect -5517 -2035 -5483 -2019
rect -5359 1957 -5325 1973
rect -5359 -2035 -5325 -2019
rect -5239 1957 -5205 1973
rect -5239 -2035 -5205 -2019
rect -5081 1957 -5047 1973
rect -5081 -2035 -5047 -2019
rect -4961 1957 -4927 1973
rect -4961 -2035 -4927 -2019
rect -4803 1957 -4769 1973
rect -4803 -2035 -4769 -2019
rect -4683 1957 -4649 1973
rect -4683 -2035 -4649 -2019
rect -4525 1957 -4491 1973
rect -4525 -2035 -4491 -2019
rect -4405 1957 -4371 1973
rect -4405 -2035 -4371 -2019
rect -4247 1957 -4213 1973
rect -4247 -2035 -4213 -2019
rect -4127 1957 -4093 1973
rect -4127 -2035 -4093 -2019
rect -3969 1957 -3935 1973
rect -3969 -2035 -3935 -2019
rect -3849 1957 -3815 1973
rect -3849 -2035 -3815 -2019
rect -3691 1957 -3657 1973
rect -3691 -2035 -3657 -2019
rect -3571 1957 -3537 1973
rect -3571 -2035 -3537 -2019
rect -3413 1957 -3379 1973
rect -3413 -2035 -3379 -2019
rect -3293 1957 -3259 1973
rect -3293 -2035 -3259 -2019
rect -3135 1957 -3101 1973
rect -3135 -2035 -3101 -2019
rect -3015 1957 -2981 1973
rect -3015 -2035 -2981 -2019
rect -2857 1957 -2823 1973
rect -2857 -2035 -2823 -2019
rect -2737 1957 -2703 1973
rect -2737 -2035 -2703 -2019
rect -2579 1957 -2545 1973
rect -2579 -2035 -2545 -2019
rect -2459 1957 -2425 1973
rect -2459 -2035 -2425 -2019
rect -2301 1957 -2267 1973
rect -2301 -2035 -2267 -2019
rect -2181 1957 -2147 1973
rect -2181 -2035 -2147 -2019
rect -2023 1957 -1989 1973
rect -2023 -2035 -1989 -2019
rect -1903 1957 -1869 1973
rect -1903 -2035 -1869 -2019
rect -1745 1957 -1711 1973
rect -1745 -2035 -1711 -2019
rect -1625 1957 -1591 1973
rect -1625 -2035 -1591 -2019
rect -1467 1957 -1433 1973
rect -1467 -2035 -1433 -2019
rect -1347 1957 -1313 1973
rect -1347 -2035 -1313 -2019
rect -1189 1957 -1155 1973
rect -1189 -2035 -1155 -2019
rect -1069 1957 -1035 1973
rect -1069 -2035 -1035 -2019
rect -911 1957 -877 1973
rect -911 -2035 -877 -2019
rect -791 1957 -757 1973
rect -791 -2035 -757 -2019
rect -633 1957 -599 1973
rect -633 -2035 -599 -2019
rect -513 1957 -479 1973
rect -513 -2035 -479 -2019
rect -355 1957 -321 1973
rect -355 -2035 -321 -2019
rect -235 1957 -201 1973
rect -235 -2035 -201 -2019
rect -77 1957 -43 1973
rect -77 -2035 -43 -2019
rect 43 1957 77 1973
rect 43 -2035 77 -2019
rect 201 1957 235 1973
rect 201 -2035 235 -2019
rect 321 1957 355 1973
rect 321 -2035 355 -2019
rect 479 1957 513 1973
rect 479 -2035 513 -2019
rect 599 1957 633 1973
rect 599 -2035 633 -2019
rect 757 1957 791 1973
rect 757 -2035 791 -2019
rect 877 1957 911 1973
rect 877 -2035 911 -2019
rect 1035 1957 1069 1973
rect 1035 -2035 1069 -2019
rect 1155 1957 1189 1973
rect 1155 -2035 1189 -2019
rect 1313 1957 1347 1973
rect 1313 -2035 1347 -2019
rect 1433 1957 1467 1973
rect 1433 -2035 1467 -2019
rect 1591 1957 1625 1973
rect 1591 -2035 1625 -2019
rect 1711 1957 1745 1973
rect 1711 -2035 1745 -2019
rect 1869 1957 1903 1973
rect 1869 -2035 1903 -2019
rect 1989 1957 2023 1973
rect 1989 -2035 2023 -2019
rect 2147 1957 2181 1973
rect 2147 -2035 2181 -2019
rect 2267 1957 2301 1973
rect 2267 -2035 2301 -2019
rect 2425 1957 2459 1973
rect 2425 -2035 2459 -2019
rect 2545 1957 2579 1973
rect 2545 -2035 2579 -2019
rect 2703 1957 2737 1973
rect 2703 -2035 2737 -2019
rect 2823 1957 2857 1973
rect 2823 -2035 2857 -2019
rect 2981 1957 3015 1973
rect 2981 -2035 3015 -2019
rect 3101 1957 3135 1973
rect 3101 -2035 3135 -2019
rect 3259 1957 3293 1973
rect 3259 -2035 3293 -2019
rect 3379 1957 3413 1973
rect 3379 -2035 3413 -2019
rect 3537 1957 3571 1973
rect 3537 -2035 3571 -2019
rect 3657 1957 3691 1973
rect 3657 -2035 3691 -2019
rect 3815 1957 3849 1973
rect 3815 -2035 3849 -2019
rect 3935 1957 3969 1973
rect 3935 -2035 3969 -2019
rect 4093 1957 4127 1973
rect 4093 -2035 4127 -2019
rect 4213 1957 4247 1973
rect 4213 -2035 4247 -2019
rect 4371 1957 4405 1973
rect 4371 -2035 4405 -2019
rect 4491 1957 4525 1973
rect 4491 -2035 4525 -2019
rect 4649 1957 4683 1973
rect 4649 -2035 4683 -2019
rect 4769 1957 4803 1973
rect 4769 -2035 4803 -2019
rect 4927 1957 4961 1973
rect 4927 -2035 4961 -2019
rect 5047 1957 5081 1973
rect 5047 -2035 5081 -2019
rect 5205 1957 5239 1973
rect 5205 -2035 5239 -2019
rect 5325 1957 5359 1973
rect 5325 -2035 5359 -2019
rect 5483 1957 5517 1973
rect 5483 -2035 5517 -2019
rect 5603 1957 5637 1973
rect 5603 -2035 5637 -2019
rect 5761 1957 5795 1973
rect 5761 -2035 5795 -2019
rect 5881 1957 5915 1973
rect 5881 -2035 5915 -2019
rect 6039 1957 6073 1973
rect 6039 -2035 6073 -2019
rect 6159 1957 6193 1973
rect 6159 -2035 6193 -2019
rect 6317 1957 6351 1973
rect 6317 -2035 6351 -2019
rect 6437 1957 6471 1973
rect 6437 -2035 6471 -2019
rect 6595 1957 6629 1973
rect 6595 -2035 6629 -2019
rect 6715 1957 6749 1973
rect 6715 -2035 6749 -2019
rect 6873 1957 6907 1973
rect 6873 -2035 6907 -2019
rect 6993 1957 7027 1973
rect 6993 -2035 7027 -2019
rect 7151 1957 7185 1973
rect 7151 -2035 7185 -2019
rect 7271 1957 7305 1973
rect 7271 -2035 7305 -2019
rect 7429 1957 7463 1973
rect 7429 -2035 7463 -2019
rect 7549 1957 7583 1973
rect 7549 -2035 7583 -2019
rect 7707 1957 7741 1973
rect 7707 -2035 7741 -2019
rect 7827 1957 7861 1973
rect 7827 -2035 7861 -2019
rect 7985 1957 8019 1973
rect 7985 -2035 8019 -2019
rect 8105 1957 8139 1973
rect 8105 -2035 8139 -2019
rect 8263 1957 8297 1973
rect 8263 -2035 8297 -2019
rect 8383 1957 8417 1973
rect 8383 -2035 8417 -2019
rect 8541 1957 8575 1973
rect 8541 -2035 8575 -2019
rect 8661 1957 8695 1973
rect 8661 -2035 8695 -2019
rect 8819 1957 8853 1973
rect 8819 -2035 8853 -2019
rect 8939 1957 8973 1973
rect 8939 -2035 8973 -2019
rect 9097 1957 9131 1973
rect 9097 -2035 9131 -2019
rect 9217 1957 9251 1973
rect 9217 -2035 9251 -2019
rect 9375 1957 9409 1973
rect 9375 -2035 9409 -2019
rect 9495 1957 9529 1973
rect 9495 -2035 9529 -2019
rect 9653 1957 9687 1973
rect 9653 -2035 9687 -2019
rect 9773 1957 9807 1973
rect 9773 -2035 9807 -2019
rect 9931 1957 9965 1973
rect 9931 -2035 9965 -2019
rect 10051 1957 10085 1973
rect 10051 -2035 10085 -2019
rect 10209 1957 10243 1973
rect 10209 -2035 10243 -2019
rect 10329 1957 10363 1973
rect 10329 -2035 10363 -2019
rect 10487 1957 10521 1973
rect 10487 -2035 10521 -2019
rect 10607 1957 10641 1973
rect 10607 -2035 10641 -2019
rect 10765 1957 10799 1973
rect 10765 -2035 10799 -2019
rect 10885 1957 10919 1973
rect 10885 -2035 10919 -2019
rect 11043 1957 11077 1973
rect 11043 -2035 11077 -2019
rect 11163 1957 11197 1973
rect 11163 -2035 11197 -2019
rect 11321 1957 11355 1973
rect 11321 -2035 11355 -2019
rect 11441 1957 11475 1973
rect 11441 -2035 11475 -2019
rect 11599 1957 11633 1973
rect 11599 -2035 11633 -2019
rect 11719 1957 11753 1973
rect 11719 -2035 11753 -2019
rect 11877 1957 11911 1973
rect 11877 -2035 11911 -2019
rect 11997 1957 12031 1973
rect 11997 -2035 12031 -2019
rect 12155 1957 12189 1973
rect 12155 -2035 12189 -2019
rect 12275 1957 12309 1973
rect 12275 -2035 12309 -2019
rect 12433 1957 12467 1973
rect 12433 -2035 12467 -2019
rect 12553 1957 12587 1973
rect 12553 -2035 12587 -2019
rect 12711 1957 12745 1973
rect 12711 -2035 12745 -2019
rect 12831 1957 12865 1973
rect 12831 -2035 12865 -2019
rect 12989 1957 13023 1973
rect 12989 -2035 13023 -2019
rect 13109 1957 13143 1973
rect 13109 -2035 13143 -2019
rect 13267 1957 13301 1973
rect 13267 -2035 13301 -2019
rect 13387 1957 13421 1973
rect 13387 -2035 13421 -2019
rect 13545 1957 13579 1973
rect 13545 -2035 13579 -2019
rect 13665 1957 13699 1973
rect 13665 -2035 13699 -2019
rect 13823 1957 13857 1973
rect 13823 -2035 13857 -2019
rect 13943 1957 13977 1973
rect 13943 -2035 13977 -2019
rect 14101 1957 14135 1973
rect 14101 -2035 14135 -2019
rect 14221 1957 14255 1973
rect 14221 -2035 14255 -2019
rect 14379 1957 14413 1973
rect 14379 -2035 14413 -2019
rect 14499 1957 14533 1973
rect 14499 -2035 14533 -2019
rect 14657 1957 14691 1973
rect 14657 -2035 14691 -2019
rect 14777 1957 14811 1973
rect 14777 -2035 14811 -2019
rect 14935 1957 14969 1973
rect 14935 -2035 14969 -2019
rect 15055 1957 15089 1973
rect 15055 -2035 15089 -2019
rect 15213 1957 15247 1973
rect 15213 -2035 15247 -2019
rect 15333 1957 15367 1973
rect 15333 -2035 15367 -2019
rect 15491 1957 15525 1973
rect 15491 -2035 15525 -2019
rect 15611 1957 15645 1973
rect 15611 -2035 15645 -2019
rect 15769 1957 15803 1973
rect 15769 -2035 15803 -2019
rect 15889 1957 15923 1973
rect 15889 -2035 15923 -2019
rect 16047 1957 16081 1973
rect 16047 -2035 16081 -2019
rect 16167 1957 16201 1973
rect 16167 -2035 16201 -2019
rect 16325 1957 16359 1973
rect 16325 -2035 16359 -2019
rect 16445 1957 16479 1973
rect 16445 -2035 16479 -2019
rect 16603 1957 16637 1973
rect 16603 -2035 16637 -2019
rect 16723 1957 16757 1973
rect 16723 -2035 16757 -2019
rect 16881 1957 16915 1973
rect 16881 -2035 16915 -2019
rect 17001 1957 17035 1973
rect 17001 -2035 17035 -2019
rect 17159 1957 17193 1973
rect 17159 -2035 17193 -2019
rect 17279 1957 17313 1973
rect 17279 -2035 17313 -2019
rect 17437 1957 17471 1973
rect 17437 -2035 17471 -2019
rect 17557 1957 17591 1973
rect 17557 -2035 17591 -2019
rect 17715 1957 17749 1973
rect 17715 -2035 17749 -2019
<< viali >>
rect -17687 2007 -17619 2041
rect -17409 2007 -17341 2041
rect -17131 2007 -17063 2041
rect -16853 2007 -16785 2041
rect -16575 2007 -16507 2041
rect -16297 2007 -16229 2041
rect -16019 2007 -15951 2041
rect -15741 2007 -15673 2041
rect -15463 2007 -15395 2041
rect -15185 2007 -15117 2041
rect -14907 2007 -14839 2041
rect -14629 2007 -14561 2041
rect -14351 2007 -14283 2041
rect -14073 2007 -14005 2041
rect -13795 2007 -13727 2041
rect -13517 2007 -13449 2041
rect -13239 2007 -13171 2041
rect -12961 2007 -12893 2041
rect -12683 2007 -12615 2041
rect -12405 2007 -12337 2041
rect -12127 2007 -12059 2041
rect -11849 2007 -11781 2041
rect -11571 2007 -11503 2041
rect -11293 2007 -11225 2041
rect -11015 2007 -10947 2041
rect -10737 2007 -10669 2041
rect -10459 2007 -10391 2041
rect -10181 2007 -10113 2041
rect -9903 2007 -9835 2041
rect -9625 2007 -9557 2041
rect -9347 2007 -9279 2041
rect -9069 2007 -9001 2041
rect -8791 2007 -8723 2041
rect -8513 2007 -8445 2041
rect -8235 2007 -8167 2041
rect -7957 2007 -7889 2041
rect -7679 2007 -7611 2041
rect -7401 2007 -7333 2041
rect -7123 2007 -7055 2041
rect -6845 2007 -6777 2041
rect -6567 2007 -6499 2041
rect -6289 2007 -6221 2041
rect -6011 2007 -5943 2041
rect -5733 2007 -5665 2041
rect -5455 2007 -5387 2041
rect -5177 2007 -5109 2041
rect -4899 2007 -4831 2041
rect -4621 2007 -4553 2041
rect -4343 2007 -4275 2041
rect -4065 2007 -3997 2041
rect -3787 2007 -3719 2041
rect -3509 2007 -3441 2041
rect -3231 2007 -3163 2041
rect -2953 2007 -2885 2041
rect -2675 2007 -2607 2041
rect -2397 2007 -2329 2041
rect -2119 2007 -2051 2041
rect -1841 2007 -1773 2041
rect -1563 2007 -1495 2041
rect -1285 2007 -1217 2041
rect -1007 2007 -939 2041
rect -729 2007 -661 2041
rect -451 2007 -383 2041
rect -173 2007 -105 2041
rect 105 2007 173 2041
rect 383 2007 451 2041
rect 661 2007 729 2041
rect 939 2007 1007 2041
rect 1217 2007 1285 2041
rect 1495 2007 1563 2041
rect 1773 2007 1841 2041
rect 2051 2007 2119 2041
rect 2329 2007 2397 2041
rect 2607 2007 2675 2041
rect 2885 2007 2953 2041
rect 3163 2007 3231 2041
rect 3441 2007 3509 2041
rect 3719 2007 3787 2041
rect 3997 2007 4065 2041
rect 4275 2007 4343 2041
rect 4553 2007 4621 2041
rect 4831 2007 4899 2041
rect 5109 2007 5177 2041
rect 5387 2007 5455 2041
rect 5665 2007 5733 2041
rect 5943 2007 6011 2041
rect 6221 2007 6289 2041
rect 6499 2007 6567 2041
rect 6777 2007 6845 2041
rect 7055 2007 7123 2041
rect 7333 2007 7401 2041
rect 7611 2007 7679 2041
rect 7889 2007 7957 2041
rect 8167 2007 8235 2041
rect 8445 2007 8513 2041
rect 8723 2007 8791 2041
rect 9001 2007 9069 2041
rect 9279 2007 9347 2041
rect 9557 2007 9625 2041
rect 9835 2007 9903 2041
rect 10113 2007 10181 2041
rect 10391 2007 10459 2041
rect 10669 2007 10737 2041
rect 10947 2007 11015 2041
rect 11225 2007 11293 2041
rect 11503 2007 11571 2041
rect 11781 2007 11849 2041
rect 12059 2007 12127 2041
rect 12337 2007 12405 2041
rect 12615 2007 12683 2041
rect 12893 2007 12961 2041
rect 13171 2007 13239 2041
rect 13449 2007 13517 2041
rect 13727 2007 13795 2041
rect 14005 2007 14073 2041
rect 14283 2007 14351 2041
rect 14561 2007 14629 2041
rect 14839 2007 14907 2041
rect 15117 2007 15185 2041
rect 15395 2007 15463 2041
rect 15673 2007 15741 2041
rect 15951 2007 16019 2041
rect 16229 2007 16297 2041
rect 16507 2007 16575 2041
rect 16785 2007 16853 2041
rect 17063 2007 17131 2041
rect 17341 2007 17409 2041
rect 17619 2007 17687 2041
rect -17749 -2019 -17715 1957
rect -17591 -2019 -17557 1957
rect -17471 -2019 -17437 1957
rect -17313 -2019 -17279 1957
rect -17193 -2019 -17159 1957
rect -17035 -2019 -17001 1957
rect -16915 -2019 -16881 1957
rect -16757 -2019 -16723 1957
rect -16637 -2019 -16603 1957
rect -16479 -2019 -16445 1957
rect -16359 -2019 -16325 1957
rect -16201 -2019 -16167 1957
rect -16081 -2019 -16047 1957
rect -15923 -2019 -15889 1957
rect -15803 -2019 -15769 1957
rect -15645 -2019 -15611 1957
rect -15525 -2019 -15491 1957
rect -15367 -2019 -15333 1957
rect -15247 -2019 -15213 1957
rect -15089 -2019 -15055 1957
rect -14969 -2019 -14935 1957
rect -14811 -2019 -14777 1957
rect -14691 -2019 -14657 1957
rect -14533 -2019 -14499 1957
rect -14413 -2019 -14379 1957
rect -14255 -2019 -14221 1957
rect -14135 -2019 -14101 1957
rect -13977 -2019 -13943 1957
rect -13857 -2019 -13823 1957
rect -13699 -2019 -13665 1957
rect -13579 -2019 -13545 1957
rect -13421 -2019 -13387 1957
rect -13301 -2019 -13267 1957
rect -13143 -2019 -13109 1957
rect -13023 -2019 -12989 1957
rect -12865 -2019 -12831 1957
rect -12745 -2019 -12711 1957
rect -12587 -2019 -12553 1957
rect -12467 -2019 -12433 1957
rect -12309 -2019 -12275 1957
rect -12189 -2019 -12155 1957
rect -12031 -2019 -11997 1957
rect -11911 -2019 -11877 1957
rect -11753 -2019 -11719 1957
rect -11633 -2019 -11599 1957
rect -11475 -2019 -11441 1957
rect -11355 -2019 -11321 1957
rect -11197 -2019 -11163 1957
rect -11077 -2019 -11043 1957
rect -10919 -2019 -10885 1957
rect -10799 -2019 -10765 1957
rect -10641 -2019 -10607 1957
rect -10521 -2019 -10487 1957
rect -10363 -2019 -10329 1957
rect -10243 -2019 -10209 1957
rect -10085 -2019 -10051 1957
rect -9965 -2019 -9931 1957
rect -9807 -2019 -9773 1957
rect -9687 -2019 -9653 1957
rect -9529 -2019 -9495 1957
rect -9409 -2019 -9375 1957
rect -9251 -2019 -9217 1957
rect -9131 -2019 -9097 1957
rect -8973 -2019 -8939 1957
rect -8853 -2019 -8819 1957
rect -8695 -2019 -8661 1957
rect -8575 -2019 -8541 1957
rect -8417 -2019 -8383 1957
rect -8297 -2019 -8263 1957
rect -8139 -2019 -8105 1957
rect -8019 -2019 -7985 1957
rect -7861 -2019 -7827 1957
rect -7741 -2019 -7707 1957
rect -7583 -2019 -7549 1957
rect -7463 -2019 -7429 1957
rect -7305 -2019 -7271 1957
rect -7185 -2019 -7151 1957
rect -7027 -2019 -6993 1957
rect -6907 -2019 -6873 1957
rect -6749 -2019 -6715 1957
rect -6629 -2019 -6595 1957
rect -6471 -2019 -6437 1957
rect -6351 -2019 -6317 1957
rect -6193 -2019 -6159 1957
rect -6073 -2019 -6039 1957
rect -5915 -2019 -5881 1957
rect -5795 -2019 -5761 1957
rect -5637 -2019 -5603 1957
rect -5517 -2019 -5483 1957
rect -5359 -2019 -5325 1957
rect -5239 -2019 -5205 1957
rect -5081 -2019 -5047 1957
rect -4961 -2019 -4927 1957
rect -4803 -2019 -4769 1957
rect -4683 -2019 -4649 1957
rect -4525 -2019 -4491 1957
rect -4405 -2019 -4371 1957
rect -4247 -2019 -4213 1957
rect -4127 -2019 -4093 1957
rect -3969 -2019 -3935 1957
rect -3849 -2019 -3815 1957
rect -3691 -2019 -3657 1957
rect -3571 -2019 -3537 1957
rect -3413 -2019 -3379 1957
rect -3293 -2019 -3259 1957
rect -3135 -2019 -3101 1957
rect -3015 -2019 -2981 1957
rect -2857 -2019 -2823 1957
rect -2737 -2019 -2703 1957
rect -2579 -2019 -2545 1957
rect -2459 -2019 -2425 1957
rect -2301 -2019 -2267 1957
rect -2181 -2019 -2147 1957
rect -2023 -2019 -1989 1957
rect -1903 -2019 -1869 1957
rect -1745 -2019 -1711 1957
rect -1625 -2019 -1591 1957
rect -1467 -2019 -1433 1957
rect -1347 -2019 -1313 1957
rect -1189 -2019 -1155 1957
rect -1069 -2019 -1035 1957
rect -911 -2019 -877 1957
rect -791 -2019 -757 1957
rect -633 -2019 -599 1957
rect -513 -2019 -479 1957
rect -355 -2019 -321 1957
rect -235 -2019 -201 1957
rect -77 -2019 -43 1957
rect 43 -2019 77 1957
rect 201 -2019 235 1957
rect 321 -2019 355 1957
rect 479 -2019 513 1957
rect 599 -2019 633 1957
rect 757 -2019 791 1957
rect 877 -2019 911 1957
rect 1035 -2019 1069 1957
rect 1155 -2019 1189 1957
rect 1313 -2019 1347 1957
rect 1433 -2019 1467 1957
rect 1591 -2019 1625 1957
rect 1711 -2019 1745 1957
rect 1869 -2019 1903 1957
rect 1989 -2019 2023 1957
rect 2147 -2019 2181 1957
rect 2267 -2019 2301 1957
rect 2425 -2019 2459 1957
rect 2545 -2019 2579 1957
rect 2703 -2019 2737 1957
rect 2823 -2019 2857 1957
rect 2981 -2019 3015 1957
rect 3101 -2019 3135 1957
rect 3259 -2019 3293 1957
rect 3379 -2019 3413 1957
rect 3537 -2019 3571 1957
rect 3657 -2019 3691 1957
rect 3815 -2019 3849 1957
rect 3935 -2019 3969 1957
rect 4093 -2019 4127 1957
rect 4213 -2019 4247 1957
rect 4371 -2019 4405 1957
rect 4491 -2019 4525 1957
rect 4649 -2019 4683 1957
rect 4769 -2019 4803 1957
rect 4927 -2019 4961 1957
rect 5047 -2019 5081 1957
rect 5205 -2019 5239 1957
rect 5325 -2019 5359 1957
rect 5483 -2019 5517 1957
rect 5603 -2019 5637 1957
rect 5761 -2019 5795 1957
rect 5881 -2019 5915 1957
rect 6039 -2019 6073 1957
rect 6159 -2019 6193 1957
rect 6317 -2019 6351 1957
rect 6437 -2019 6471 1957
rect 6595 -2019 6629 1957
rect 6715 -2019 6749 1957
rect 6873 -2019 6907 1957
rect 6993 -2019 7027 1957
rect 7151 -2019 7185 1957
rect 7271 -2019 7305 1957
rect 7429 -2019 7463 1957
rect 7549 -2019 7583 1957
rect 7707 -2019 7741 1957
rect 7827 -2019 7861 1957
rect 7985 -2019 8019 1957
rect 8105 -2019 8139 1957
rect 8263 -2019 8297 1957
rect 8383 -2019 8417 1957
rect 8541 -2019 8575 1957
rect 8661 -2019 8695 1957
rect 8819 -2019 8853 1957
rect 8939 -2019 8973 1957
rect 9097 -2019 9131 1957
rect 9217 -2019 9251 1957
rect 9375 -2019 9409 1957
rect 9495 -2019 9529 1957
rect 9653 -2019 9687 1957
rect 9773 -2019 9807 1957
rect 9931 -2019 9965 1957
rect 10051 -2019 10085 1957
rect 10209 -2019 10243 1957
rect 10329 -2019 10363 1957
rect 10487 -2019 10521 1957
rect 10607 -2019 10641 1957
rect 10765 -2019 10799 1957
rect 10885 -2019 10919 1957
rect 11043 -2019 11077 1957
rect 11163 -2019 11197 1957
rect 11321 -2019 11355 1957
rect 11441 -2019 11475 1957
rect 11599 -2019 11633 1957
rect 11719 -2019 11753 1957
rect 11877 -2019 11911 1957
rect 11997 -2019 12031 1957
rect 12155 -2019 12189 1957
rect 12275 -2019 12309 1957
rect 12433 -2019 12467 1957
rect 12553 -2019 12587 1957
rect 12711 -2019 12745 1957
rect 12831 -2019 12865 1957
rect 12989 -2019 13023 1957
rect 13109 -2019 13143 1957
rect 13267 -2019 13301 1957
rect 13387 -2019 13421 1957
rect 13545 -2019 13579 1957
rect 13665 -2019 13699 1957
rect 13823 -2019 13857 1957
rect 13943 -2019 13977 1957
rect 14101 -2019 14135 1957
rect 14221 -2019 14255 1957
rect 14379 -2019 14413 1957
rect 14499 -2019 14533 1957
rect 14657 -2019 14691 1957
rect 14777 -2019 14811 1957
rect 14935 -2019 14969 1957
rect 15055 -2019 15089 1957
rect 15213 -2019 15247 1957
rect 15333 -2019 15367 1957
rect 15491 -2019 15525 1957
rect 15611 -2019 15645 1957
rect 15769 -2019 15803 1957
rect 15889 -2019 15923 1957
rect 16047 -2019 16081 1957
rect 16167 -2019 16201 1957
rect 16325 -2019 16359 1957
rect 16445 -2019 16479 1957
rect 16603 -2019 16637 1957
rect 16723 -2019 16757 1957
rect 16881 -2019 16915 1957
rect 17001 -2019 17035 1957
rect 17159 -2019 17193 1957
rect 17279 -2019 17313 1957
rect 17437 -2019 17471 1957
rect 17557 -2019 17591 1957
rect 17715 -2019 17749 1957
<< metal1 >>
rect -17699 2041 -17607 2047
rect -17699 2007 -17687 2041
rect -17619 2007 -17607 2041
rect -17699 2001 -17607 2007
rect -17421 2041 -17329 2047
rect -17421 2007 -17409 2041
rect -17341 2007 -17329 2041
rect -17421 2001 -17329 2007
rect -17143 2041 -17051 2047
rect -17143 2007 -17131 2041
rect -17063 2007 -17051 2041
rect -17143 2001 -17051 2007
rect -16865 2041 -16773 2047
rect -16865 2007 -16853 2041
rect -16785 2007 -16773 2041
rect -16865 2001 -16773 2007
rect -16587 2041 -16495 2047
rect -16587 2007 -16575 2041
rect -16507 2007 -16495 2041
rect -16587 2001 -16495 2007
rect -16309 2041 -16217 2047
rect -16309 2007 -16297 2041
rect -16229 2007 -16217 2041
rect -16309 2001 -16217 2007
rect -16031 2041 -15939 2047
rect -16031 2007 -16019 2041
rect -15951 2007 -15939 2041
rect -16031 2001 -15939 2007
rect -15753 2041 -15661 2047
rect -15753 2007 -15741 2041
rect -15673 2007 -15661 2041
rect -15753 2001 -15661 2007
rect -15475 2041 -15383 2047
rect -15475 2007 -15463 2041
rect -15395 2007 -15383 2041
rect -15475 2001 -15383 2007
rect -15197 2041 -15105 2047
rect -15197 2007 -15185 2041
rect -15117 2007 -15105 2041
rect -15197 2001 -15105 2007
rect -14919 2041 -14827 2047
rect -14919 2007 -14907 2041
rect -14839 2007 -14827 2041
rect -14919 2001 -14827 2007
rect -14641 2041 -14549 2047
rect -14641 2007 -14629 2041
rect -14561 2007 -14549 2041
rect -14641 2001 -14549 2007
rect -14363 2041 -14271 2047
rect -14363 2007 -14351 2041
rect -14283 2007 -14271 2041
rect -14363 2001 -14271 2007
rect -14085 2041 -13993 2047
rect -14085 2007 -14073 2041
rect -14005 2007 -13993 2041
rect -14085 2001 -13993 2007
rect -13807 2041 -13715 2047
rect -13807 2007 -13795 2041
rect -13727 2007 -13715 2041
rect -13807 2001 -13715 2007
rect -13529 2041 -13437 2047
rect -13529 2007 -13517 2041
rect -13449 2007 -13437 2041
rect -13529 2001 -13437 2007
rect -13251 2041 -13159 2047
rect -13251 2007 -13239 2041
rect -13171 2007 -13159 2041
rect -13251 2001 -13159 2007
rect -12973 2041 -12881 2047
rect -12973 2007 -12961 2041
rect -12893 2007 -12881 2041
rect -12973 2001 -12881 2007
rect -12695 2041 -12603 2047
rect -12695 2007 -12683 2041
rect -12615 2007 -12603 2041
rect -12695 2001 -12603 2007
rect -12417 2041 -12325 2047
rect -12417 2007 -12405 2041
rect -12337 2007 -12325 2041
rect -12417 2001 -12325 2007
rect -12139 2041 -12047 2047
rect -12139 2007 -12127 2041
rect -12059 2007 -12047 2041
rect -12139 2001 -12047 2007
rect -11861 2041 -11769 2047
rect -11861 2007 -11849 2041
rect -11781 2007 -11769 2041
rect -11861 2001 -11769 2007
rect -11583 2041 -11491 2047
rect -11583 2007 -11571 2041
rect -11503 2007 -11491 2041
rect -11583 2001 -11491 2007
rect -11305 2041 -11213 2047
rect -11305 2007 -11293 2041
rect -11225 2007 -11213 2041
rect -11305 2001 -11213 2007
rect -11027 2041 -10935 2047
rect -11027 2007 -11015 2041
rect -10947 2007 -10935 2041
rect -11027 2001 -10935 2007
rect -10749 2041 -10657 2047
rect -10749 2007 -10737 2041
rect -10669 2007 -10657 2041
rect -10749 2001 -10657 2007
rect -10471 2041 -10379 2047
rect -10471 2007 -10459 2041
rect -10391 2007 -10379 2041
rect -10471 2001 -10379 2007
rect -10193 2041 -10101 2047
rect -10193 2007 -10181 2041
rect -10113 2007 -10101 2041
rect -10193 2001 -10101 2007
rect -9915 2041 -9823 2047
rect -9915 2007 -9903 2041
rect -9835 2007 -9823 2041
rect -9915 2001 -9823 2007
rect -9637 2041 -9545 2047
rect -9637 2007 -9625 2041
rect -9557 2007 -9545 2041
rect -9637 2001 -9545 2007
rect -9359 2041 -9267 2047
rect -9359 2007 -9347 2041
rect -9279 2007 -9267 2041
rect -9359 2001 -9267 2007
rect -9081 2041 -8989 2047
rect -9081 2007 -9069 2041
rect -9001 2007 -8989 2041
rect -9081 2001 -8989 2007
rect -8803 2041 -8711 2047
rect -8803 2007 -8791 2041
rect -8723 2007 -8711 2041
rect -8803 2001 -8711 2007
rect -8525 2041 -8433 2047
rect -8525 2007 -8513 2041
rect -8445 2007 -8433 2041
rect -8525 2001 -8433 2007
rect -8247 2041 -8155 2047
rect -8247 2007 -8235 2041
rect -8167 2007 -8155 2041
rect -8247 2001 -8155 2007
rect -7969 2041 -7877 2047
rect -7969 2007 -7957 2041
rect -7889 2007 -7877 2041
rect -7969 2001 -7877 2007
rect -7691 2041 -7599 2047
rect -7691 2007 -7679 2041
rect -7611 2007 -7599 2041
rect -7691 2001 -7599 2007
rect -7413 2041 -7321 2047
rect -7413 2007 -7401 2041
rect -7333 2007 -7321 2041
rect -7413 2001 -7321 2007
rect -7135 2041 -7043 2047
rect -7135 2007 -7123 2041
rect -7055 2007 -7043 2041
rect -7135 2001 -7043 2007
rect -6857 2041 -6765 2047
rect -6857 2007 -6845 2041
rect -6777 2007 -6765 2041
rect -6857 2001 -6765 2007
rect -6579 2041 -6487 2047
rect -6579 2007 -6567 2041
rect -6499 2007 -6487 2041
rect -6579 2001 -6487 2007
rect -6301 2041 -6209 2047
rect -6301 2007 -6289 2041
rect -6221 2007 -6209 2041
rect -6301 2001 -6209 2007
rect -6023 2041 -5931 2047
rect -6023 2007 -6011 2041
rect -5943 2007 -5931 2041
rect -6023 2001 -5931 2007
rect -5745 2041 -5653 2047
rect -5745 2007 -5733 2041
rect -5665 2007 -5653 2041
rect -5745 2001 -5653 2007
rect -5467 2041 -5375 2047
rect -5467 2007 -5455 2041
rect -5387 2007 -5375 2041
rect -5467 2001 -5375 2007
rect -5189 2041 -5097 2047
rect -5189 2007 -5177 2041
rect -5109 2007 -5097 2041
rect -5189 2001 -5097 2007
rect -4911 2041 -4819 2047
rect -4911 2007 -4899 2041
rect -4831 2007 -4819 2041
rect -4911 2001 -4819 2007
rect -4633 2041 -4541 2047
rect -4633 2007 -4621 2041
rect -4553 2007 -4541 2041
rect -4633 2001 -4541 2007
rect -4355 2041 -4263 2047
rect -4355 2007 -4343 2041
rect -4275 2007 -4263 2041
rect -4355 2001 -4263 2007
rect -4077 2041 -3985 2047
rect -4077 2007 -4065 2041
rect -3997 2007 -3985 2041
rect -4077 2001 -3985 2007
rect -3799 2041 -3707 2047
rect -3799 2007 -3787 2041
rect -3719 2007 -3707 2041
rect -3799 2001 -3707 2007
rect -3521 2041 -3429 2047
rect -3521 2007 -3509 2041
rect -3441 2007 -3429 2041
rect -3521 2001 -3429 2007
rect -3243 2041 -3151 2047
rect -3243 2007 -3231 2041
rect -3163 2007 -3151 2041
rect -3243 2001 -3151 2007
rect -2965 2041 -2873 2047
rect -2965 2007 -2953 2041
rect -2885 2007 -2873 2041
rect -2965 2001 -2873 2007
rect -2687 2041 -2595 2047
rect -2687 2007 -2675 2041
rect -2607 2007 -2595 2041
rect -2687 2001 -2595 2007
rect -2409 2041 -2317 2047
rect -2409 2007 -2397 2041
rect -2329 2007 -2317 2041
rect -2409 2001 -2317 2007
rect -2131 2041 -2039 2047
rect -2131 2007 -2119 2041
rect -2051 2007 -2039 2041
rect -2131 2001 -2039 2007
rect -1853 2041 -1761 2047
rect -1853 2007 -1841 2041
rect -1773 2007 -1761 2041
rect -1853 2001 -1761 2007
rect -1575 2041 -1483 2047
rect -1575 2007 -1563 2041
rect -1495 2007 -1483 2041
rect -1575 2001 -1483 2007
rect -1297 2041 -1205 2047
rect -1297 2007 -1285 2041
rect -1217 2007 -1205 2041
rect -1297 2001 -1205 2007
rect -1019 2041 -927 2047
rect -1019 2007 -1007 2041
rect -939 2007 -927 2041
rect -1019 2001 -927 2007
rect -741 2041 -649 2047
rect -741 2007 -729 2041
rect -661 2007 -649 2041
rect -741 2001 -649 2007
rect -463 2041 -371 2047
rect -463 2007 -451 2041
rect -383 2007 -371 2041
rect -463 2001 -371 2007
rect -185 2041 -93 2047
rect -185 2007 -173 2041
rect -105 2007 -93 2041
rect -185 2001 -93 2007
rect 93 2041 185 2047
rect 93 2007 105 2041
rect 173 2007 185 2041
rect 93 2001 185 2007
rect 371 2041 463 2047
rect 371 2007 383 2041
rect 451 2007 463 2041
rect 371 2001 463 2007
rect 649 2041 741 2047
rect 649 2007 661 2041
rect 729 2007 741 2041
rect 649 2001 741 2007
rect 927 2041 1019 2047
rect 927 2007 939 2041
rect 1007 2007 1019 2041
rect 927 2001 1019 2007
rect 1205 2041 1297 2047
rect 1205 2007 1217 2041
rect 1285 2007 1297 2041
rect 1205 2001 1297 2007
rect 1483 2041 1575 2047
rect 1483 2007 1495 2041
rect 1563 2007 1575 2041
rect 1483 2001 1575 2007
rect 1761 2041 1853 2047
rect 1761 2007 1773 2041
rect 1841 2007 1853 2041
rect 1761 2001 1853 2007
rect 2039 2041 2131 2047
rect 2039 2007 2051 2041
rect 2119 2007 2131 2041
rect 2039 2001 2131 2007
rect 2317 2041 2409 2047
rect 2317 2007 2329 2041
rect 2397 2007 2409 2041
rect 2317 2001 2409 2007
rect 2595 2041 2687 2047
rect 2595 2007 2607 2041
rect 2675 2007 2687 2041
rect 2595 2001 2687 2007
rect 2873 2041 2965 2047
rect 2873 2007 2885 2041
rect 2953 2007 2965 2041
rect 2873 2001 2965 2007
rect 3151 2041 3243 2047
rect 3151 2007 3163 2041
rect 3231 2007 3243 2041
rect 3151 2001 3243 2007
rect 3429 2041 3521 2047
rect 3429 2007 3441 2041
rect 3509 2007 3521 2041
rect 3429 2001 3521 2007
rect 3707 2041 3799 2047
rect 3707 2007 3719 2041
rect 3787 2007 3799 2041
rect 3707 2001 3799 2007
rect 3985 2041 4077 2047
rect 3985 2007 3997 2041
rect 4065 2007 4077 2041
rect 3985 2001 4077 2007
rect 4263 2041 4355 2047
rect 4263 2007 4275 2041
rect 4343 2007 4355 2041
rect 4263 2001 4355 2007
rect 4541 2041 4633 2047
rect 4541 2007 4553 2041
rect 4621 2007 4633 2041
rect 4541 2001 4633 2007
rect 4819 2041 4911 2047
rect 4819 2007 4831 2041
rect 4899 2007 4911 2041
rect 4819 2001 4911 2007
rect 5097 2041 5189 2047
rect 5097 2007 5109 2041
rect 5177 2007 5189 2041
rect 5097 2001 5189 2007
rect 5375 2041 5467 2047
rect 5375 2007 5387 2041
rect 5455 2007 5467 2041
rect 5375 2001 5467 2007
rect 5653 2041 5745 2047
rect 5653 2007 5665 2041
rect 5733 2007 5745 2041
rect 5653 2001 5745 2007
rect 5931 2041 6023 2047
rect 5931 2007 5943 2041
rect 6011 2007 6023 2041
rect 5931 2001 6023 2007
rect 6209 2041 6301 2047
rect 6209 2007 6221 2041
rect 6289 2007 6301 2041
rect 6209 2001 6301 2007
rect 6487 2041 6579 2047
rect 6487 2007 6499 2041
rect 6567 2007 6579 2041
rect 6487 2001 6579 2007
rect 6765 2041 6857 2047
rect 6765 2007 6777 2041
rect 6845 2007 6857 2041
rect 6765 2001 6857 2007
rect 7043 2041 7135 2047
rect 7043 2007 7055 2041
rect 7123 2007 7135 2041
rect 7043 2001 7135 2007
rect 7321 2041 7413 2047
rect 7321 2007 7333 2041
rect 7401 2007 7413 2041
rect 7321 2001 7413 2007
rect 7599 2041 7691 2047
rect 7599 2007 7611 2041
rect 7679 2007 7691 2041
rect 7599 2001 7691 2007
rect 7877 2041 7969 2047
rect 7877 2007 7889 2041
rect 7957 2007 7969 2041
rect 7877 2001 7969 2007
rect 8155 2041 8247 2047
rect 8155 2007 8167 2041
rect 8235 2007 8247 2041
rect 8155 2001 8247 2007
rect 8433 2041 8525 2047
rect 8433 2007 8445 2041
rect 8513 2007 8525 2041
rect 8433 2001 8525 2007
rect 8711 2041 8803 2047
rect 8711 2007 8723 2041
rect 8791 2007 8803 2041
rect 8711 2001 8803 2007
rect 8989 2041 9081 2047
rect 8989 2007 9001 2041
rect 9069 2007 9081 2041
rect 8989 2001 9081 2007
rect 9267 2041 9359 2047
rect 9267 2007 9279 2041
rect 9347 2007 9359 2041
rect 9267 2001 9359 2007
rect 9545 2041 9637 2047
rect 9545 2007 9557 2041
rect 9625 2007 9637 2041
rect 9545 2001 9637 2007
rect 9823 2041 9915 2047
rect 9823 2007 9835 2041
rect 9903 2007 9915 2041
rect 9823 2001 9915 2007
rect 10101 2041 10193 2047
rect 10101 2007 10113 2041
rect 10181 2007 10193 2041
rect 10101 2001 10193 2007
rect 10379 2041 10471 2047
rect 10379 2007 10391 2041
rect 10459 2007 10471 2041
rect 10379 2001 10471 2007
rect 10657 2041 10749 2047
rect 10657 2007 10669 2041
rect 10737 2007 10749 2041
rect 10657 2001 10749 2007
rect 10935 2041 11027 2047
rect 10935 2007 10947 2041
rect 11015 2007 11027 2041
rect 10935 2001 11027 2007
rect 11213 2041 11305 2047
rect 11213 2007 11225 2041
rect 11293 2007 11305 2041
rect 11213 2001 11305 2007
rect 11491 2041 11583 2047
rect 11491 2007 11503 2041
rect 11571 2007 11583 2041
rect 11491 2001 11583 2007
rect 11769 2041 11861 2047
rect 11769 2007 11781 2041
rect 11849 2007 11861 2041
rect 11769 2001 11861 2007
rect 12047 2041 12139 2047
rect 12047 2007 12059 2041
rect 12127 2007 12139 2041
rect 12047 2001 12139 2007
rect 12325 2041 12417 2047
rect 12325 2007 12337 2041
rect 12405 2007 12417 2041
rect 12325 2001 12417 2007
rect 12603 2041 12695 2047
rect 12603 2007 12615 2041
rect 12683 2007 12695 2041
rect 12603 2001 12695 2007
rect 12881 2041 12973 2047
rect 12881 2007 12893 2041
rect 12961 2007 12973 2041
rect 12881 2001 12973 2007
rect 13159 2041 13251 2047
rect 13159 2007 13171 2041
rect 13239 2007 13251 2041
rect 13159 2001 13251 2007
rect 13437 2041 13529 2047
rect 13437 2007 13449 2041
rect 13517 2007 13529 2041
rect 13437 2001 13529 2007
rect 13715 2041 13807 2047
rect 13715 2007 13727 2041
rect 13795 2007 13807 2041
rect 13715 2001 13807 2007
rect 13993 2041 14085 2047
rect 13993 2007 14005 2041
rect 14073 2007 14085 2041
rect 13993 2001 14085 2007
rect 14271 2041 14363 2047
rect 14271 2007 14283 2041
rect 14351 2007 14363 2041
rect 14271 2001 14363 2007
rect 14549 2041 14641 2047
rect 14549 2007 14561 2041
rect 14629 2007 14641 2041
rect 14549 2001 14641 2007
rect 14827 2041 14919 2047
rect 14827 2007 14839 2041
rect 14907 2007 14919 2041
rect 14827 2001 14919 2007
rect 15105 2041 15197 2047
rect 15105 2007 15117 2041
rect 15185 2007 15197 2041
rect 15105 2001 15197 2007
rect 15383 2041 15475 2047
rect 15383 2007 15395 2041
rect 15463 2007 15475 2041
rect 15383 2001 15475 2007
rect 15661 2041 15753 2047
rect 15661 2007 15673 2041
rect 15741 2007 15753 2041
rect 15661 2001 15753 2007
rect 15939 2041 16031 2047
rect 15939 2007 15951 2041
rect 16019 2007 16031 2041
rect 15939 2001 16031 2007
rect 16217 2041 16309 2047
rect 16217 2007 16229 2041
rect 16297 2007 16309 2041
rect 16217 2001 16309 2007
rect 16495 2041 16587 2047
rect 16495 2007 16507 2041
rect 16575 2007 16587 2041
rect 16495 2001 16587 2007
rect 16773 2041 16865 2047
rect 16773 2007 16785 2041
rect 16853 2007 16865 2041
rect 16773 2001 16865 2007
rect 17051 2041 17143 2047
rect 17051 2007 17063 2041
rect 17131 2007 17143 2041
rect 17051 2001 17143 2007
rect 17329 2041 17421 2047
rect 17329 2007 17341 2041
rect 17409 2007 17421 2041
rect 17329 2001 17421 2007
rect 17607 2041 17699 2047
rect 17607 2007 17619 2041
rect 17687 2007 17699 2041
rect 17607 2001 17699 2007
rect -17755 1957 -17709 1969
rect -17755 -2019 -17749 1957
rect -17715 -2019 -17709 1957
rect -17755 -2031 -17709 -2019
rect -17597 1957 -17551 1969
rect -17597 -2019 -17591 1957
rect -17557 -2019 -17551 1957
rect -17597 -2031 -17551 -2019
rect -17477 1957 -17431 1969
rect -17477 -2019 -17471 1957
rect -17437 -2019 -17431 1957
rect -17477 -2031 -17431 -2019
rect -17319 1957 -17273 1969
rect -17319 -2019 -17313 1957
rect -17279 -2019 -17273 1957
rect -17319 -2031 -17273 -2019
rect -17199 1957 -17153 1969
rect -17199 -2019 -17193 1957
rect -17159 -2019 -17153 1957
rect -17199 -2031 -17153 -2019
rect -17041 1957 -16995 1969
rect -17041 -2019 -17035 1957
rect -17001 -2019 -16995 1957
rect -17041 -2031 -16995 -2019
rect -16921 1957 -16875 1969
rect -16921 -2019 -16915 1957
rect -16881 -2019 -16875 1957
rect -16921 -2031 -16875 -2019
rect -16763 1957 -16717 1969
rect -16763 -2019 -16757 1957
rect -16723 -2019 -16717 1957
rect -16763 -2031 -16717 -2019
rect -16643 1957 -16597 1969
rect -16643 -2019 -16637 1957
rect -16603 -2019 -16597 1957
rect -16643 -2031 -16597 -2019
rect -16485 1957 -16439 1969
rect -16485 -2019 -16479 1957
rect -16445 -2019 -16439 1957
rect -16485 -2031 -16439 -2019
rect -16365 1957 -16319 1969
rect -16365 -2019 -16359 1957
rect -16325 -2019 -16319 1957
rect -16365 -2031 -16319 -2019
rect -16207 1957 -16161 1969
rect -16207 -2019 -16201 1957
rect -16167 -2019 -16161 1957
rect -16207 -2031 -16161 -2019
rect -16087 1957 -16041 1969
rect -16087 -2019 -16081 1957
rect -16047 -2019 -16041 1957
rect -16087 -2031 -16041 -2019
rect -15929 1957 -15883 1969
rect -15929 -2019 -15923 1957
rect -15889 -2019 -15883 1957
rect -15929 -2031 -15883 -2019
rect -15809 1957 -15763 1969
rect -15809 -2019 -15803 1957
rect -15769 -2019 -15763 1957
rect -15809 -2031 -15763 -2019
rect -15651 1957 -15605 1969
rect -15651 -2019 -15645 1957
rect -15611 -2019 -15605 1957
rect -15651 -2031 -15605 -2019
rect -15531 1957 -15485 1969
rect -15531 -2019 -15525 1957
rect -15491 -2019 -15485 1957
rect -15531 -2031 -15485 -2019
rect -15373 1957 -15327 1969
rect -15373 -2019 -15367 1957
rect -15333 -2019 -15327 1957
rect -15373 -2031 -15327 -2019
rect -15253 1957 -15207 1969
rect -15253 -2019 -15247 1957
rect -15213 -2019 -15207 1957
rect -15253 -2031 -15207 -2019
rect -15095 1957 -15049 1969
rect -15095 -2019 -15089 1957
rect -15055 -2019 -15049 1957
rect -15095 -2031 -15049 -2019
rect -14975 1957 -14929 1969
rect -14975 -2019 -14969 1957
rect -14935 -2019 -14929 1957
rect -14975 -2031 -14929 -2019
rect -14817 1957 -14771 1969
rect -14817 -2019 -14811 1957
rect -14777 -2019 -14771 1957
rect -14817 -2031 -14771 -2019
rect -14697 1957 -14651 1969
rect -14697 -2019 -14691 1957
rect -14657 -2019 -14651 1957
rect -14697 -2031 -14651 -2019
rect -14539 1957 -14493 1969
rect -14539 -2019 -14533 1957
rect -14499 -2019 -14493 1957
rect -14539 -2031 -14493 -2019
rect -14419 1957 -14373 1969
rect -14419 -2019 -14413 1957
rect -14379 -2019 -14373 1957
rect -14419 -2031 -14373 -2019
rect -14261 1957 -14215 1969
rect -14261 -2019 -14255 1957
rect -14221 -2019 -14215 1957
rect -14261 -2031 -14215 -2019
rect -14141 1957 -14095 1969
rect -14141 -2019 -14135 1957
rect -14101 -2019 -14095 1957
rect -14141 -2031 -14095 -2019
rect -13983 1957 -13937 1969
rect -13983 -2019 -13977 1957
rect -13943 -2019 -13937 1957
rect -13983 -2031 -13937 -2019
rect -13863 1957 -13817 1969
rect -13863 -2019 -13857 1957
rect -13823 -2019 -13817 1957
rect -13863 -2031 -13817 -2019
rect -13705 1957 -13659 1969
rect -13705 -2019 -13699 1957
rect -13665 -2019 -13659 1957
rect -13705 -2031 -13659 -2019
rect -13585 1957 -13539 1969
rect -13585 -2019 -13579 1957
rect -13545 -2019 -13539 1957
rect -13585 -2031 -13539 -2019
rect -13427 1957 -13381 1969
rect -13427 -2019 -13421 1957
rect -13387 -2019 -13381 1957
rect -13427 -2031 -13381 -2019
rect -13307 1957 -13261 1969
rect -13307 -2019 -13301 1957
rect -13267 -2019 -13261 1957
rect -13307 -2031 -13261 -2019
rect -13149 1957 -13103 1969
rect -13149 -2019 -13143 1957
rect -13109 -2019 -13103 1957
rect -13149 -2031 -13103 -2019
rect -13029 1957 -12983 1969
rect -13029 -2019 -13023 1957
rect -12989 -2019 -12983 1957
rect -13029 -2031 -12983 -2019
rect -12871 1957 -12825 1969
rect -12871 -2019 -12865 1957
rect -12831 -2019 -12825 1957
rect -12871 -2031 -12825 -2019
rect -12751 1957 -12705 1969
rect -12751 -2019 -12745 1957
rect -12711 -2019 -12705 1957
rect -12751 -2031 -12705 -2019
rect -12593 1957 -12547 1969
rect -12593 -2019 -12587 1957
rect -12553 -2019 -12547 1957
rect -12593 -2031 -12547 -2019
rect -12473 1957 -12427 1969
rect -12473 -2019 -12467 1957
rect -12433 -2019 -12427 1957
rect -12473 -2031 -12427 -2019
rect -12315 1957 -12269 1969
rect -12315 -2019 -12309 1957
rect -12275 -2019 -12269 1957
rect -12315 -2031 -12269 -2019
rect -12195 1957 -12149 1969
rect -12195 -2019 -12189 1957
rect -12155 -2019 -12149 1957
rect -12195 -2031 -12149 -2019
rect -12037 1957 -11991 1969
rect -12037 -2019 -12031 1957
rect -11997 -2019 -11991 1957
rect -12037 -2031 -11991 -2019
rect -11917 1957 -11871 1969
rect -11917 -2019 -11911 1957
rect -11877 -2019 -11871 1957
rect -11917 -2031 -11871 -2019
rect -11759 1957 -11713 1969
rect -11759 -2019 -11753 1957
rect -11719 -2019 -11713 1957
rect -11759 -2031 -11713 -2019
rect -11639 1957 -11593 1969
rect -11639 -2019 -11633 1957
rect -11599 -2019 -11593 1957
rect -11639 -2031 -11593 -2019
rect -11481 1957 -11435 1969
rect -11481 -2019 -11475 1957
rect -11441 -2019 -11435 1957
rect -11481 -2031 -11435 -2019
rect -11361 1957 -11315 1969
rect -11361 -2019 -11355 1957
rect -11321 -2019 -11315 1957
rect -11361 -2031 -11315 -2019
rect -11203 1957 -11157 1969
rect -11203 -2019 -11197 1957
rect -11163 -2019 -11157 1957
rect -11203 -2031 -11157 -2019
rect -11083 1957 -11037 1969
rect -11083 -2019 -11077 1957
rect -11043 -2019 -11037 1957
rect -11083 -2031 -11037 -2019
rect -10925 1957 -10879 1969
rect -10925 -2019 -10919 1957
rect -10885 -2019 -10879 1957
rect -10925 -2031 -10879 -2019
rect -10805 1957 -10759 1969
rect -10805 -2019 -10799 1957
rect -10765 -2019 -10759 1957
rect -10805 -2031 -10759 -2019
rect -10647 1957 -10601 1969
rect -10647 -2019 -10641 1957
rect -10607 -2019 -10601 1957
rect -10647 -2031 -10601 -2019
rect -10527 1957 -10481 1969
rect -10527 -2019 -10521 1957
rect -10487 -2019 -10481 1957
rect -10527 -2031 -10481 -2019
rect -10369 1957 -10323 1969
rect -10369 -2019 -10363 1957
rect -10329 -2019 -10323 1957
rect -10369 -2031 -10323 -2019
rect -10249 1957 -10203 1969
rect -10249 -2019 -10243 1957
rect -10209 -2019 -10203 1957
rect -10249 -2031 -10203 -2019
rect -10091 1957 -10045 1969
rect -10091 -2019 -10085 1957
rect -10051 -2019 -10045 1957
rect -10091 -2031 -10045 -2019
rect -9971 1957 -9925 1969
rect -9971 -2019 -9965 1957
rect -9931 -2019 -9925 1957
rect -9971 -2031 -9925 -2019
rect -9813 1957 -9767 1969
rect -9813 -2019 -9807 1957
rect -9773 -2019 -9767 1957
rect -9813 -2031 -9767 -2019
rect -9693 1957 -9647 1969
rect -9693 -2019 -9687 1957
rect -9653 -2019 -9647 1957
rect -9693 -2031 -9647 -2019
rect -9535 1957 -9489 1969
rect -9535 -2019 -9529 1957
rect -9495 -2019 -9489 1957
rect -9535 -2031 -9489 -2019
rect -9415 1957 -9369 1969
rect -9415 -2019 -9409 1957
rect -9375 -2019 -9369 1957
rect -9415 -2031 -9369 -2019
rect -9257 1957 -9211 1969
rect -9257 -2019 -9251 1957
rect -9217 -2019 -9211 1957
rect -9257 -2031 -9211 -2019
rect -9137 1957 -9091 1969
rect -9137 -2019 -9131 1957
rect -9097 -2019 -9091 1957
rect -9137 -2031 -9091 -2019
rect -8979 1957 -8933 1969
rect -8979 -2019 -8973 1957
rect -8939 -2019 -8933 1957
rect -8979 -2031 -8933 -2019
rect -8859 1957 -8813 1969
rect -8859 -2019 -8853 1957
rect -8819 -2019 -8813 1957
rect -8859 -2031 -8813 -2019
rect -8701 1957 -8655 1969
rect -8701 -2019 -8695 1957
rect -8661 -2019 -8655 1957
rect -8701 -2031 -8655 -2019
rect -8581 1957 -8535 1969
rect -8581 -2019 -8575 1957
rect -8541 -2019 -8535 1957
rect -8581 -2031 -8535 -2019
rect -8423 1957 -8377 1969
rect -8423 -2019 -8417 1957
rect -8383 -2019 -8377 1957
rect -8423 -2031 -8377 -2019
rect -8303 1957 -8257 1969
rect -8303 -2019 -8297 1957
rect -8263 -2019 -8257 1957
rect -8303 -2031 -8257 -2019
rect -8145 1957 -8099 1969
rect -8145 -2019 -8139 1957
rect -8105 -2019 -8099 1957
rect -8145 -2031 -8099 -2019
rect -8025 1957 -7979 1969
rect -8025 -2019 -8019 1957
rect -7985 -2019 -7979 1957
rect -8025 -2031 -7979 -2019
rect -7867 1957 -7821 1969
rect -7867 -2019 -7861 1957
rect -7827 -2019 -7821 1957
rect -7867 -2031 -7821 -2019
rect -7747 1957 -7701 1969
rect -7747 -2019 -7741 1957
rect -7707 -2019 -7701 1957
rect -7747 -2031 -7701 -2019
rect -7589 1957 -7543 1969
rect -7589 -2019 -7583 1957
rect -7549 -2019 -7543 1957
rect -7589 -2031 -7543 -2019
rect -7469 1957 -7423 1969
rect -7469 -2019 -7463 1957
rect -7429 -2019 -7423 1957
rect -7469 -2031 -7423 -2019
rect -7311 1957 -7265 1969
rect -7311 -2019 -7305 1957
rect -7271 -2019 -7265 1957
rect -7311 -2031 -7265 -2019
rect -7191 1957 -7145 1969
rect -7191 -2019 -7185 1957
rect -7151 -2019 -7145 1957
rect -7191 -2031 -7145 -2019
rect -7033 1957 -6987 1969
rect -7033 -2019 -7027 1957
rect -6993 -2019 -6987 1957
rect -7033 -2031 -6987 -2019
rect -6913 1957 -6867 1969
rect -6913 -2019 -6907 1957
rect -6873 -2019 -6867 1957
rect -6913 -2031 -6867 -2019
rect -6755 1957 -6709 1969
rect -6755 -2019 -6749 1957
rect -6715 -2019 -6709 1957
rect -6755 -2031 -6709 -2019
rect -6635 1957 -6589 1969
rect -6635 -2019 -6629 1957
rect -6595 -2019 -6589 1957
rect -6635 -2031 -6589 -2019
rect -6477 1957 -6431 1969
rect -6477 -2019 -6471 1957
rect -6437 -2019 -6431 1957
rect -6477 -2031 -6431 -2019
rect -6357 1957 -6311 1969
rect -6357 -2019 -6351 1957
rect -6317 -2019 -6311 1957
rect -6357 -2031 -6311 -2019
rect -6199 1957 -6153 1969
rect -6199 -2019 -6193 1957
rect -6159 -2019 -6153 1957
rect -6199 -2031 -6153 -2019
rect -6079 1957 -6033 1969
rect -6079 -2019 -6073 1957
rect -6039 -2019 -6033 1957
rect -6079 -2031 -6033 -2019
rect -5921 1957 -5875 1969
rect -5921 -2019 -5915 1957
rect -5881 -2019 -5875 1957
rect -5921 -2031 -5875 -2019
rect -5801 1957 -5755 1969
rect -5801 -2019 -5795 1957
rect -5761 -2019 -5755 1957
rect -5801 -2031 -5755 -2019
rect -5643 1957 -5597 1969
rect -5643 -2019 -5637 1957
rect -5603 -2019 -5597 1957
rect -5643 -2031 -5597 -2019
rect -5523 1957 -5477 1969
rect -5523 -2019 -5517 1957
rect -5483 -2019 -5477 1957
rect -5523 -2031 -5477 -2019
rect -5365 1957 -5319 1969
rect -5365 -2019 -5359 1957
rect -5325 -2019 -5319 1957
rect -5365 -2031 -5319 -2019
rect -5245 1957 -5199 1969
rect -5245 -2019 -5239 1957
rect -5205 -2019 -5199 1957
rect -5245 -2031 -5199 -2019
rect -5087 1957 -5041 1969
rect -5087 -2019 -5081 1957
rect -5047 -2019 -5041 1957
rect -5087 -2031 -5041 -2019
rect -4967 1957 -4921 1969
rect -4967 -2019 -4961 1957
rect -4927 -2019 -4921 1957
rect -4967 -2031 -4921 -2019
rect -4809 1957 -4763 1969
rect -4809 -2019 -4803 1957
rect -4769 -2019 -4763 1957
rect -4809 -2031 -4763 -2019
rect -4689 1957 -4643 1969
rect -4689 -2019 -4683 1957
rect -4649 -2019 -4643 1957
rect -4689 -2031 -4643 -2019
rect -4531 1957 -4485 1969
rect -4531 -2019 -4525 1957
rect -4491 -2019 -4485 1957
rect -4531 -2031 -4485 -2019
rect -4411 1957 -4365 1969
rect -4411 -2019 -4405 1957
rect -4371 -2019 -4365 1957
rect -4411 -2031 -4365 -2019
rect -4253 1957 -4207 1969
rect -4253 -2019 -4247 1957
rect -4213 -2019 -4207 1957
rect -4253 -2031 -4207 -2019
rect -4133 1957 -4087 1969
rect -4133 -2019 -4127 1957
rect -4093 -2019 -4087 1957
rect -4133 -2031 -4087 -2019
rect -3975 1957 -3929 1969
rect -3975 -2019 -3969 1957
rect -3935 -2019 -3929 1957
rect -3975 -2031 -3929 -2019
rect -3855 1957 -3809 1969
rect -3855 -2019 -3849 1957
rect -3815 -2019 -3809 1957
rect -3855 -2031 -3809 -2019
rect -3697 1957 -3651 1969
rect -3697 -2019 -3691 1957
rect -3657 -2019 -3651 1957
rect -3697 -2031 -3651 -2019
rect -3577 1957 -3531 1969
rect -3577 -2019 -3571 1957
rect -3537 -2019 -3531 1957
rect -3577 -2031 -3531 -2019
rect -3419 1957 -3373 1969
rect -3419 -2019 -3413 1957
rect -3379 -2019 -3373 1957
rect -3419 -2031 -3373 -2019
rect -3299 1957 -3253 1969
rect -3299 -2019 -3293 1957
rect -3259 -2019 -3253 1957
rect -3299 -2031 -3253 -2019
rect -3141 1957 -3095 1969
rect -3141 -2019 -3135 1957
rect -3101 -2019 -3095 1957
rect -3141 -2031 -3095 -2019
rect -3021 1957 -2975 1969
rect -3021 -2019 -3015 1957
rect -2981 -2019 -2975 1957
rect -3021 -2031 -2975 -2019
rect -2863 1957 -2817 1969
rect -2863 -2019 -2857 1957
rect -2823 -2019 -2817 1957
rect -2863 -2031 -2817 -2019
rect -2743 1957 -2697 1969
rect -2743 -2019 -2737 1957
rect -2703 -2019 -2697 1957
rect -2743 -2031 -2697 -2019
rect -2585 1957 -2539 1969
rect -2585 -2019 -2579 1957
rect -2545 -2019 -2539 1957
rect -2585 -2031 -2539 -2019
rect -2465 1957 -2419 1969
rect -2465 -2019 -2459 1957
rect -2425 -2019 -2419 1957
rect -2465 -2031 -2419 -2019
rect -2307 1957 -2261 1969
rect -2307 -2019 -2301 1957
rect -2267 -2019 -2261 1957
rect -2307 -2031 -2261 -2019
rect -2187 1957 -2141 1969
rect -2187 -2019 -2181 1957
rect -2147 -2019 -2141 1957
rect -2187 -2031 -2141 -2019
rect -2029 1957 -1983 1969
rect -2029 -2019 -2023 1957
rect -1989 -2019 -1983 1957
rect -2029 -2031 -1983 -2019
rect -1909 1957 -1863 1969
rect -1909 -2019 -1903 1957
rect -1869 -2019 -1863 1957
rect -1909 -2031 -1863 -2019
rect -1751 1957 -1705 1969
rect -1751 -2019 -1745 1957
rect -1711 -2019 -1705 1957
rect -1751 -2031 -1705 -2019
rect -1631 1957 -1585 1969
rect -1631 -2019 -1625 1957
rect -1591 -2019 -1585 1957
rect -1631 -2031 -1585 -2019
rect -1473 1957 -1427 1969
rect -1473 -2019 -1467 1957
rect -1433 -2019 -1427 1957
rect -1473 -2031 -1427 -2019
rect -1353 1957 -1307 1969
rect -1353 -2019 -1347 1957
rect -1313 -2019 -1307 1957
rect -1353 -2031 -1307 -2019
rect -1195 1957 -1149 1969
rect -1195 -2019 -1189 1957
rect -1155 -2019 -1149 1957
rect -1195 -2031 -1149 -2019
rect -1075 1957 -1029 1969
rect -1075 -2019 -1069 1957
rect -1035 -2019 -1029 1957
rect -1075 -2031 -1029 -2019
rect -917 1957 -871 1969
rect -917 -2019 -911 1957
rect -877 -2019 -871 1957
rect -917 -2031 -871 -2019
rect -797 1957 -751 1969
rect -797 -2019 -791 1957
rect -757 -2019 -751 1957
rect -797 -2031 -751 -2019
rect -639 1957 -593 1969
rect -639 -2019 -633 1957
rect -599 -2019 -593 1957
rect -639 -2031 -593 -2019
rect -519 1957 -473 1969
rect -519 -2019 -513 1957
rect -479 -2019 -473 1957
rect -519 -2031 -473 -2019
rect -361 1957 -315 1969
rect -361 -2019 -355 1957
rect -321 -2019 -315 1957
rect -361 -2031 -315 -2019
rect -241 1957 -195 1969
rect -241 -2019 -235 1957
rect -201 -2019 -195 1957
rect -241 -2031 -195 -2019
rect -83 1957 -37 1969
rect -83 -2019 -77 1957
rect -43 -2019 -37 1957
rect -83 -2031 -37 -2019
rect 37 1957 83 1969
rect 37 -2019 43 1957
rect 77 -2019 83 1957
rect 37 -2031 83 -2019
rect 195 1957 241 1969
rect 195 -2019 201 1957
rect 235 -2019 241 1957
rect 195 -2031 241 -2019
rect 315 1957 361 1969
rect 315 -2019 321 1957
rect 355 -2019 361 1957
rect 315 -2031 361 -2019
rect 473 1957 519 1969
rect 473 -2019 479 1957
rect 513 -2019 519 1957
rect 473 -2031 519 -2019
rect 593 1957 639 1969
rect 593 -2019 599 1957
rect 633 -2019 639 1957
rect 593 -2031 639 -2019
rect 751 1957 797 1969
rect 751 -2019 757 1957
rect 791 -2019 797 1957
rect 751 -2031 797 -2019
rect 871 1957 917 1969
rect 871 -2019 877 1957
rect 911 -2019 917 1957
rect 871 -2031 917 -2019
rect 1029 1957 1075 1969
rect 1029 -2019 1035 1957
rect 1069 -2019 1075 1957
rect 1029 -2031 1075 -2019
rect 1149 1957 1195 1969
rect 1149 -2019 1155 1957
rect 1189 -2019 1195 1957
rect 1149 -2031 1195 -2019
rect 1307 1957 1353 1969
rect 1307 -2019 1313 1957
rect 1347 -2019 1353 1957
rect 1307 -2031 1353 -2019
rect 1427 1957 1473 1969
rect 1427 -2019 1433 1957
rect 1467 -2019 1473 1957
rect 1427 -2031 1473 -2019
rect 1585 1957 1631 1969
rect 1585 -2019 1591 1957
rect 1625 -2019 1631 1957
rect 1585 -2031 1631 -2019
rect 1705 1957 1751 1969
rect 1705 -2019 1711 1957
rect 1745 -2019 1751 1957
rect 1705 -2031 1751 -2019
rect 1863 1957 1909 1969
rect 1863 -2019 1869 1957
rect 1903 -2019 1909 1957
rect 1863 -2031 1909 -2019
rect 1983 1957 2029 1969
rect 1983 -2019 1989 1957
rect 2023 -2019 2029 1957
rect 1983 -2031 2029 -2019
rect 2141 1957 2187 1969
rect 2141 -2019 2147 1957
rect 2181 -2019 2187 1957
rect 2141 -2031 2187 -2019
rect 2261 1957 2307 1969
rect 2261 -2019 2267 1957
rect 2301 -2019 2307 1957
rect 2261 -2031 2307 -2019
rect 2419 1957 2465 1969
rect 2419 -2019 2425 1957
rect 2459 -2019 2465 1957
rect 2419 -2031 2465 -2019
rect 2539 1957 2585 1969
rect 2539 -2019 2545 1957
rect 2579 -2019 2585 1957
rect 2539 -2031 2585 -2019
rect 2697 1957 2743 1969
rect 2697 -2019 2703 1957
rect 2737 -2019 2743 1957
rect 2697 -2031 2743 -2019
rect 2817 1957 2863 1969
rect 2817 -2019 2823 1957
rect 2857 -2019 2863 1957
rect 2817 -2031 2863 -2019
rect 2975 1957 3021 1969
rect 2975 -2019 2981 1957
rect 3015 -2019 3021 1957
rect 2975 -2031 3021 -2019
rect 3095 1957 3141 1969
rect 3095 -2019 3101 1957
rect 3135 -2019 3141 1957
rect 3095 -2031 3141 -2019
rect 3253 1957 3299 1969
rect 3253 -2019 3259 1957
rect 3293 -2019 3299 1957
rect 3253 -2031 3299 -2019
rect 3373 1957 3419 1969
rect 3373 -2019 3379 1957
rect 3413 -2019 3419 1957
rect 3373 -2031 3419 -2019
rect 3531 1957 3577 1969
rect 3531 -2019 3537 1957
rect 3571 -2019 3577 1957
rect 3531 -2031 3577 -2019
rect 3651 1957 3697 1969
rect 3651 -2019 3657 1957
rect 3691 -2019 3697 1957
rect 3651 -2031 3697 -2019
rect 3809 1957 3855 1969
rect 3809 -2019 3815 1957
rect 3849 -2019 3855 1957
rect 3809 -2031 3855 -2019
rect 3929 1957 3975 1969
rect 3929 -2019 3935 1957
rect 3969 -2019 3975 1957
rect 3929 -2031 3975 -2019
rect 4087 1957 4133 1969
rect 4087 -2019 4093 1957
rect 4127 -2019 4133 1957
rect 4087 -2031 4133 -2019
rect 4207 1957 4253 1969
rect 4207 -2019 4213 1957
rect 4247 -2019 4253 1957
rect 4207 -2031 4253 -2019
rect 4365 1957 4411 1969
rect 4365 -2019 4371 1957
rect 4405 -2019 4411 1957
rect 4365 -2031 4411 -2019
rect 4485 1957 4531 1969
rect 4485 -2019 4491 1957
rect 4525 -2019 4531 1957
rect 4485 -2031 4531 -2019
rect 4643 1957 4689 1969
rect 4643 -2019 4649 1957
rect 4683 -2019 4689 1957
rect 4643 -2031 4689 -2019
rect 4763 1957 4809 1969
rect 4763 -2019 4769 1957
rect 4803 -2019 4809 1957
rect 4763 -2031 4809 -2019
rect 4921 1957 4967 1969
rect 4921 -2019 4927 1957
rect 4961 -2019 4967 1957
rect 4921 -2031 4967 -2019
rect 5041 1957 5087 1969
rect 5041 -2019 5047 1957
rect 5081 -2019 5087 1957
rect 5041 -2031 5087 -2019
rect 5199 1957 5245 1969
rect 5199 -2019 5205 1957
rect 5239 -2019 5245 1957
rect 5199 -2031 5245 -2019
rect 5319 1957 5365 1969
rect 5319 -2019 5325 1957
rect 5359 -2019 5365 1957
rect 5319 -2031 5365 -2019
rect 5477 1957 5523 1969
rect 5477 -2019 5483 1957
rect 5517 -2019 5523 1957
rect 5477 -2031 5523 -2019
rect 5597 1957 5643 1969
rect 5597 -2019 5603 1957
rect 5637 -2019 5643 1957
rect 5597 -2031 5643 -2019
rect 5755 1957 5801 1969
rect 5755 -2019 5761 1957
rect 5795 -2019 5801 1957
rect 5755 -2031 5801 -2019
rect 5875 1957 5921 1969
rect 5875 -2019 5881 1957
rect 5915 -2019 5921 1957
rect 5875 -2031 5921 -2019
rect 6033 1957 6079 1969
rect 6033 -2019 6039 1957
rect 6073 -2019 6079 1957
rect 6033 -2031 6079 -2019
rect 6153 1957 6199 1969
rect 6153 -2019 6159 1957
rect 6193 -2019 6199 1957
rect 6153 -2031 6199 -2019
rect 6311 1957 6357 1969
rect 6311 -2019 6317 1957
rect 6351 -2019 6357 1957
rect 6311 -2031 6357 -2019
rect 6431 1957 6477 1969
rect 6431 -2019 6437 1957
rect 6471 -2019 6477 1957
rect 6431 -2031 6477 -2019
rect 6589 1957 6635 1969
rect 6589 -2019 6595 1957
rect 6629 -2019 6635 1957
rect 6589 -2031 6635 -2019
rect 6709 1957 6755 1969
rect 6709 -2019 6715 1957
rect 6749 -2019 6755 1957
rect 6709 -2031 6755 -2019
rect 6867 1957 6913 1969
rect 6867 -2019 6873 1957
rect 6907 -2019 6913 1957
rect 6867 -2031 6913 -2019
rect 6987 1957 7033 1969
rect 6987 -2019 6993 1957
rect 7027 -2019 7033 1957
rect 6987 -2031 7033 -2019
rect 7145 1957 7191 1969
rect 7145 -2019 7151 1957
rect 7185 -2019 7191 1957
rect 7145 -2031 7191 -2019
rect 7265 1957 7311 1969
rect 7265 -2019 7271 1957
rect 7305 -2019 7311 1957
rect 7265 -2031 7311 -2019
rect 7423 1957 7469 1969
rect 7423 -2019 7429 1957
rect 7463 -2019 7469 1957
rect 7423 -2031 7469 -2019
rect 7543 1957 7589 1969
rect 7543 -2019 7549 1957
rect 7583 -2019 7589 1957
rect 7543 -2031 7589 -2019
rect 7701 1957 7747 1969
rect 7701 -2019 7707 1957
rect 7741 -2019 7747 1957
rect 7701 -2031 7747 -2019
rect 7821 1957 7867 1969
rect 7821 -2019 7827 1957
rect 7861 -2019 7867 1957
rect 7821 -2031 7867 -2019
rect 7979 1957 8025 1969
rect 7979 -2019 7985 1957
rect 8019 -2019 8025 1957
rect 7979 -2031 8025 -2019
rect 8099 1957 8145 1969
rect 8099 -2019 8105 1957
rect 8139 -2019 8145 1957
rect 8099 -2031 8145 -2019
rect 8257 1957 8303 1969
rect 8257 -2019 8263 1957
rect 8297 -2019 8303 1957
rect 8257 -2031 8303 -2019
rect 8377 1957 8423 1969
rect 8377 -2019 8383 1957
rect 8417 -2019 8423 1957
rect 8377 -2031 8423 -2019
rect 8535 1957 8581 1969
rect 8535 -2019 8541 1957
rect 8575 -2019 8581 1957
rect 8535 -2031 8581 -2019
rect 8655 1957 8701 1969
rect 8655 -2019 8661 1957
rect 8695 -2019 8701 1957
rect 8655 -2031 8701 -2019
rect 8813 1957 8859 1969
rect 8813 -2019 8819 1957
rect 8853 -2019 8859 1957
rect 8813 -2031 8859 -2019
rect 8933 1957 8979 1969
rect 8933 -2019 8939 1957
rect 8973 -2019 8979 1957
rect 8933 -2031 8979 -2019
rect 9091 1957 9137 1969
rect 9091 -2019 9097 1957
rect 9131 -2019 9137 1957
rect 9091 -2031 9137 -2019
rect 9211 1957 9257 1969
rect 9211 -2019 9217 1957
rect 9251 -2019 9257 1957
rect 9211 -2031 9257 -2019
rect 9369 1957 9415 1969
rect 9369 -2019 9375 1957
rect 9409 -2019 9415 1957
rect 9369 -2031 9415 -2019
rect 9489 1957 9535 1969
rect 9489 -2019 9495 1957
rect 9529 -2019 9535 1957
rect 9489 -2031 9535 -2019
rect 9647 1957 9693 1969
rect 9647 -2019 9653 1957
rect 9687 -2019 9693 1957
rect 9647 -2031 9693 -2019
rect 9767 1957 9813 1969
rect 9767 -2019 9773 1957
rect 9807 -2019 9813 1957
rect 9767 -2031 9813 -2019
rect 9925 1957 9971 1969
rect 9925 -2019 9931 1957
rect 9965 -2019 9971 1957
rect 9925 -2031 9971 -2019
rect 10045 1957 10091 1969
rect 10045 -2019 10051 1957
rect 10085 -2019 10091 1957
rect 10045 -2031 10091 -2019
rect 10203 1957 10249 1969
rect 10203 -2019 10209 1957
rect 10243 -2019 10249 1957
rect 10203 -2031 10249 -2019
rect 10323 1957 10369 1969
rect 10323 -2019 10329 1957
rect 10363 -2019 10369 1957
rect 10323 -2031 10369 -2019
rect 10481 1957 10527 1969
rect 10481 -2019 10487 1957
rect 10521 -2019 10527 1957
rect 10481 -2031 10527 -2019
rect 10601 1957 10647 1969
rect 10601 -2019 10607 1957
rect 10641 -2019 10647 1957
rect 10601 -2031 10647 -2019
rect 10759 1957 10805 1969
rect 10759 -2019 10765 1957
rect 10799 -2019 10805 1957
rect 10759 -2031 10805 -2019
rect 10879 1957 10925 1969
rect 10879 -2019 10885 1957
rect 10919 -2019 10925 1957
rect 10879 -2031 10925 -2019
rect 11037 1957 11083 1969
rect 11037 -2019 11043 1957
rect 11077 -2019 11083 1957
rect 11037 -2031 11083 -2019
rect 11157 1957 11203 1969
rect 11157 -2019 11163 1957
rect 11197 -2019 11203 1957
rect 11157 -2031 11203 -2019
rect 11315 1957 11361 1969
rect 11315 -2019 11321 1957
rect 11355 -2019 11361 1957
rect 11315 -2031 11361 -2019
rect 11435 1957 11481 1969
rect 11435 -2019 11441 1957
rect 11475 -2019 11481 1957
rect 11435 -2031 11481 -2019
rect 11593 1957 11639 1969
rect 11593 -2019 11599 1957
rect 11633 -2019 11639 1957
rect 11593 -2031 11639 -2019
rect 11713 1957 11759 1969
rect 11713 -2019 11719 1957
rect 11753 -2019 11759 1957
rect 11713 -2031 11759 -2019
rect 11871 1957 11917 1969
rect 11871 -2019 11877 1957
rect 11911 -2019 11917 1957
rect 11871 -2031 11917 -2019
rect 11991 1957 12037 1969
rect 11991 -2019 11997 1957
rect 12031 -2019 12037 1957
rect 11991 -2031 12037 -2019
rect 12149 1957 12195 1969
rect 12149 -2019 12155 1957
rect 12189 -2019 12195 1957
rect 12149 -2031 12195 -2019
rect 12269 1957 12315 1969
rect 12269 -2019 12275 1957
rect 12309 -2019 12315 1957
rect 12269 -2031 12315 -2019
rect 12427 1957 12473 1969
rect 12427 -2019 12433 1957
rect 12467 -2019 12473 1957
rect 12427 -2031 12473 -2019
rect 12547 1957 12593 1969
rect 12547 -2019 12553 1957
rect 12587 -2019 12593 1957
rect 12547 -2031 12593 -2019
rect 12705 1957 12751 1969
rect 12705 -2019 12711 1957
rect 12745 -2019 12751 1957
rect 12705 -2031 12751 -2019
rect 12825 1957 12871 1969
rect 12825 -2019 12831 1957
rect 12865 -2019 12871 1957
rect 12825 -2031 12871 -2019
rect 12983 1957 13029 1969
rect 12983 -2019 12989 1957
rect 13023 -2019 13029 1957
rect 12983 -2031 13029 -2019
rect 13103 1957 13149 1969
rect 13103 -2019 13109 1957
rect 13143 -2019 13149 1957
rect 13103 -2031 13149 -2019
rect 13261 1957 13307 1969
rect 13261 -2019 13267 1957
rect 13301 -2019 13307 1957
rect 13261 -2031 13307 -2019
rect 13381 1957 13427 1969
rect 13381 -2019 13387 1957
rect 13421 -2019 13427 1957
rect 13381 -2031 13427 -2019
rect 13539 1957 13585 1969
rect 13539 -2019 13545 1957
rect 13579 -2019 13585 1957
rect 13539 -2031 13585 -2019
rect 13659 1957 13705 1969
rect 13659 -2019 13665 1957
rect 13699 -2019 13705 1957
rect 13659 -2031 13705 -2019
rect 13817 1957 13863 1969
rect 13817 -2019 13823 1957
rect 13857 -2019 13863 1957
rect 13817 -2031 13863 -2019
rect 13937 1957 13983 1969
rect 13937 -2019 13943 1957
rect 13977 -2019 13983 1957
rect 13937 -2031 13983 -2019
rect 14095 1957 14141 1969
rect 14095 -2019 14101 1957
rect 14135 -2019 14141 1957
rect 14095 -2031 14141 -2019
rect 14215 1957 14261 1969
rect 14215 -2019 14221 1957
rect 14255 -2019 14261 1957
rect 14215 -2031 14261 -2019
rect 14373 1957 14419 1969
rect 14373 -2019 14379 1957
rect 14413 -2019 14419 1957
rect 14373 -2031 14419 -2019
rect 14493 1957 14539 1969
rect 14493 -2019 14499 1957
rect 14533 -2019 14539 1957
rect 14493 -2031 14539 -2019
rect 14651 1957 14697 1969
rect 14651 -2019 14657 1957
rect 14691 -2019 14697 1957
rect 14651 -2031 14697 -2019
rect 14771 1957 14817 1969
rect 14771 -2019 14777 1957
rect 14811 -2019 14817 1957
rect 14771 -2031 14817 -2019
rect 14929 1957 14975 1969
rect 14929 -2019 14935 1957
rect 14969 -2019 14975 1957
rect 14929 -2031 14975 -2019
rect 15049 1957 15095 1969
rect 15049 -2019 15055 1957
rect 15089 -2019 15095 1957
rect 15049 -2031 15095 -2019
rect 15207 1957 15253 1969
rect 15207 -2019 15213 1957
rect 15247 -2019 15253 1957
rect 15207 -2031 15253 -2019
rect 15327 1957 15373 1969
rect 15327 -2019 15333 1957
rect 15367 -2019 15373 1957
rect 15327 -2031 15373 -2019
rect 15485 1957 15531 1969
rect 15485 -2019 15491 1957
rect 15525 -2019 15531 1957
rect 15485 -2031 15531 -2019
rect 15605 1957 15651 1969
rect 15605 -2019 15611 1957
rect 15645 -2019 15651 1957
rect 15605 -2031 15651 -2019
rect 15763 1957 15809 1969
rect 15763 -2019 15769 1957
rect 15803 -2019 15809 1957
rect 15763 -2031 15809 -2019
rect 15883 1957 15929 1969
rect 15883 -2019 15889 1957
rect 15923 -2019 15929 1957
rect 15883 -2031 15929 -2019
rect 16041 1957 16087 1969
rect 16041 -2019 16047 1957
rect 16081 -2019 16087 1957
rect 16041 -2031 16087 -2019
rect 16161 1957 16207 1969
rect 16161 -2019 16167 1957
rect 16201 -2019 16207 1957
rect 16161 -2031 16207 -2019
rect 16319 1957 16365 1969
rect 16319 -2019 16325 1957
rect 16359 -2019 16365 1957
rect 16319 -2031 16365 -2019
rect 16439 1957 16485 1969
rect 16439 -2019 16445 1957
rect 16479 -2019 16485 1957
rect 16439 -2031 16485 -2019
rect 16597 1957 16643 1969
rect 16597 -2019 16603 1957
rect 16637 -2019 16643 1957
rect 16597 -2031 16643 -2019
rect 16717 1957 16763 1969
rect 16717 -2019 16723 1957
rect 16757 -2019 16763 1957
rect 16717 -2031 16763 -2019
rect 16875 1957 16921 1969
rect 16875 -2019 16881 1957
rect 16915 -2019 16921 1957
rect 16875 -2031 16921 -2019
rect 16995 1957 17041 1969
rect 16995 -2019 17001 1957
rect 17035 -2019 17041 1957
rect 16995 -2031 17041 -2019
rect 17153 1957 17199 1969
rect 17153 -2019 17159 1957
rect 17193 -2019 17199 1957
rect 17153 -2031 17199 -2019
rect 17273 1957 17319 1969
rect 17273 -2019 17279 1957
rect 17313 -2019 17319 1957
rect 17273 -2031 17319 -2019
rect 17431 1957 17477 1969
rect 17431 -2019 17437 1957
rect 17471 -2019 17477 1957
rect 17431 -2031 17477 -2019
rect 17551 1957 17597 1969
rect 17551 -2019 17557 1957
rect 17591 -2019 17597 1957
rect 17551 -2031 17597 -2019
rect 17709 1957 17755 1969
rect 17709 -2019 17715 1957
rect 17749 -2019 17755 1957
rect 17709 -2031 17755 -2019
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 20.0 l 0.5 m 1 nf 128 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
