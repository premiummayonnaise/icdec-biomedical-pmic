magic
tech sky130A
magscale 1 2
timestamp 1769135993
<< nwell >>
rect -1940 -259 1940 293
<< pmos >>
rect -1846 -159 -1696 231
rect -1524 -159 -1374 231
rect -1202 -159 -1052 231
rect -880 -159 -730 231
rect -558 -159 -408 231
rect -236 -159 -86 231
rect 86 -159 236 231
rect 408 -159 558 231
rect 730 -159 880 231
rect 1052 -159 1202 231
rect 1374 -159 1524 231
rect 1696 -159 1846 231
<< pdiff >>
rect -1904 219 -1846 231
rect -1904 -147 -1892 219
rect -1858 -147 -1846 219
rect -1904 -159 -1846 -147
rect -1696 219 -1638 231
rect -1696 -147 -1684 219
rect -1650 -147 -1638 219
rect -1696 -159 -1638 -147
rect -1582 219 -1524 231
rect -1582 -147 -1570 219
rect -1536 -147 -1524 219
rect -1582 -159 -1524 -147
rect -1374 219 -1316 231
rect -1374 -147 -1362 219
rect -1328 -147 -1316 219
rect -1374 -159 -1316 -147
rect -1260 219 -1202 231
rect -1260 -147 -1248 219
rect -1214 -147 -1202 219
rect -1260 -159 -1202 -147
rect -1052 219 -994 231
rect -1052 -147 -1040 219
rect -1006 -147 -994 219
rect -1052 -159 -994 -147
rect -938 219 -880 231
rect -938 -147 -926 219
rect -892 -147 -880 219
rect -938 -159 -880 -147
rect -730 219 -672 231
rect -730 -147 -718 219
rect -684 -147 -672 219
rect -730 -159 -672 -147
rect -616 219 -558 231
rect -616 -147 -604 219
rect -570 -147 -558 219
rect -616 -159 -558 -147
rect -408 219 -350 231
rect -408 -147 -396 219
rect -362 -147 -350 219
rect -408 -159 -350 -147
rect -294 219 -236 231
rect -294 -147 -282 219
rect -248 -147 -236 219
rect -294 -159 -236 -147
rect -86 219 -28 231
rect -86 -147 -74 219
rect -40 -147 -28 219
rect -86 -159 -28 -147
rect 28 219 86 231
rect 28 -147 40 219
rect 74 -147 86 219
rect 28 -159 86 -147
rect 236 219 294 231
rect 236 -147 248 219
rect 282 -147 294 219
rect 236 -159 294 -147
rect 350 219 408 231
rect 350 -147 362 219
rect 396 -147 408 219
rect 350 -159 408 -147
rect 558 219 616 231
rect 558 -147 570 219
rect 604 -147 616 219
rect 558 -159 616 -147
rect 672 219 730 231
rect 672 -147 684 219
rect 718 -147 730 219
rect 672 -159 730 -147
rect 880 219 938 231
rect 880 -147 892 219
rect 926 -147 938 219
rect 880 -159 938 -147
rect 994 219 1052 231
rect 994 -147 1006 219
rect 1040 -147 1052 219
rect 994 -159 1052 -147
rect 1202 219 1260 231
rect 1202 -147 1214 219
rect 1248 -147 1260 219
rect 1202 -159 1260 -147
rect 1316 219 1374 231
rect 1316 -147 1328 219
rect 1362 -147 1374 219
rect 1316 -159 1374 -147
rect 1524 219 1582 231
rect 1524 -147 1536 219
rect 1570 -147 1582 219
rect 1524 -159 1582 -147
rect 1638 219 1696 231
rect 1638 -147 1650 219
rect 1684 -147 1696 219
rect 1638 -159 1696 -147
rect 1846 219 1904 231
rect 1846 -147 1858 219
rect 1892 -147 1904 219
rect 1846 -159 1904 -147
<< pdiffc >>
rect -1892 -147 -1858 219
rect -1684 -147 -1650 219
rect -1570 -147 -1536 219
rect -1362 -147 -1328 219
rect -1248 -147 -1214 219
rect -1040 -147 -1006 219
rect -926 -147 -892 219
rect -718 -147 -684 219
rect -604 -147 -570 219
rect -396 -147 -362 219
rect -282 -147 -248 219
rect -74 -147 -40 219
rect 40 -147 74 219
rect 248 -147 282 219
rect 362 -147 396 219
rect 570 -147 604 219
rect 684 -147 718 219
rect 892 -147 926 219
rect 1006 -147 1040 219
rect 1214 -147 1248 219
rect 1328 -147 1362 219
rect 1536 -147 1570 219
rect 1650 -147 1684 219
rect 1858 -147 1892 219
<< poly >>
rect -1846 231 -1696 257
rect -1524 231 -1374 257
rect -1202 231 -1052 257
rect -880 231 -730 257
rect -558 231 -408 257
rect -236 231 -86 257
rect 86 231 236 257
rect 408 231 558 257
rect 730 231 880 257
rect 1052 231 1202 257
rect 1374 231 1524 257
rect 1696 231 1846 257
rect -1846 -206 -1696 -159
rect -1846 -240 -1830 -206
rect -1712 -240 -1696 -206
rect -1846 -256 -1696 -240
rect -1524 -206 -1374 -159
rect -1524 -240 -1508 -206
rect -1390 -240 -1374 -206
rect -1524 -256 -1374 -240
rect -1202 -206 -1052 -159
rect -1202 -240 -1186 -206
rect -1068 -240 -1052 -206
rect -1202 -256 -1052 -240
rect -880 -206 -730 -159
rect -880 -240 -864 -206
rect -746 -240 -730 -206
rect -880 -256 -730 -240
rect -558 -206 -408 -159
rect -558 -240 -542 -206
rect -424 -240 -408 -206
rect -558 -256 -408 -240
rect -236 -206 -86 -159
rect -236 -240 -220 -206
rect -102 -240 -86 -206
rect -236 -256 -86 -240
rect 86 -206 236 -159
rect 86 -240 102 -206
rect 220 -240 236 -206
rect 86 -256 236 -240
rect 408 -206 558 -159
rect 408 -240 424 -206
rect 542 -240 558 -206
rect 408 -256 558 -240
rect 730 -206 880 -159
rect 730 -240 746 -206
rect 864 -240 880 -206
rect 730 -256 880 -240
rect 1052 -206 1202 -159
rect 1052 -240 1068 -206
rect 1186 -240 1202 -206
rect 1052 -256 1202 -240
rect 1374 -206 1524 -159
rect 1374 -240 1390 -206
rect 1508 -240 1524 -206
rect 1374 -256 1524 -240
rect 1696 -206 1846 -159
rect 1696 -240 1712 -206
rect 1830 -240 1846 -206
rect 1696 -256 1846 -240
<< polycont >>
rect -1830 -240 -1712 -206
rect -1508 -240 -1390 -206
rect -1186 -240 -1068 -206
rect -864 -240 -746 -206
rect -542 -240 -424 -206
rect -220 -240 -102 -206
rect 102 -240 220 -206
rect 424 -240 542 -206
rect 746 -240 864 -206
rect 1068 -240 1186 -206
rect 1390 -240 1508 -206
rect 1712 -240 1830 -206
<< locali >>
rect -1892 219 -1858 235
rect -1892 -163 -1858 -147
rect -1684 219 -1650 235
rect -1684 -163 -1650 -147
rect -1570 219 -1536 235
rect -1570 -163 -1536 -147
rect -1362 219 -1328 235
rect -1362 -163 -1328 -147
rect -1248 219 -1214 235
rect -1248 -163 -1214 -147
rect -1040 219 -1006 235
rect -1040 -163 -1006 -147
rect -926 219 -892 235
rect -926 -163 -892 -147
rect -718 219 -684 235
rect -718 -163 -684 -147
rect -604 219 -570 235
rect -604 -163 -570 -147
rect -396 219 -362 235
rect -396 -163 -362 -147
rect -282 219 -248 235
rect -282 -163 -248 -147
rect -74 219 -40 235
rect -74 -163 -40 -147
rect 40 219 74 235
rect 40 -163 74 -147
rect 248 219 282 235
rect 248 -163 282 -147
rect 362 219 396 235
rect 362 -163 396 -147
rect 570 219 604 235
rect 570 -163 604 -147
rect 684 219 718 235
rect 684 -163 718 -147
rect 892 219 926 235
rect 892 -163 926 -147
rect 1006 219 1040 235
rect 1006 -163 1040 -147
rect 1214 219 1248 235
rect 1214 -163 1248 -147
rect 1328 219 1362 235
rect 1328 -163 1362 -147
rect 1536 219 1570 235
rect 1536 -163 1570 -147
rect 1650 219 1684 235
rect 1650 -163 1684 -147
rect 1858 219 1892 235
rect 1858 -163 1892 -147
rect -1846 -240 -1830 -206
rect -1712 -240 -1696 -206
rect -1524 -240 -1508 -206
rect -1390 -240 -1374 -206
rect -1202 -240 -1186 -206
rect -1068 -240 -1052 -206
rect -880 -240 -864 -206
rect -746 -240 -730 -206
rect -558 -240 -542 -206
rect -424 -240 -408 -206
rect -236 -240 -220 -206
rect -102 -240 -86 -206
rect 86 -240 102 -206
rect 220 -240 236 -206
rect 408 -240 424 -206
rect 542 -240 558 -206
rect 730 -240 746 -206
rect 864 -240 880 -206
rect 1052 -240 1068 -206
rect 1186 -240 1202 -206
rect 1374 -240 1390 -206
rect 1508 -240 1524 -206
rect 1696 -240 1712 -206
rect 1830 -240 1846 -206
<< viali >>
rect -1892 -147 -1858 219
rect -1684 -147 -1650 219
rect -1570 -147 -1536 219
rect -1362 -147 -1328 219
rect -1248 -147 -1214 219
rect -1040 -147 -1006 219
rect -926 -147 -892 219
rect -718 -147 -684 219
rect -604 -147 -570 219
rect -396 -147 -362 219
rect -282 -147 -248 219
rect -74 -147 -40 219
rect 40 -147 74 219
rect 248 -147 282 219
rect 362 -147 396 219
rect 570 -147 604 219
rect 684 -147 718 219
rect 892 -147 926 219
rect 1006 -147 1040 219
rect 1214 -147 1248 219
rect 1328 -147 1362 219
rect 1536 -147 1570 219
rect 1650 -147 1684 219
rect 1858 -147 1892 219
rect -1830 -240 -1712 -206
rect -1508 -240 -1390 -206
rect -1186 -240 -1068 -206
rect -864 -240 -746 -206
rect -542 -240 -424 -206
rect -220 -240 -102 -206
rect 102 -240 220 -206
rect 424 -240 542 -206
rect 746 -240 864 -206
rect 1068 -240 1186 -206
rect 1390 -240 1508 -206
rect 1712 -240 1830 -206
<< metal1 >>
rect -1898 219 -1852 231
rect -1898 -147 -1892 219
rect -1858 -147 -1852 219
rect -1898 -159 -1852 -147
rect -1690 219 -1644 231
rect -1690 -147 -1684 219
rect -1650 -147 -1644 219
rect -1690 -159 -1644 -147
rect -1576 219 -1530 231
rect -1576 -147 -1570 219
rect -1536 -147 -1530 219
rect -1576 -159 -1530 -147
rect -1368 219 -1322 231
rect -1368 -147 -1362 219
rect -1328 -147 -1322 219
rect -1368 -159 -1322 -147
rect -1254 219 -1208 231
rect -1254 -147 -1248 219
rect -1214 -147 -1208 219
rect -1254 -159 -1208 -147
rect -1046 219 -1000 231
rect -1046 -147 -1040 219
rect -1006 -147 -1000 219
rect -1046 -159 -1000 -147
rect -932 219 -886 231
rect -932 -147 -926 219
rect -892 -147 -886 219
rect -932 -159 -886 -147
rect -724 219 -678 231
rect -724 -147 -718 219
rect -684 -147 -678 219
rect -724 -159 -678 -147
rect -610 219 -564 231
rect -610 -147 -604 219
rect -570 -147 -564 219
rect -610 -159 -564 -147
rect -402 219 -356 231
rect -402 -147 -396 219
rect -362 -147 -356 219
rect -402 -159 -356 -147
rect -288 219 -242 231
rect -288 -147 -282 219
rect -248 -147 -242 219
rect -288 -159 -242 -147
rect -80 219 -34 231
rect -80 -147 -74 219
rect -40 -147 -34 219
rect -80 -159 -34 -147
rect 34 219 80 231
rect 34 -147 40 219
rect 74 -147 80 219
rect 34 -159 80 -147
rect 242 219 288 231
rect 242 -147 248 219
rect 282 -147 288 219
rect 242 -159 288 -147
rect 356 219 402 231
rect 356 -147 362 219
rect 396 -147 402 219
rect 356 -159 402 -147
rect 564 219 610 231
rect 564 -147 570 219
rect 604 -147 610 219
rect 564 -159 610 -147
rect 678 219 724 231
rect 678 -147 684 219
rect 718 -147 724 219
rect 678 -159 724 -147
rect 886 219 932 231
rect 886 -147 892 219
rect 926 -147 932 219
rect 886 -159 932 -147
rect 1000 219 1046 231
rect 1000 -147 1006 219
rect 1040 -147 1046 219
rect 1000 -159 1046 -147
rect 1208 219 1254 231
rect 1208 -147 1214 219
rect 1248 -147 1254 219
rect 1208 -159 1254 -147
rect 1322 219 1368 231
rect 1322 -147 1328 219
rect 1362 -147 1368 219
rect 1322 -159 1368 -147
rect 1530 219 1576 231
rect 1530 -147 1536 219
rect 1570 -147 1576 219
rect 1530 -159 1576 -147
rect 1644 219 1690 231
rect 1644 -147 1650 219
rect 1684 -147 1690 219
rect 1644 -159 1690 -147
rect 1852 219 1898 231
rect 1852 -147 1858 219
rect 1892 -147 1898 219
rect 1852 -159 1898 -147
rect -1842 -206 -1700 -200
rect -1842 -240 -1830 -206
rect -1712 -240 -1700 -206
rect -1842 -246 -1700 -240
rect -1520 -206 -1378 -200
rect -1520 -240 -1508 -206
rect -1390 -240 -1378 -206
rect -1520 -246 -1378 -240
rect -1198 -206 -1056 -200
rect -1198 -240 -1186 -206
rect -1068 -240 -1056 -206
rect -1198 -246 -1056 -240
rect -876 -206 -734 -200
rect -876 -240 -864 -206
rect -746 -240 -734 -206
rect -876 -246 -734 -240
rect -554 -206 -412 -200
rect -554 -240 -542 -206
rect -424 -240 -412 -206
rect -554 -246 -412 -240
rect -232 -206 -90 -200
rect -232 -240 -220 -206
rect -102 -240 -90 -206
rect -232 -246 -90 -240
rect 90 -206 232 -200
rect 90 -240 102 -206
rect 220 -240 232 -206
rect 90 -246 232 -240
rect 412 -206 554 -200
rect 412 -240 424 -206
rect 542 -240 554 -206
rect 412 -246 554 -240
rect 734 -206 876 -200
rect 734 -240 746 -206
rect 864 -240 876 -206
rect 734 -246 876 -240
rect 1056 -206 1198 -200
rect 1056 -240 1068 -206
rect 1186 -240 1198 -206
rect 1056 -246 1198 -240
rect 1378 -206 1520 -200
rect 1378 -240 1390 -206
rect 1508 -240 1520 -206
rect 1378 -246 1520 -240
rect 1700 -206 1842 -200
rect 1700 -240 1712 -206
rect 1830 -240 1842 -206
rect 1700 -246 1842 -240
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.95 l 0.75 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
