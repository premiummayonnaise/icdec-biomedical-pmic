magic
tech sky130A
magscale 1 2
timestamp 1769410403
<< nwell >>
rect -3200 -27780 14980 -26000
rect -2840 -27800 14980 -27780
<< pwell >>
rect -3200 -27800 -2840 -27780
rect -3200 -30700 14980 -27800
rect -3200 -30820 3000 -30700
rect 5100 -30820 14920 -30700
rect 14960 -30740 14980 -30700
rect -3200 -30880 12820 -30820
rect 14940 -30880 14980 -30740
rect -3200 -32300 14980 -30880
<< psubdiff >>
rect -3000 -28040 -600 -28000
rect -3000 -28160 -2800 -28040
rect -800 -28160 -600 -28040
rect -3000 -28200 -600 -28160
rect -3000 -30600 -2960 -28200
rect -2840 -30600 -2800 -28200
rect -800 -30600 -760 -28200
rect -640 -30600 -600 -28200
rect -200 -28040 1000 -28000
rect -200 -28160 0 -28040
rect 800 -28160 1000 -28040
rect -200 -28200 1000 -28160
rect -200 -28800 -160 -28200
rect -40 -28800 0 -28200
rect 800 -28800 820 -28200
rect 960 -28800 1000 -28200
rect -200 -28840 1000 -28800
rect -200 -28960 0 -28840
rect 800 -28960 1000 -28840
rect 1400 -28040 3000 -28000
rect 1400 -28160 1600 -28040
rect 2800 -28160 3000 -28040
rect 1400 -28200 3000 -28160
rect 1400 -28800 1440 -28200
rect 1560 -28800 1600 -28200
rect 2800 -28800 2840 -28200
rect 2960 -28800 3000 -28200
rect 1400 -28840 3000 -28800
rect 1400 -28960 1600 -28840
rect 2800 -28960 3000 -28840
rect -204 -29000 1004 -28960
rect 1400 -29000 3000 -28960
rect -204 -29200 1 -29000
rect 799 -29200 1004 -29000
rect 1600 -29200 1802 -29000
rect 2598 -29200 2801 -29000
rect -3000 -30640 -600 -30600
rect -3000 -30760 -2800 -30640
rect -800 -30760 -600 -30640
rect -3000 -30800 -600 -30760
rect -400 -29240 1200 -29200
rect -400 -29360 -200 -29240
rect 1000 -29360 1200 -29240
rect -400 -29400 1200 -29360
rect -400 -30600 -360 -29400
rect -240 -30600 -200 -29400
rect 1000 -30600 1040 -29400
rect 1160 -30600 1200 -29400
rect -400 -30640 1200 -30600
rect -400 -30760 -200 -30640
rect 1000 -30760 1200 -30640
rect -400 -30800 1200 -30760
rect 1600 -29240 2801 -29200
rect 1600 -29360 1800 -29240
rect 2600 -29360 2800 -29240
rect 1600 -29400 2800 -29360
rect 1600 -30600 1640 -29400
rect 1760 -30600 1800 -29400
rect 2600 -30600 2640 -29400
rect 2760 -30600 2800 -29400
rect 1600 -30640 2800 -30600
rect 1600 -30760 1800 -30640
rect 2600 -30760 2800 -30640
rect 1600 -30800 2800 -30760
rect 12820 -29440 14920 -29400
rect 12820 -29560 13020 -29440
rect 14720 -29560 14920 -29440
rect 12820 -29600 14920 -29560
rect 12820 -30600 12860 -29600
rect 12980 -30600 13020 -29600
rect 14720 -30600 14760 -29600
rect 14880 -30600 14920 -29600
rect 12820 -30640 14920 -30600
rect 12820 -30760 13020 -30640
rect 14720 -30760 14920 -30640
rect 12820 -30800 14920 -30760
<< nsubdiff >>
rect -3000 -26240 400 -26200
rect -3000 -26360 -2800 -26240
rect 200 -26360 400 -26240
rect -3000 -26400 400 -26360
rect -3000 -27400 -2960 -26400
rect -2840 -27400 -2800 -26400
rect 200 -27400 240 -26400
rect 360 -27400 400 -26400
rect -3000 -27440 400 -27400
rect -3000 -27560 -2800 -27440
rect 200 -27560 400 -27440
rect -3000 -27600 400 -27560
rect 600 -26240 4000 -26200
rect 600 -26360 800 -26240
rect 3800 -26360 4000 -26240
rect 600 -26400 4000 -26360
rect 600 -27400 640 -26400
rect 760 -27400 800 -26400
rect 3800 -27400 3840 -26400
rect 3960 -27400 4000 -26400
rect 600 -27440 4000 -27400
rect 600 -27560 800 -27440
rect 3800 -27560 4000 -27440
rect 600 -27600 4000 -27560
rect 4200 -26240 14900 -26200
rect 4200 -26360 4400 -26240
rect 14700 -26360 14900 -26240
rect 4200 -26400 14900 -26360
rect 4200 -27500 4240 -26400
rect 4360 -27500 4400 -26400
rect 14700 -27500 14740 -26400
rect 14860 -27500 14900 -26400
rect 4200 -27540 14900 -27500
rect 4200 -27660 4400 -27540
rect 14700 -27660 14900 -27540
rect 4200 -27700 14900 -27660
<< psubdiffcont >>
rect -2800 -28160 -800 -28040
rect -2960 -30600 -2840 -28200
rect -760 -30600 -640 -28200
rect 0 -28160 800 -28040
rect -160 -28800 -40 -28200
rect 820 -28800 960 -28200
rect 0 -28960 800 -28840
rect 1600 -28160 2800 -28040
rect 1440 -28800 1560 -28200
rect 2840 -28800 2960 -28200
rect 1600 -28960 2800 -28840
rect -2800 -30760 -800 -30640
rect -200 -29360 1000 -29240
rect -360 -30600 -240 -29400
rect 1040 -30600 1160 -29400
rect -200 -30760 1000 -30640
rect 1800 -29360 2600 -29240
rect 1640 -30600 1760 -29400
rect 2640 -30600 2760 -29400
rect 1800 -30760 2600 -30640
rect 13020 -29560 14720 -29440
rect 12860 -30600 12980 -29600
rect 14760 -30600 14880 -29600
rect 13020 -30760 14720 -30640
<< nsubdiffcont >>
rect -2800 -26360 200 -26240
rect -2960 -27400 -2840 -26400
rect 240 -27400 360 -26400
rect -2800 -27560 200 -27440
rect 800 -26360 3800 -26240
rect 640 -27400 760 -26400
rect 3840 -27400 3960 -26400
rect 800 -27560 3800 -27440
rect 4400 -26360 14700 -26240
rect 4240 -27500 4360 -26400
rect 14740 -27500 14860 -26400
rect 4400 -27660 14700 -27540
<< locali >>
rect -3200 -24800 14980 -24600
rect -3200 -25400 -3000 -24800
rect -2400 -25400 -2200 -24800
rect -1600 -25400 -1400 -24800
rect -800 -25400 -600 -24800
rect 0 -25400 200 -24800
rect 800 -25400 1000 -24800
rect 1600 -25400 1800 -24800
rect 2400 -25400 2600 -24800
rect 3200 -25400 3400 -24800
rect 4000 -25400 4200 -24800
rect 4800 -25400 5000 -24800
rect 5600 -25400 5800 -24800
rect 6400 -25400 6600 -24800
rect 7200 -25400 7400 -24800
rect 8000 -25400 8200 -24800
rect 8800 -25400 9000 -24800
rect 9600 -25400 9800 -24800
rect 10400 -25400 10600 -24800
rect 11200 -25400 11400 -24800
rect 12000 -25400 12200 -24800
rect 12800 -25400 13000 -24800
rect 13600 -25400 13800 -24800
rect 14400 -25400 14980 -24800
rect -3200 -25600 14980 -25400
rect -3200 -26200 -3000 -25600
rect -2400 -26200 -2200 -25600
rect -1600 -26200 -1400 -25600
rect -800 -26200 -600 -25600
rect 0 -26200 200 -25600
rect 800 -26200 1000 -25600
rect 1600 -26200 1800 -25600
rect 2400 -26200 2600 -25600
rect 3200 -26200 3400 -25600
rect 4000 -26200 4200 -25600
rect 4800 -26200 5000 -25600
rect 5600 -26200 5800 -25600
rect 6400 -26200 6600 -25600
rect 7200 -26200 7400 -25600
rect 8000 -26200 8200 -25600
rect 8800 -26200 9000 -25600
rect 9600 -26200 9800 -25600
rect 10400 -26200 10600 -25600
rect 11200 -26200 11400 -25600
rect 12000 -26200 12200 -25600
rect 12800 -26200 13000 -25600
rect 13600 -26200 13800 -25600
rect 14400 -26200 14980 -25600
rect -3200 -26240 14980 -26200
rect -3200 -26300 -2800 -26240
rect -3000 -26360 -2800 -26300
rect 200 -26300 800 -26240
rect 200 -26360 400 -26300
rect -3000 -26400 400 -26360
rect -3000 -27400 -2960 -26400
rect -2840 -27400 -2800 -26400
rect -2600 -27162 -2499 -26555
rect -2278 -27097 -2179 -26400
rect -1661 -27099 -1562 -26400
rect -1341 -27162 -1262 -26560
rect -1046 -27101 -947 -26400
rect -430 -27097 -331 -26400
rect -124 -27146 -19 -26559
rect -170 -27162 -19 -27146
rect -2600 -27180 -19 -27162
rect -2600 -27240 -100 -27180
rect -40 -27240 -19 -27180
rect -2600 -27259 -19 -27240
rect -2560 -27260 -19 -27259
rect -2560 -27261 -70 -27260
rect 200 -27400 240 -26400
rect 360 -27400 400 -26400
rect -3000 -27440 400 -27400
rect -3000 -27560 -2800 -27440
rect 200 -27560 400 -27440
rect -3000 -27600 400 -27560
rect 600 -26360 800 -26300
rect 3800 -26300 4400 -26240
rect 3800 -26360 4000 -26300
rect 600 -26400 4000 -26360
rect 600 -27400 640 -26400
rect 760 -27400 800 -26400
rect 1321 -27101 1421 -26400
rect 1938 -27105 2038 -26400
rect 2555 -27105 2655 -26400
rect 3170 -27100 3270 -26400
rect 999 -27160 3447 -27146
rect 999 -27201 1020 -27160
rect 997 -27220 1020 -27201
rect 1079 -27220 3447 -27160
rect 997 -27240 3447 -27220
rect 997 -27260 1100 -27240
rect 997 -27320 1020 -27260
rect 1079 -27320 1100 -27260
rect 997 -27340 1100 -27320
rect 3800 -27400 3840 -26400
rect 3960 -27400 4000 -26400
rect 600 -27440 4000 -27400
rect 600 -27560 800 -27440
rect 3800 -27560 4000 -27440
rect 600 -27600 4000 -27560
rect 4200 -26360 4400 -26300
rect 14700 -26300 14980 -26240
rect 14700 -26360 14900 -26300
rect 4200 -26400 14900 -26360
rect 4200 -27500 4240 -26400
rect 4360 -27500 4400 -26400
rect 4919 -27318 5022 -26400
rect 5535 -27319 5638 -26400
rect 6151 -27316 6254 -26400
rect 6769 -27319 6872 -26400
rect 7387 -27319 7490 -26400
rect 8000 -27321 8103 -26400
rect 8618 -27323 8721 -26400
rect 9231 -27319 9334 -26400
rect 9847 -27319 9950 -26400
rect 10466 -27318 10569 -26400
rect 11077 -27318 11180 -26400
rect 11697 -27318 11800 -26400
rect 12311 -27321 12414 -26400
rect 12927 -27321 13030 -26400
rect 13546 -27323 13649 -26400
rect 14162 -27318 14265 -26400
rect 4518 -27360 4673 -27359
rect 4518 -27380 14440 -27360
rect 4518 -27438 4540 -27380
rect 4601 -27438 4639 -27380
rect 4518 -27439 4639 -27438
rect 4700 -27439 14440 -27380
rect 4518 -27460 14440 -27439
rect 4518 -27461 4673 -27460
rect 14700 -27500 14740 -26400
rect 14860 -27500 14900 -26400
rect 4200 -27540 14900 -27500
rect 4200 -27660 4400 -27540
rect 14700 -27660 14900 -27540
rect 4200 -27700 14900 -27660
rect -3000 -28040 -600 -28000
rect -3000 -28160 -2800 -28040
rect -800 -28160 -600 -28040
rect -3000 -28200 -600 -28160
rect -3000 -30600 -2960 -28200
rect -2840 -30600 -2800 -28200
rect -800 -30600 -760 -28200
rect -640 -30600 -600 -28200
rect -200 -28040 1000 -28000
rect -200 -28160 0 -28040
rect 800 -28160 1000 -28040
rect -200 -28200 1000 -28160
rect -200 -28800 -160 -28200
rect -40 -28800 0 -28200
rect 800 -28800 820 -28200
rect 960 -28800 1000 -28200
rect 1400 -28040 3000 -28000
rect 1400 -28160 1600 -28040
rect 2800 -28160 3000 -28040
rect 1400 -28200 3000 -28160
rect 1400 -28800 1440 -28200
rect 1560 -28800 1600 -28200
rect 2800 -28800 2840 -28200
rect 2960 -28800 3000 -28200
rect -204 -28840 1004 -28800
rect -204 -28960 0 -28840
rect 800 -28960 1004 -28840
rect -204 -29000 1004 -28960
rect 1400 -28840 3000 -28800
rect 1400 -28960 1600 -28840
rect 2800 -28960 3000 -28840
rect 1400 -29000 3000 -28960
rect -204 -29200 1 -29000
rect 799 -29200 1004 -29000
rect 1600 -29200 1802 -29000
rect 2598 -29200 2801 -29000
rect -3000 -30640 -600 -30600
rect -3000 -30700 -2800 -30640
rect -3200 -30760 -2800 -30700
rect -800 -30700 -600 -30640
rect -400 -29240 1200 -29200
rect -400 -29360 -200 -29240
rect 1000 -29360 1200 -29240
rect -400 -29400 1200 -29360
rect -400 -30600 -360 -29400
rect -240 -30600 -200 -29400
rect 1000 -30600 1040 -29400
rect 1160 -30600 1200 -29400
rect -400 -30640 1200 -30600
rect -400 -30700 -200 -30640
rect -800 -30760 -200 -30700
rect 1000 -30700 1200 -30640
rect 1600 -29240 2801 -29200
rect 1600 -29360 1800 -29240
rect 2600 -29360 2801 -29240
rect 1600 -29386 2801 -29360
rect 1600 -29400 2800 -29386
rect 1600 -30600 1640 -29400
rect 1760 -30600 1800 -29400
rect 2321 -30600 2420 -29699
rect 2600 -30600 2640 -29400
rect 2760 -30600 2800 -29400
rect 1600 -30640 2800 -30600
rect 1600 -30700 1800 -30640
rect 1000 -30760 1800 -30700
rect 2600 -30700 2800 -30640
rect 12820 -29440 14920 -29400
rect 12820 -29560 13020 -29440
rect 14720 -29560 14920 -29440
rect 12820 -29600 14920 -29560
rect 12820 -30600 12860 -29600
rect 12980 -30600 13020 -29600
rect 13507 -30600 13611 -29872
rect 14121 -30600 14225 -29870
rect 14720 -30600 14760 -29600
rect 14880 -30600 14920 -29600
rect 12820 -30640 14920 -30600
rect 12820 -30700 13020 -30640
rect 2600 -30760 13020 -30700
rect 14720 -30700 14920 -30640
rect 14720 -30760 14980 -30700
rect -3200 -30800 14980 -30760
rect -3200 -31400 -3000 -30800
rect -2400 -31400 -2200 -30800
rect -1600 -31400 -1400 -30800
rect -800 -31400 -600 -30800
rect 0 -31400 200 -30800
rect 800 -31400 1000 -30800
rect 1600 -31400 1800 -30800
rect 2400 -31400 2600 -30800
rect 3200 -31400 3400 -30800
rect 4000 -31400 4200 -30800
rect 4800 -31400 5000 -30800
rect 5600 -31400 5800 -30800
rect 6400 -31400 6600 -30800
rect 7200 -31400 7400 -30800
rect 8000 -31400 8200 -30800
rect 8800 -31400 9000 -30800
rect 9600 -31400 9800 -30800
rect 10400 -31400 10600 -30800
rect 11200 -31400 11400 -30800
rect 12000 -31400 12200 -30800
rect 12800 -31400 13000 -30800
rect 13600 -31400 13800 -30800
rect 14400 -31400 14980 -30800
rect -3200 -31600 14980 -31400
rect -3200 -32200 -3000 -31600
rect -2400 -32200 -2200 -31600
rect -1600 -32200 -1400 -31600
rect -800 -32200 -600 -31600
rect 0 -32200 200 -31600
rect 800 -32200 1000 -31600
rect 1600 -32200 1800 -31600
rect 2400 -32200 2600 -31600
rect 3200 -32200 3400 -31600
rect 4000 -32200 4200 -31600
rect 4800 -32200 5000 -31600
rect 5600 -32200 5800 -31600
rect 6400 -32200 6600 -31600
rect 7200 -32200 7400 -31600
rect 8000 -32200 8200 -31600
rect 8800 -32200 9000 -31600
rect 9600 -32200 9800 -31600
rect 10400 -32200 10600 -31600
rect 11200 -32200 11400 -31600
rect 12000 -32200 12200 -31600
rect 12800 -32200 13000 -31600
rect 13600 -32200 13800 -31600
rect 14400 -32200 14980 -31600
rect -3200 -32400 14980 -32200
<< viali >>
rect -3000 -25400 -2400 -24800
rect -2200 -25400 -1600 -24800
rect -1400 -25400 -800 -24800
rect -600 -25400 0 -24800
rect 200 -25400 800 -24800
rect 1000 -25400 1600 -24800
rect 1800 -25400 2400 -24800
rect 2600 -25400 3200 -24800
rect 3400 -25400 4000 -24800
rect 4200 -25400 4800 -24800
rect 5000 -25400 5600 -24800
rect 5800 -25400 6400 -24800
rect 6600 -25400 7200 -24800
rect 7400 -25400 8000 -24800
rect 8200 -25400 8800 -24800
rect 9000 -25400 9600 -24800
rect 9800 -25400 10400 -24800
rect 10600 -25400 11200 -24800
rect 11400 -25400 12000 -24800
rect 12200 -25400 12800 -24800
rect 13000 -25400 13600 -24800
rect 13800 -25400 14400 -24800
rect -3000 -26200 -2400 -25600
rect -2200 -26200 -1600 -25600
rect -1400 -26200 -800 -25600
rect -600 -26200 0 -25600
rect 200 -26200 800 -25600
rect 1000 -26200 1600 -25600
rect 1800 -26200 2400 -25600
rect 2600 -26200 3200 -25600
rect 3400 -26200 4000 -25600
rect 4200 -26200 4800 -25600
rect 5000 -26200 5600 -25600
rect 5800 -26200 6400 -25600
rect 6600 -26200 7200 -25600
rect 7400 -26200 8000 -25600
rect 8200 -26200 8800 -25600
rect 9000 -26200 9600 -25600
rect 9800 -26200 10400 -25600
rect 10600 -26200 11200 -25600
rect 11400 -26200 12000 -25600
rect 12200 -26200 12800 -25600
rect 13000 -26200 13600 -25600
rect 13800 -26200 14400 -25600
rect -100 -27240 -40 -27180
rect 1020 -27220 1079 -27160
rect 1020 -27320 1079 -27260
rect 4540 -27438 4601 -27380
rect 4639 -27439 4700 -27380
rect -3000 -31400 -2400 -30800
rect -2200 -31400 -1600 -30800
rect -1400 -31400 -800 -30800
rect -600 -31400 0 -30800
rect 200 -31400 800 -30800
rect 1000 -31400 1600 -30800
rect 1800 -31400 2400 -30800
rect 2600 -31400 3200 -30800
rect 3400 -31400 4000 -30800
rect 4200 -31400 4800 -30800
rect 5000 -31400 5600 -30800
rect 5800 -31400 6400 -30800
rect 6600 -31400 7200 -30800
rect 7400 -31400 8000 -30800
rect 8200 -31400 8800 -30800
rect 9000 -31400 9600 -30800
rect 9800 -31400 10400 -30800
rect 10600 -31400 11200 -30800
rect 11400 -31400 12000 -30800
rect 12200 -31400 12800 -30800
rect 13000 -31400 13600 -30800
rect 13800 -31400 14400 -30800
rect -3000 -32200 -2400 -31600
rect -2200 -32200 -1600 -31600
rect -1400 -32200 -800 -31600
rect -600 -32200 0 -31600
rect 200 -32200 800 -31600
rect 1000 -32200 1600 -31600
rect 1800 -32200 2400 -31600
rect 2600 -32200 3200 -31600
rect 3400 -32200 4000 -31600
rect 4200 -32200 4800 -31600
rect 5000 -32200 5600 -31600
rect 5800 -32200 6400 -31600
rect 6600 -32200 7200 -31600
rect 7400 -32200 8000 -31600
rect 8200 -32200 8800 -31600
rect 9000 -32200 9600 -31600
rect 9800 -32200 10400 -31600
rect 10600 -32200 11200 -31600
rect 11400 -32200 12000 -31600
rect 12200 -32200 12800 -31600
rect 13000 -32200 13600 -31600
rect 13800 -32200 14400 -31600
<< metal1 >>
rect -3200 -24800 14980 -24600
rect -3200 -25400 -3000 -24800
rect -2400 -25400 -2200 -24800
rect -1600 -25400 -1400 -24800
rect -800 -25400 -600 -24800
rect 0 -25400 200 -24800
rect 800 -25400 1000 -24800
rect 1600 -25400 1800 -24800
rect 2400 -25400 2600 -24800
rect 3200 -25400 3400 -24800
rect 4000 -25400 4200 -24800
rect 4800 -25400 5000 -24800
rect 5600 -25400 5800 -24800
rect 6400 -25400 6600 -24800
rect 7200 -25400 7400 -24800
rect 8000 -25400 8200 -24800
rect 8800 -25400 9000 -24800
rect 9600 -25400 9800 -24800
rect 10400 -25400 10600 -24800
rect 11200 -25400 11400 -24800
rect 12000 -25400 12200 -24800
rect 12800 -25400 13000 -24800
rect 13600 -25400 13800 -24800
rect 14400 -25400 14980 -24800
rect -3200 -25600 14980 -25400
rect -3200 -26200 -3000 -25600
rect -2400 -26200 -2200 -25600
rect -1600 -26200 -1400 -25600
rect -800 -26200 -600 -25600
rect 0 -26200 200 -25600
rect 800 -26200 1000 -25600
rect 1600 -26200 1800 -25600
rect 2400 -26200 2600 -25600
rect 3200 -26200 3400 -25600
rect 4000 -26200 4200 -25600
rect 4800 -26200 5000 -25600
rect 5600 -26200 5800 -25600
rect 6400 -26200 6600 -25600
rect 7200 -26200 7400 -25600
rect 8000 -26200 8200 -25600
rect 8800 -26200 9000 -25600
rect 9600 -26200 9800 -25600
rect 10400 -26200 10600 -25600
rect 11200 -26200 11400 -25600
rect 12000 -26200 12200 -25600
rect 12800 -26200 13000 -25600
rect 13600 -26200 13800 -25600
rect 14400 -26200 14980 -25600
rect -3200 -26300 14980 -26200
rect -1964 -27492 -1870 -26559
rect -736 -27492 -642 -26559
rect -122 -27180 -16 -26559
rect -122 -27240 -100 -27180
rect -40 -27240 -16 -27180
rect -1965 -27590 -419 -27492
rect -3123 -28455 -2694 -28452
rect -3123 -28737 -2140 -28455
rect -1532 -28608 -1104 -28459
rect -3123 -30700 -2694 -28737
rect -2581 -28959 -2153 -28868
rect -2592 -29430 -2153 -28959
rect -1532 -29079 -1095 -28608
rect -1532 -29152 -1104 -29079
rect -1532 -29330 -1104 -29266
rect -2581 -29561 -2153 -29430
rect -2581 -29752 -2153 -29681
rect -2592 -30223 -2153 -29752
rect -1537 -29801 -1101 -29330
rect -1532 -29959 -1104 -29801
rect -560 -30038 -460 -27590
rect -122 -27922 -16 -27240
rect 996 -27160 1100 -26541
rect 996 -27220 1020 -27160
rect 1079 -27220 1100 -27160
rect 996 -27260 1100 -27220
rect 996 -27320 1020 -27260
rect 1079 -27320 1100 -27260
rect 1630 -27240 1730 -26553
rect 2243 -26621 2351 -26558
rect 2243 -26701 2259 -26621
rect 2339 -26701 2351 -26621
rect 2243 -26719 2351 -26701
rect 2243 -26799 2260 -26719
rect 2340 -26799 2351 -26719
rect 2243 -26820 2351 -26799
rect 2243 -26900 2259 -26820
rect 2339 -26900 2351 -26820
rect 2243 -26920 2351 -26900
rect 2243 -27000 2259 -26920
rect 2339 -27000 2351 -26920
rect 2243 -27020 2351 -27000
rect 2243 -27100 2260 -27020
rect 2340 -27100 2351 -27020
rect 2243 -27120 2351 -27100
rect 2860 -27240 2960 -26555
rect 1630 -27263 2960 -27240
rect 1630 -27273 1924 -27263
rect 1632 -27310 1924 -27273
rect 996 -27400 1100 -27320
rect 1631 -27322 1924 -27310
rect 1984 -27322 2030 -27263
rect 2090 -27310 2960 -27263
rect 2090 -27322 2961 -27310
rect 1631 -27342 2961 -27322
rect 2238 -27394 2354 -27374
rect 2238 -27400 2268 -27394
rect 994 -27421 2268 -27400
rect 994 -27480 1700 -27421
rect 1760 -27480 1819 -27421
rect 1879 -27450 2268 -27421
rect 2322 -27400 2354 -27394
rect 3492 -27400 3596 -26540
rect 4600 -26820 4720 -26760
rect 4600 -26900 4620 -26820
rect 4700 -26900 4720 -26820
rect 4600 -26940 4720 -26900
rect 4600 -27020 4620 -26940
rect 4700 -27020 4720 -26940
rect 4600 -27060 4720 -27020
rect 4600 -27140 4620 -27060
rect 4700 -27140 4720 -27060
rect 4600 -27160 4720 -27140
rect 5220 -26820 5340 -26760
rect 5220 -26900 5240 -26820
rect 5320 -26900 5340 -26820
rect 5220 -26940 5340 -26900
rect 5220 -27020 5240 -26940
rect 5320 -27020 5340 -26940
rect 5220 -27060 5340 -27020
rect 5220 -27140 5240 -27060
rect 5320 -27140 5340 -27060
rect 5220 -27160 5340 -27140
rect 5840 -26820 5960 -26760
rect 5840 -26900 5860 -26820
rect 5940 -26900 5960 -26820
rect 5840 -26940 5960 -26900
rect 5840 -27020 5860 -26940
rect 5940 -27020 5960 -26940
rect 5840 -27060 5960 -27020
rect 5840 -27140 5860 -27060
rect 5940 -27140 5960 -27060
rect 5840 -27160 5960 -27140
rect 6460 -26820 6580 -26760
rect 6460 -26900 6480 -26820
rect 6560 -26900 6580 -26820
rect 6460 -26940 6580 -26900
rect 6460 -27020 6480 -26940
rect 6560 -27020 6580 -26940
rect 6460 -27060 6580 -27020
rect 6460 -27140 6480 -27060
rect 6560 -27140 6580 -27060
rect 6460 -27160 6580 -27140
rect 7060 -26820 7180 -26760
rect 7060 -26900 7080 -26820
rect 7160 -26900 7180 -26820
rect 7060 -26940 7180 -26900
rect 7060 -27020 7080 -26940
rect 7160 -27020 7180 -26940
rect 7060 -27060 7180 -27020
rect 7060 -27140 7080 -27060
rect 7160 -27140 7180 -27060
rect 7060 -27160 7180 -27140
rect 7680 -26820 7800 -26760
rect 7680 -26900 7700 -26820
rect 7780 -26900 7800 -26820
rect 7680 -26940 7800 -26900
rect 7680 -27020 7700 -26940
rect 7780 -27020 7800 -26940
rect 7680 -27060 7800 -27020
rect 7680 -27140 7700 -27060
rect 7780 -27140 7800 -27060
rect 7680 -27160 7800 -27140
rect 8300 -26820 8420 -26760
rect 8300 -26900 8320 -26820
rect 8400 -26900 8420 -26820
rect 8300 -26940 8420 -26900
rect 8300 -27020 8320 -26940
rect 8400 -27020 8420 -26940
rect 8300 -27060 8420 -27020
rect 8300 -27140 8320 -27060
rect 8400 -27140 8420 -27060
rect 8300 -27160 8420 -27140
rect 8920 -26820 9040 -26760
rect 8920 -26900 8940 -26820
rect 9020 -26900 9040 -26820
rect 8920 -26940 9040 -26900
rect 8920 -27020 8940 -26940
rect 9020 -27020 9040 -26940
rect 8920 -27060 9040 -27020
rect 8920 -27140 8940 -27060
rect 9020 -27140 9040 -27060
rect 8920 -27160 9040 -27140
rect 9540 -26820 9660 -26760
rect 9540 -26900 9560 -26820
rect 9640 -26900 9660 -26820
rect 9540 -26940 9660 -26900
rect 9540 -27020 9560 -26940
rect 9640 -27020 9660 -26940
rect 9540 -27060 9660 -27020
rect 9540 -27140 9560 -27060
rect 9640 -27140 9660 -27060
rect 9540 -27160 9660 -27140
rect 10140 -26820 10260 -26760
rect 10140 -26900 10160 -26820
rect 10240 -26900 10260 -26820
rect 10140 -26940 10260 -26900
rect 10140 -27020 10160 -26940
rect 10240 -27020 10260 -26940
rect 10140 -27060 10260 -27020
rect 10140 -27140 10160 -27060
rect 10240 -27140 10260 -27060
rect 10140 -27160 10260 -27140
rect 10760 -26820 10880 -26760
rect 10760 -26900 10780 -26820
rect 10860 -26900 10880 -26820
rect 10760 -26940 10880 -26900
rect 10760 -27020 10780 -26940
rect 10860 -27020 10880 -26940
rect 10760 -27060 10880 -27020
rect 10760 -27140 10780 -27060
rect 10860 -27140 10880 -27060
rect 10760 -27160 10880 -27140
rect 11380 -26820 11500 -26760
rect 11380 -26900 11400 -26820
rect 11480 -26900 11500 -26820
rect 11380 -26940 11500 -26900
rect 11380 -27020 11400 -26940
rect 11480 -27020 11500 -26940
rect 11380 -27060 11500 -27020
rect 11380 -27140 11400 -27060
rect 11480 -27140 11500 -27060
rect 11380 -27160 11500 -27140
rect 12000 -26820 12120 -26760
rect 12000 -26900 12020 -26820
rect 12100 -26900 12120 -26820
rect 12000 -26940 12120 -26900
rect 12000 -27020 12020 -26940
rect 12100 -27020 12120 -26940
rect 12000 -27060 12120 -27020
rect 12000 -27140 12020 -27060
rect 12100 -27140 12120 -27060
rect 12000 -27160 12120 -27140
rect 12600 -26820 12720 -26760
rect 12600 -26900 12620 -26820
rect 12700 -26900 12720 -26820
rect 12600 -26940 12720 -26900
rect 12600 -27020 12620 -26940
rect 12700 -27020 12720 -26940
rect 12600 -27060 12720 -27020
rect 12600 -27140 12620 -27060
rect 12700 -27140 12720 -27060
rect 12600 -27160 12720 -27140
rect 13220 -26820 13340 -26760
rect 13220 -26900 13240 -26820
rect 13320 -26900 13340 -26820
rect 13220 -26940 13340 -26900
rect 13220 -27020 13240 -26940
rect 13320 -27020 13340 -26940
rect 13220 -27060 13340 -27020
rect 13220 -27140 13240 -27060
rect 13320 -27140 13340 -27060
rect 13220 -27160 13340 -27140
rect 13840 -26820 13960 -26760
rect 13840 -26900 13860 -26820
rect 13940 -26900 13960 -26820
rect 13840 -26940 13960 -26900
rect 13840 -27020 13860 -26940
rect 13940 -27020 13960 -26940
rect 13840 -27060 13960 -27020
rect 13840 -27140 13860 -27060
rect 13940 -27140 13960 -27060
rect 13840 -27160 13960 -27140
rect 14460 -26820 14580 -26760
rect 14460 -26900 14480 -26820
rect 14560 -26900 14580 -26820
rect 14460 -26940 14580 -26900
rect 14460 -27020 14480 -26940
rect 14560 -27020 14580 -26940
rect 14460 -27060 14580 -27020
rect 14460 -27140 14480 -27060
rect 14560 -27140 14580 -27060
rect 14460 -27160 14580 -27140
rect 4518 -27360 4673 -27359
rect 4518 -27374 4724 -27360
rect 4518 -27380 4626 -27374
rect 2322 -27422 3597 -27400
rect 2322 -27450 2507 -27422
rect 1879 -27480 2507 -27450
rect 994 -27481 2507 -27480
rect 2567 -27481 2631 -27422
rect 2691 -27481 3597 -27422
rect 4518 -27438 4540 -27380
rect 4601 -27438 4626 -27380
rect 4518 -27461 4626 -27438
rect 4618 -27469 4626 -27461
rect 4712 -27469 4724 -27374
rect 4618 -27481 4724 -27469
rect 994 -27504 3597 -27481
rect 4619 -27517 4723 -27481
rect 2144 -27620 2257 -27596
rect 2144 -27697 2160 -27620
rect 2238 -27697 2257 -27620
rect 2144 -27741 2257 -27697
rect 2144 -27818 2160 -27741
rect 2238 -27818 2257 -27741
rect 4619 -27612 4626 -27517
rect 4712 -27612 4723 -27517
rect 4619 -27654 4723 -27612
rect 4619 -27749 4628 -27654
rect 4714 -27749 4723 -27654
rect 4619 -27761 4723 -27749
rect 2144 -27826 2257 -27818
rect -126 -27964 218 -27922
rect -126 -28024 -98 -27964
rect -38 -28024 0 -27964
rect 60 -28024 112 -27964
rect 172 -28024 218 -27964
rect -126 -28058 218 -28024
rect -122 -28385 -16 -28058
rect 2268 -28141 2447 -28140
rect 1899 -28146 2120 -28141
rect 1899 -28205 1929 -28146
rect 1988 -28205 2048 -28146
rect 2107 -28205 2120 -28146
rect 1899 -28212 2120 -28205
rect 1960 -28213 2120 -28212
rect 2038 -28215 2120 -28213
rect 2268 -28146 2537 -28141
rect 2268 -28205 2368 -28146
rect 2427 -28205 2461 -28146
rect 2520 -28205 2537 -28146
rect 2268 -28213 2537 -28205
rect 2268 -28215 2447 -28213
rect 1836 -28280 2009 -28279
rect 1807 -28287 2009 -28280
rect 1807 -28351 1846 -28287
rect 1908 -28351 1937 -28287
rect 1999 -28351 2009 -28287
rect 1807 -28361 2009 -28351
rect 2040 -28360 2120 -28215
rect 2270 -28360 2350 -28215
rect 2380 -28279 2562 -28278
rect 2380 -28287 2585 -28279
rect 14560 -28280 14880 -28260
rect 2380 -28351 2390 -28287
rect 2452 -28351 2489 -28287
rect 2551 -28351 2585 -28287
rect 2380 -28359 2585 -28351
rect 2400 -28360 2585 -28359
rect 14559 -28360 14580 -28280
rect 14660 -28360 14780 -28280
rect 14860 -28360 14880 -28280
rect -122 -28600 376 -28385
rect 427 -28560 777 -28390
rect 1688 -28448 1796 -28403
rect 1688 -28508 1709 -28448
rect 1769 -28508 1796 -28448
rect 1688 -28520 1796 -28508
rect -122 -28660 460 -28600
rect -122 -28663 376 -28660
rect 617 -29480 725 -28560
rect 1688 -28580 1709 -28520
rect 1769 -28580 1796 -28520
rect 1688 -28594 1796 -28580
rect 1688 -28654 1709 -28594
rect 1769 -28654 1796 -28594
rect 1688 -28668 1796 -28654
rect 1920 -28795 2020 -28404
rect 2150 -28426 2255 -28397
rect 14559 -28400 14880 -28360
rect 2150 -28486 2164 -28426
rect 2224 -28486 2255 -28426
rect 2150 -28502 2255 -28486
rect 2150 -28562 2166 -28502
rect 2226 -28562 2255 -28502
rect 2150 -28578 2255 -28562
rect 2150 -28638 2166 -28578
rect 2226 -28638 2255 -28578
rect 2150 -28652 2255 -28638
rect 1920 -28800 2043 -28795
rect 2379 -28800 2481 -28405
rect 2606 -28445 2712 -28401
rect 2606 -28505 2629 -28445
rect 2689 -28505 2712 -28445
rect 2606 -28518 2712 -28505
rect 2606 -28578 2629 -28518
rect 2689 -28578 2712 -28518
rect 2606 -28592 2712 -28578
rect 2606 -28652 2630 -28592
rect 2690 -28652 2712 -28592
rect 2606 -28664 2712 -28652
rect 14559 -28480 14580 -28400
rect 14660 -28480 14780 -28400
rect 14860 -28401 14880 -28400
rect 15400 -28401 15600 -28400
rect 14860 -28480 15600 -28401
rect 14559 -28520 15600 -28480
rect 14559 -28600 14580 -28520
rect 14660 -28600 14780 -28520
rect 14860 -28600 15600 -28520
rect 14559 -28601 15599 -28600
rect 14559 -28640 14880 -28601
rect 14559 -28720 14580 -28640
rect 14660 -28720 14780 -28640
rect 14860 -28720 14880 -28640
rect 14559 -28733 14880 -28720
rect 1920 -28901 2481 -28800
rect 60 -29528 616 -29527
rect -12 -29633 616 -29528
rect -12 -29640 726 -29633
rect -12 -30038 132 -29640
rect 617 -29641 725 -29640
rect -2581 -30374 -2153 -30223
rect -1538 -30437 -1102 -30083
rect -560 -30138 132 -30038
rect -12 -30384 132 -30138
rect 288 -30437 389 -29694
rect 600 -29760 700 -29700
rect 600 -29820 620 -29760
rect 680 -29820 700 -29760
rect 600 -29840 700 -29820
rect 600 -29900 620 -29840
rect 680 -29900 700 -29840
rect 600 -29920 700 -29900
rect 600 -29980 620 -29920
rect 680 -29980 700 -29920
rect 600 -30000 700 -29980
rect 600 -30060 620 -30000
rect 680 -30060 700 -30000
rect 600 -30080 700 -30060
rect 600 -30140 620 -30080
rect 680 -30140 700 -30080
rect 600 -30160 700 -30140
rect 600 -30220 620 -30160
rect 680 -30220 700 -30160
rect 600 -30240 700 -30220
rect 600 -30300 620 -30240
rect 680 -30300 700 -30240
rect 600 -30320 700 -30300
rect 600 -30380 620 -30320
rect 680 -30380 700 -30320
rect 600 -30400 700 -30380
rect 1941 -30381 2043 -28901
rect 2120 -29600 2280 -29560
rect 2120 -29660 2140 -29600
rect 2200 -29660 2220 -29600
rect 2120 -29680 2280 -29660
rect 13332 -29620 14400 -29563
rect 13332 -29700 13360 -29620
rect 13440 -29700 13460 -29620
rect 13540 -29700 13560 -29620
rect 13640 -29700 13660 -29620
rect 13740 -29700 13760 -29620
rect 13840 -29700 13860 -29620
rect 13940 -29700 13960 -29620
rect 14040 -29700 14060 -29620
rect 14140 -29700 14160 -29620
rect 14240 -29700 14260 -29620
rect 14340 -29700 14400 -29620
rect 13332 -29720 14400 -29700
rect 13332 -29800 13360 -29720
rect 13440 -29800 13460 -29720
rect 13540 -29800 13560 -29720
rect 13640 -29800 13660 -29720
rect 13740 -29800 13760 -29720
rect 13840 -29800 13860 -29720
rect 13940 -29800 13960 -29720
rect 14040 -29800 14060 -29720
rect 14140 -29800 14160 -29720
rect 14240 -29800 14260 -29720
rect 14340 -29800 14400 -29720
rect 13332 -29843 14400 -29800
rect 13180 -29980 13300 -29920
rect 13180 -30060 13200 -29980
rect 13280 -30060 13300 -29980
rect 13180 -30100 13300 -30060
rect 13180 -30180 13200 -30100
rect 13280 -30180 13300 -30100
rect 13180 -30220 13300 -30180
rect 13180 -30300 13200 -30220
rect 13280 -30300 13300 -30220
rect 13180 -30320 13300 -30300
rect 13800 -29980 13920 -29920
rect 13800 -30060 13820 -29980
rect 13900 -30060 13920 -29980
rect 13800 -30100 13920 -30060
rect 13800 -30180 13820 -30100
rect 13900 -30180 13920 -30100
rect 13800 -30220 13920 -30180
rect 13800 -30300 13820 -30220
rect 13900 -30300 13920 -30220
rect 13800 -30320 13920 -30300
rect 14420 -29980 14540 -29920
rect 14420 -30060 14440 -29980
rect 14520 -30060 14540 -29980
rect 14420 -30100 14540 -30060
rect 14420 -30180 14440 -30100
rect 14520 -30180 14540 -30100
rect 14420 -30220 14540 -30180
rect 14420 -30300 14440 -30220
rect 14520 -30300 14540 -30220
rect 14420 -30320 14540 -30300
rect -1538 -30554 422 -30437
rect -1537 -30560 422 -30554
rect -3200 -30800 14980 -30700
rect -3200 -31400 -3000 -30800
rect -2400 -31400 -2200 -30800
rect -1600 -31400 -1400 -30800
rect -800 -31400 -600 -30800
rect 0 -31400 200 -30800
rect 800 -31400 1000 -30800
rect 1600 -31400 1800 -30800
rect 2400 -31400 2600 -30800
rect 3200 -31400 3400 -30800
rect 4000 -31400 4200 -30800
rect 4800 -31400 5000 -30800
rect 5600 -31400 5800 -30800
rect 6400 -31400 6600 -30800
rect 7200 -31400 7400 -30800
rect 8000 -31400 8200 -30800
rect 8800 -31400 9000 -30800
rect 9600 -31400 9800 -30800
rect 10400 -31400 10600 -30800
rect 11200 -31400 11400 -30800
rect 12000 -31400 12200 -30800
rect 12800 -31400 13000 -30800
rect 13600 -31400 13800 -30800
rect 14400 -31400 14980 -30800
rect -3200 -31600 14980 -31400
rect -3200 -32200 -3000 -31600
rect -2400 -32200 -2200 -31600
rect -1600 -32200 -1400 -31600
rect -800 -32200 -600 -31600
rect 0 -32200 200 -31600
rect 800 -32200 1000 -31600
rect 1600 -32200 1800 -31600
rect 2400 -32200 2600 -31600
rect 3200 -32200 3400 -31600
rect 4000 -32200 4200 -31600
rect 4800 -32200 5000 -31600
rect 5600 -32200 5800 -31600
rect 6400 -32200 6600 -31600
rect 7200 -32200 7400 -31600
rect 8000 -32200 8200 -31600
rect 8800 -32200 9000 -31600
rect 9600 -32200 9800 -31600
rect 10400 -32200 10600 -31600
rect 11200 -32200 11400 -31600
rect 12000 -32200 12200 -31600
rect 12800 -32200 13000 -31600
rect 13600 -32200 13800 -31600
rect 14400 -32200 14980 -31600
rect -3200 -32400 14980 -32200
rect 1200 -32620 1400 -32600
rect 1200 -32680 1220 -32620
rect 1280 -32680 1320 -32620
rect 1380 -32680 1400 -32620
rect 1200 -32720 1400 -32680
rect 1200 -32780 1220 -32720
rect 1280 -32780 1320 -32720
rect 1380 -32780 1400 -32720
rect 1200 -32800 1400 -32780
rect 3000 -32620 3200 -32600
rect 3000 -32680 3020 -32620
rect 3080 -32680 3120 -32620
rect 3180 -32680 3200 -32620
rect 3000 -32720 3200 -32680
rect 3000 -32780 3020 -32720
rect 3080 -32780 3120 -32720
rect 3180 -32780 3200 -32720
rect 3000 -32800 3200 -32780
<< rmetal1 >>
rect 616 -29633 726 -29480
<< via1 >>
rect 2259 -26701 2339 -26621
rect 2260 -26799 2340 -26719
rect 2259 -26900 2339 -26820
rect 2259 -27000 2339 -26920
rect 2260 -27100 2340 -27020
rect 1924 -27322 1984 -27263
rect 2030 -27322 2090 -27263
rect 1700 -27480 1760 -27421
rect 1819 -27480 1879 -27421
rect 2268 -27450 2322 -27394
rect 4620 -26900 4700 -26820
rect 4620 -27020 4700 -26940
rect 4620 -27140 4700 -27060
rect 5240 -26900 5320 -26820
rect 5240 -27020 5320 -26940
rect 5240 -27140 5320 -27060
rect 5860 -26900 5940 -26820
rect 5860 -27020 5940 -26940
rect 5860 -27140 5940 -27060
rect 6480 -26900 6560 -26820
rect 6480 -27020 6560 -26940
rect 6480 -27140 6560 -27060
rect 7080 -26900 7160 -26820
rect 7080 -27020 7160 -26940
rect 7080 -27140 7160 -27060
rect 7700 -26900 7780 -26820
rect 7700 -27020 7780 -26940
rect 7700 -27140 7780 -27060
rect 8320 -26900 8400 -26820
rect 8320 -27020 8400 -26940
rect 8320 -27140 8400 -27060
rect 8940 -26900 9020 -26820
rect 8940 -27020 9020 -26940
rect 8940 -27140 9020 -27060
rect 9560 -26900 9640 -26820
rect 9560 -27020 9640 -26940
rect 9560 -27140 9640 -27060
rect 10160 -26900 10240 -26820
rect 10160 -27020 10240 -26940
rect 10160 -27140 10240 -27060
rect 10780 -26900 10860 -26820
rect 10780 -27020 10860 -26940
rect 10780 -27140 10860 -27060
rect 11400 -26900 11480 -26820
rect 11400 -27020 11480 -26940
rect 11400 -27140 11480 -27060
rect 12020 -26900 12100 -26820
rect 12020 -27020 12100 -26940
rect 12020 -27140 12100 -27060
rect 12620 -26900 12700 -26820
rect 12620 -27020 12700 -26940
rect 12620 -27140 12700 -27060
rect 13240 -26900 13320 -26820
rect 13240 -27020 13320 -26940
rect 13240 -27140 13320 -27060
rect 13860 -26900 13940 -26820
rect 13860 -27020 13940 -26940
rect 13860 -27140 13940 -27060
rect 14480 -26900 14560 -26820
rect 14480 -27020 14560 -26940
rect 14480 -27140 14560 -27060
rect 4626 -27380 4712 -27374
rect 2507 -27481 2567 -27422
rect 2631 -27481 2691 -27422
rect 4626 -27439 4639 -27380
rect 4639 -27439 4700 -27380
rect 4700 -27439 4712 -27380
rect 4626 -27469 4712 -27439
rect 2160 -27697 2238 -27620
rect 2160 -27818 2238 -27741
rect 4626 -27612 4712 -27517
rect 4628 -27749 4714 -27654
rect -98 -28024 -38 -27964
rect 0 -28024 60 -27964
rect 112 -28024 172 -27964
rect 1929 -28205 1988 -28146
rect 2048 -28205 2107 -28146
rect 2368 -28205 2427 -28146
rect 2461 -28205 2520 -28146
rect 1846 -28351 1908 -28287
rect 1937 -28351 1999 -28287
rect 2390 -28351 2452 -28287
rect 2489 -28351 2551 -28287
rect 14580 -28360 14660 -28280
rect 14780 -28360 14860 -28280
rect 1709 -28508 1769 -28448
rect 1709 -28580 1769 -28520
rect 1709 -28654 1769 -28594
rect 2164 -28486 2224 -28426
rect 2166 -28562 2226 -28502
rect 2166 -28638 2226 -28578
rect 2629 -28505 2689 -28445
rect 2629 -28578 2689 -28518
rect 2630 -28652 2690 -28592
rect 14580 -28480 14660 -28400
rect 14780 -28480 14860 -28400
rect 14580 -28600 14660 -28520
rect 14780 -28600 14860 -28520
rect 14580 -28720 14660 -28640
rect 14780 -28720 14860 -28640
rect 620 -29820 680 -29760
rect 620 -29900 680 -29840
rect 620 -29980 680 -29920
rect 620 -30060 680 -30000
rect 620 -30140 680 -30080
rect 620 -30220 680 -30160
rect 620 -30300 680 -30240
rect 620 -30380 680 -30320
rect 2140 -29660 2200 -29600
rect 2220 -29660 2280 -29600
rect 13360 -29700 13440 -29620
rect 13460 -29700 13540 -29620
rect 13560 -29700 13640 -29620
rect 13660 -29700 13740 -29620
rect 13760 -29700 13840 -29620
rect 13860 -29700 13940 -29620
rect 13960 -29700 14040 -29620
rect 14060 -29700 14140 -29620
rect 14160 -29700 14240 -29620
rect 14260 -29700 14340 -29620
rect 13360 -29800 13440 -29720
rect 13460 -29800 13540 -29720
rect 13560 -29800 13640 -29720
rect 13660 -29800 13740 -29720
rect 13760 -29800 13840 -29720
rect 13860 -29800 13940 -29720
rect 13960 -29800 14040 -29720
rect 14060 -29800 14140 -29720
rect 14160 -29800 14240 -29720
rect 14260 -29800 14340 -29720
rect 13200 -30060 13280 -29980
rect 13200 -30180 13280 -30100
rect 13200 -30300 13280 -30220
rect 13820 -30060 13900 -29980
rect 13820 -30180 13900 -30100
rect 13820 -30300 13900 -30220
rect 14440 -30060 14520 -29980
rect 14440 -30180 14520 -30100
rect 14440 -30300 14520 -30220
rect 1220 -32680 1280 -32620
rect 1320 -32680 1380 -32620
rect 1220 -32780 1280 -32720
rect 1320 -32780 1380 -32720
rect 3020 -32680 3080 -32620
rect 3120 -32680 3180 -32620
rect 3020 -32780 3080 -32720
rect 3120 -32780 3180 -32720
<< metal2 >>
rect 2245 -26621 2351 -26559
rect 2245 -26701 2259 -26621
rect 2339 -26701 2351 -26621
rect 2245 -26719 2351 -26701
rect 2245 -26799 2260 -26719
rect 2340 -26799 2351 -26719
rect 2245 -26820 2351 -26799
rect 2245 -26900 2259 -26820
rect 2339 -26900 2351 -26820
rect 2245 -26920 2351 -26900
rect 2245 -27000 2259 -26920
rect 2339 -27000 2351 -26920
rect 2245 -27020 2351 -27000
rect 2245 -27100 2260 -27020
rect 2340 -27100 2351 -27020
rect 2245 -27102 2351 -27100
rect 4600 -26820 4720 -26760
rect 4600 -26900 4620 -26820
rect 4700 -26900 4720 -26820
rect 4600 -26940 4720 -26900
rect 4600 -27020 4620 -26940
rect 4700 -27020 4720 -26940
rect 4600 -27060 4720 -27020
rect 1894 -27263 2124 -27240
rect 1894 -27322 1924 -27263
rect 1984 -27322 2030 -27263
rect 2090 -27322 2124 -27263
rect 1894 -27342 2124 -27322
rect 1688 -27400 1804 -27399
rect 1688 -27420 1900 -27400
rect 1688 -27482 1700 -27420
rect 1762 -27482 1818 -27420
rect 1880 -27482 1900 -27420
rect 1688 -27502 1900 -27482
rect 1689 -27504 1900 -27502
rect 2010 -27502 2124 -27342
rect 2240 -27374 2354 -27102
rect 4600 -27140 4620 -27060
rect 4700 -27140 4720 -27060
rect 4600 -27160 4720 -27140
rect 5220 -26820 5340 -26760
rect 5220 -26900 5240 -26820
rect 5320 -26900 5340 -26820
rect 5220 -26940 5340 -26900
rect 5220 -27020 5240 -26940
rect 5320 -27020 5340 -26940
rect 5220 -27060 5340 -27020
rect 5220 -27140 5240 -27060
rect 5320 -27140 5340 -27060
rect 5220 -27160 5340 -27140
rect 5840 -26820 5960 -26760
rect 5840 -26900 5860 -26820
rect 5940 -26900 5960 -26820
rect 5840 -26940 5960 -26900
rect 5840 -27020 5860 -26940
rect 5940 -27020 5960 -26940
rect 5840 -27060 5960 -27020
rect 5840 -27140 5860 -27060
rect 5940 -27140 5960 -27060
rect 5840 -27160 5960 -27140
rect 6460 -26820 6580 -26760
rect 6460 -26900 6480 -26820
rect 6560 -26900 6580 -26820
rect 6460 -26940 6580 -26900
rect 6460 -27020 6480 -26940
rect 6560 -27020 6580 -26940
rect 6460 -27060 6580 -27020
rect 6460 -27140 6480 -27060
rect 6560 -27140 6580 -27060
rect 6460 -27160 6580 -27140
rect 7060 -26820 7180 -26760
rect 7060 -26900 7080 -26820
rect 7160 -26900 7180 -26820
rect 7060 -26940 7180 -26900
rect 7060 -27020 7080 -26940
rect 7160 -27020 7180 -26940
rect 7060 -27060 7180 -27020
rect 7060 -27140 7080 -27060
rect 7160 -27140 7180 -27060
rect 7060 -27160 7180 -27140
rect 7680 -26820 7800 -26760
rect 7680 -26900 7700 -26820
rect 7780 -26900 7800 -26820
rect 7680 -26940 7800 -26900
rect 7680 -27020 7700 -26940
rect 7780 -27020 7800 -26940
rect 7680 -27060 7800 -27020
rect 7680 -27140 7700 -27060
rect 7780 -27140 7800 -27060
rect 7680 -27160 7800 -27140
rect 8300 -26820 8420 -26760
rect 8300 -26900 8320 -26820
rect 8400 -26900 8420 -26820
rect 8300 -26940 8420 -26900
rect 8300 -27020 8320 -26940
rect 8400 -27020 8420 -26940
rect 8300 -27060 8420 -27020
rect 8300 -27140 8320 -27060
rect 8400 -27140 8420 -27060
rect 8300 -27160 8420 -27140
rect 8920 -26820 9040 -26760
rect 8920 -26900 8940 -26820
rect 9020 -26900 9040 -26820
rect 8920 -26940 9040 -26900
rect 8920 -27020 8940 -26940
rect 9020 -27020 9040 -26940
rect 8920 -27060 9040 -27020
rect 8920 -27140 8940 -27060
rect 9020 -27140 9040 -27060
rect 8920 -27160 9040 -27140
rect 9540 -26820 9660 -26760
rect 9540 -26900 9560 -26820
rect 9640 -26900 9660 -26820
rect 9540 -26940 9660 -26900
rect 9540 -27020 9560 -26940
rect 9640 -27020 9660 -26940
rect 9540 -27060 9660 -27020
rect 9540 -27140 9560 -27060
rect 9640 -27140 9660 -27060
rect 9540 -27160 9660 -27140
rect 10140 -26820 10260 -26760
rect 10140 -26900 10160 -26820
rect 10240 -26900 10260 -26820
rect 10140 -26940 10260 -26900
rect 10140 -27020 10160 -26940
rect 10240 -27020 10260 -26940
rect 10140 -27060 10260 -27020
rect 10140 -27140 10160 -27060
rect 10240 -27140 10260 -27060
rect 10140 -27160 10260 -27140
rect 10760 -26820 10880 -26760
rect 10760 -26900 10780 -26820
rect 10860 -26900 10880 -26820
rect 10760 -26940 10880 -26900
rect 10760 -27020 10780 -26940
rect 10860 -27020 10880 -26940
rect 10760 -27060 10880 -27020
rect 10760 -27140 10780 -27060
rect 10860 -27140 10880 -27060
rect 10760 -27160 10880 -27140
rect 11380 -26820 11500 -26760
rect 11380 -26900 11400 -26820
rect 11480 -26900 11500 -26820
rect 11380 -26940 11500 -26900
rect 11380 -27020 11400 -26940
rect 11480 -27020 11500 -26940
rect 11380 -27060 11500 -27020
rect 11380 -27140 11400 -27060
rect 11480 -27140 11500 -27060
rect 11380 -27160 11500 -27140
rect 12000 -26820 12120 -26760
rect 12000 -26900 12020 -26820
rect 12100 -26900 12120 -26820
rect 12000 -26940 12120 -26900
rect 12000 -27020 12020 -26940
rect 12100 -27020 12120 -26940
rect 12000 -27060 12120 -27020
rect 12000 -27140 12020 -27060
rect 12100 -27140 12120 -27060
rect 12000 -27160 12120 -27140
rect 12600 -26820 12720 -26760
rect 12600 -26900 12620 -26820
rect 12700 -26900 12720 -26820
rect 12600 -26940 12720 -26900
rect 12600 -27020 12620 -26940
rect 12700 -27020 12720 -26940
rect 12600 -27060 12720 -27020
rect 12600 -27140 12620 -27060
rect 12700 -27140 12720 -27060
rect 12600 -27160 12720 -27140
rect 13220 -26820 13340 -26760
rect 13220 -26900 13240 -26820
rect 13320 -26900 13340 -26820
rect 13220 -26940 13340 -26900
rect 13220 -27020 13240 -26940
rect 13320 -27020 13340 -26940
rect 13220 -27060 13340 -27020
rect 13220 -27140 13240 -27060
rect 13320 -27140 13340 -27060
rect 13220 -27160 13340 -27140
rect 13840 -26820 13960 -26760
rect 13840 -26900 13860 -26820
rect 13940 -26900 13960 -26820
rect 13840 -26940 13960 -26900
rect 13840 -27020 13860 -26940
rect 13940 -27020 13960 -26940
rect 13840 -27060 13960 -27020
rect 13840 -27140 13860 -27060
rect 13940 -27140 13960 -27060
rect 13840 -27160 13960 -27140
rect 14460 -26820 14580 -26760
rect 14460 -26900 14480 -26820
rect 14560 -26900 14580 -26820
rect 14460 -26940 14580 -26900
rect 14460 -27020 14480 -26940
rect 14560 -27020 14580 -26940
rect 14460 -27060 14580 -27020
rect 14460 -27140 14480 -27060
rect 14560 -27140 14580 -27060
rect 14460 -27160 14580 -27140
rect 2238 -27394 2354 -27374
rect 2238 -27446 2268 -27394
rect 2240 -27450 2268 -27446
rect 2322 -27398 2354 -27394
rect 4619 -27374 4723 -27360
rect 2322 -27400 2580 -27398
rect 2322 -27420 2710 -27400
rect 2322 -27422 2630 -27420
rect 2692 -27422 2710 -27420
rect 2322 -27424 2506 -27422
rect 2322 -27450 2366 -27424
rect 2240 -27460 2366 -27450
rect 2300 -27486 2366 -27460
rect 2428 -27484 2506 -27424
rect 2568 -27482 2630 -27422
rect 2692 -27482 2712 -27422
rect 2568 -27484 2712 -27482
rect 2428 -27486 2712 -27484
rect 2300 -27500 2712 -27486
rect -126 -27964 1072 -27926
rect -126 -28024 -98 -27964
rect -38 -28024 0 -27964
rect 60 -28024 112 -27964
rect 172 -28024 1072 -27964
rect -126 -28058 1072 -28024
rect 940 -29560 1072 -28058
rect 1690 -28448 1796 -27504
rect 2010 -27596 2256 -27502
rect 2488 -27504 2712 -27500
rect 2010 -27598 2257 -27596
rect 2144 -27620 2257 -27598
rect 2144 -27697 2160 -27620
rect 2238 -27697 2257 -27620
rect 2144 -27740 2257 -27697
rect 2144 -27818 2160 -27740
rect 2239 -27792 2257 -27740
rect 2239 -27817 2259 -27792
rect 2238 -27818 2259 -27817
rect 2144 -27822 2259 -27818
rect 2144 -27826 2257 -27822
rect 2145 -27828 2256 -27826
rect 2146 -28081 2253 -27828
rect 2146 -28127 2256 -28081
rect 1899 -28146 2120 -28141
rect 1899 -28205 1929 -28146
rect 1988 -28205 2048 -28146
rect 2107 -28205 2120 -28146
rect 1899 -28212 2120 -28205
rect 1900 -28213 2120 -28212
rect 2038 -28215 2120 -28213
rect 1836 -28287 2009 -28279
rect 1836 -28351 1846 -28287
rect 1908 -28351 1937 -28287
rect 1999 -28351 2009 -28287
rect 1836 -28361 2009 -28351
rect 1690 -28508 1709 -28448
rect 1769 -28508 1796 -28448
rect 1690 -28520 1796 -28508
rect 1690 -28580 1709 -28520
rect 1769 -28580 1796 -28520
rect 1690 -28594 1796 -28580
rect 1690 -28654 1709 -28594
rect 1769 -28654 1796 -28594
rect 2150 -28426 2256 -28127
rect 2349 -28141 2446 -28140
rect 2349 -28146 2537 -28141
rect 2349 -28205 2368 -28146
rect 2427 -28205 2461 -28146
rect 2520 -28205 2537 -28146
rect 2349 -28213 2537 -28205
rect 2380 -28287 2562 -28278
rect 2380 -28351 2390 -28287
rect 2452 -28351 2489 -28287
rect 2551 -28351 2562 -28287
rect 2380 -28359 2562 -28351
rect 2400 -28360 2562 -28359
rect 2150 -28486 2164 -28426
rect 2224 -28486 2256 -28426
rect 2150 -28502 2256 -28486
rect 2150 -28562 2166 -28502
rect 2226 -28562 2256 -28502
rect 2150 -28578 2256 -28562
rect 2150 -28638 2166 -28578
rect 2226 -28638 2256 -28578
rect 2150 -28651 2256 -28638
rect 2606 -28445 2712 -27504
rect 4619 -27469 4626 -27374
rect 4712 -27469 4723 -27374
rect 4619 -27517 4723 -27469
rect 4619 -27612 4626 -27517
rect 4713 -27612 4723 -27517
rect 4619 -27654 4723 -27612
rect 4619 -27749 4628 -27654
rect 4714 -27749 4723 -27654
rect 4619 -27761 4723 -27749
rect 14560 -28280 14880 -28260
rect 2606 -28505 2629 -28445
rect 2689 -28505 2712 -28445
rect 2606 -28518 2712 -28505
rect 2606 -28578 2629 -28518
rect 2689 -28578 2712 -28518
rect 2606 -28592 2712 -28578
rect 1690 -28666 1796 -28654
rect 2606 -28652 2630 -28592
rect 2690 -28652 2712 -28592
rect 2606 -28663 2712 -28652
rect 14559 -28360 14580 -28280
rect 14660 -28360 14780 -28280
rect 14860 -28360 14880 -28280
rect 14559 -28400 14880 -28360
rect 14559 -28480 14580 -28400
rect 14660 -28480 14780 -28400
rect 14860 -28401 14880 -28400
rect 14860 -28480 15599 -28401
rect 14559 -28520 15599 -28480
rect 14559 -28600 14580 -28520
rect 14660 -28600 14780 -28520
rect 14860 -28600 15599 -28520
rect 14559 -28601 15599 -28600
rect 14559 -28640 14880 -28601
rect 14559 -28720 14580 -28640
rect 14660 -28720 14780 -28640
rect 14860 -28720 14880 -28640
rect 14559 -28733 14880 -28720
rect 591 -29600 14480 -29560
rect 591 -29660 2140 -29600
rect 2200 -29660 2220 -29600
rect 2280 -29620 14480 -29600
rect 2280 -29660 13360 -29620
rect 591 -29678 13360 -29660
rect 591 -29760 723 -29678
rect 591 -29820 620 -29760
rect 680 -29820 723 -29760
rect 591 -29840 723 -29820
rect 13340 -29700 13360 -29678
rect 13440 -29700 13460 -29620
rect 13540 -29700 13560 -29620
rect 13640 -29700 13660 -29620
rect 13740 -29700 13760 -29620
rect 13840 -29700 13860 -29620
rect 13940 -29700 13960 -29620
rect 14040 -29700 14060 -29620
rect 14140 -29700 14160 -29620
rect 14240 -29700 14260 -29620
rect 14340 -29678 14480 -29620
rect 14340 -29700 14400 -29678
rect 13340 -29720 14400 -29700
rect 13340 -29800 13360 -29720
rect 13440 -29800 13460 -29720
rect 13540 -29800 13560 -29720
rect 13640 -29800 13660 -29720
rect 13740 -29800 13760 -29720
rect 13840 -29800 13860 -29720
rect 13940 -29800 13960 -29720
rect 14040 -29800 14060 -29720
rect 14140 -29800 14160 -29720
rect 14240 -29800 14260 -29720
rect 14340 -29800 14400 -29720
rect 13340 -29840 14400 -29800
rect 591 -29900 620 -29840
rect 680 -29900 723 -29840
rect 591 -29920 723 -29900
rect 591 -29980 620 -29920
rect 680 -29980 723 -29920
rect 591 -30000 723 -29980
rect 591 -30012 620 -30000
rect 680 -30060 723 -30000
rect 620 -30080 723 -30060
rect 591 -30140 620 -30117
rect 680 -30140 723 -30080
rect 591 -30160 723 -30140
rect 591 -30220 620 -30160
rect 680 -30220 723 -30160
rect 591 -30240 723 -30220
rect 591 -30300 620 -30240
rect 680 -30300 723 -30240
rect 591 -30320 723 -30300
rect 13180 -29980 13300 -29920
rect 13180 -30060 13200 -29980
rect 13280 -30060 13300 -29980
rect 13180 -30100 13300 -30060
rect 13180 -30180 13200 -30100
rect 13280 -30180 13300 -30100
rect 13180 -30220 13300 -30180
rect 13180 -30300 13200 -30220
rect 13280 -30300 13300 -30220
rect 13180 -30320 13300 -30300
rect 13800 -29980 13920 -29920
rect 13800 -30060 13820 -29980
rect 13900 -30060 13920 -29980
rect 13800 -30100 13920 -30060
rect 13800 -30180 13820 -30100
rect 13900 -30180 13920 -30100
rect 13800 -30220 13920 -30180
rect 13800 -30300 13820 -30220
rect 13900 -30300 13920 -30220
rect 13800 -30320 13920 -30300
rect 14420 -29980 14540 -29920
rect 14420 -30060 14440 -29980
rect 14520 -30060 14540 -29980
rect 14420 -30100 14540 -30060
rect 14420 -30180 14440 -30100
rect 14520 -30180 14540 -30100
rect 14420 -30220 14540 -30180
rect 14420 -30300 14440 -30220
rect 14520 -30300 14540 -30220
rect 14420 -30320 14540 -30300
rect 591 -30380 620 -30320
rect 680 -30380 723 -30320
rect 591 -30400 723 -30380
rect 1200 -32620 1400 -32600
rect 1200 -32680 1220 -32620
rect 1280 -32680 1320 -32620
rect 1380 -32680 1400 -32620
rect 1200 -32720 1400 -32680
rect 1200 -32780 1220 -32720
rect 1280 -32780 1320 -32720
rect 1380 -32780 1400 -32720
rect 1200 -32800 1400 -32780
rect 3000 -32620 3200 -32600
rect 3000 -32680 3020 -32620
rect 3080 -32680 3120 -32620
rect 3180 -32680 3200 -32620
rect 3000 -32720 3200 -32680
rect 3000 -32780 3020 -32720
rect 3080 -32780 3120 -32720
rect 3180 -32780 3200 -32720
rect 3000 -32800 3200 -32780
<< via2 >>
rect 4620 -26900 4700 -26820
rect 4620 -27020 4700 -26940
rect 1700 -27421 1762 -27420
rect 1700 -27480 1760 -27421
rect 1760 -27480 1762 -27421
rect 1700 -27482 1762 -27480
rect 1818 -27421 1880 -27420
rect 1818 -27480 1819 -27421
rect 1819 -27480 1879 -27421
rect 1879 -27480 1880 -27421
rect 1818 -27482 1880 -27480
rect 4620 -27140 4700 -27060
rect 5240 -26900 5320 -26820
rect 5240 -27020 5320 -26940
rect 5240 -27140 5320 -27060
rect 5860 -26900 5940 -26820
rect 5860 -27020 5940 -26940
rect 5860 -27140 5940 -27060
rect 6480 -26900 6560 -26820
rect 6480 -27020 6560 -26940
rect 6480 -27140 6560 -27060
rect 7080 -26900 7160 -26820
rect 7080 -27020 7160 -26940
rect 7080 -27140 7160 -27060
rect 7700 -26900 7780 -26820
rect 7700 -27020 7780 -26940
rect 7700 -27140 7780 -27060
rect 8320 -26900 8400 -26820
rect 8320 -27020 8400 -26940
rect 8320 -27140 8400 -27060
rect 8940 -26900 9020 -26820
rect 8940 -27020 9020 -26940
rect 8940 -27140 9020 -27060
rect 9560 -26900 9640 -26820
rect 9560 -27020 9640 -26940
rect 9560 -27140 9640 -27060
rect 10160 -26900 10240 -26820
rect 10160 -27020 10240 -26940
rect 10160 -27140 10240 -27060
rect 10780 -26900 10860 -26820
rect 10780 -27020 10860 -26940
rect 10780 -27140 10860 -27060
rect 11400 -26900 11480 -26820
rect 11400 -27020 11480 -26940
rect 11400 -27140 11480 -27060
rect 12020 -26900 12100 -26820
rect 12020 -27020 12100 -26940
rect 12020 -27140 12100 -27060
rect 12620 -26900 12700 -26820
rect 12620 -27020 12700 -26940
rect 12620 -27140 12700 -27060
rect 13240 -26900 13320 -26820
rect 13240 -27020 13320 -26940
rect 13240 -27140 13320 -27060
rect 13860 -26900 13940 -26820
rect 13860 -27020 13940 -26940
rect 13860 -27140 13940 -27060
rect 14480 -26900 14560 -26820
rect 14480 -27020 14560 -26940
rect 14480 -27140 14560 -27060
rect 2630 -27422 2692 -27420
rect 2366 -27486 2428 -27424
rect 2506 -27481 2507 -27422
rect 2507 -27481 2567 -27422
rect 2567 -27481 2568 -27422
rect 2506 -27484 2568 -27481
rect 2630 -27481 2631 -27422
rect 2631 -27481 2691 -27422
rect 2691 -27481 2692 -27422
rect 2630 -27482 2692 -27481
rect 2160 -27697 2238 -27620
rect 2160 -27741 2239 -27740
rect 2160 -27818 2238 -27741
rect 2238 -27817 2239 -27741
rect 1929 -28205 1988 -28146
rect 2048 -28205 2107 -28146
rect 1846 -28351 1908 -28287
rect 1937 -28351 1999 -28287
rect 2368 -28205 2427 -28146
rect 2461 -28205 2520 -28146
rect 2390 -28351 2452 -28287
rect 2489 -28351 2551 -28287
rect 4626 -27469 4712 -27374
rect 4626 -27612 4712 -27517
rect 4712 -27612 4713 -27517
rect 4628 -27749 4714 -27654
rect 14580 -28360 14660 -28280
rect 14780 -28360 14860 -28280
rect 14580 -28480 14660 -28400
rect 14780 -28480 14860 -28400
rect 14580 -28600 14660 -28520
rect 14780 -28600 14860 -28520
rect 14580 -28720 14660 -28640
rect 14780 -28720 14860 -28640
rect 13200 -30060 13280 -29980
rect 13200 -30180 13280 -30100
rect 13200 -30300 13280 -30220
rect 13820 -30060 13900 -29980
rect 13820 -30180 13900 -30100
rect 13820 -30300 13900 -30220
rect 14440 -30060 14520 -29980
rect 14440 -30180 14520 -30100
rect 14440 -30300 14520 -30220
rect 1220 -32680 1280 -32620
rect 1320 -32680 1380 -32620
rect 1220 -32780 1280 -32720
rect 1320 -32780 1380 -32720
rect 3020 -32680 3080 -32620
rect 3120 -32680 3180 -32620
rect 3020 -32780 3080 -32720
rect 3120 -32780 3180 -32720
<< metal3 >>
rect 14560 -26760 14880 -26360
rect 4200 -26820 14880 -26760
rect 4200 -26900 4620 -26820
rect 4700 -26900 5240 -26820
rect 5320 -26900 5860 -26820
rect 5940 -26900 6480 -26820
rect 6560 -26900 7080 -26820
rect 7160 -26900 7700 -26820
rect 7780 -26900 8320 -26820
rect 8400 -26900 8940 -26820
rect 9020 -26900 9560 -26820
rect 9640 -26900 10160 -26820
rect 10240 -26900 10780 -26820
rect 10860 -26900 11400 -26820
rect 11480 -26900 12020 -26820
rect 12100 -26900 12620 -26820
rect 12700 -26900 13240 -26820
rect 13320 -26900 13860 -26820
rect 13940 -26900 14480 -26820
rect 14560 -26900 14880 -26820
rect 4200 -26940 14880 -26900
rect 4200 -27020 4620 -26940
rect 4700 -27020 5240 -26940
rect 5320 -27020 5860 -26940
rect 5940 -27020 6480 -26940
rect 6560 -27020 7080 -26940
rect 7160 -27020 7700 -26940
rect 7780 -27020 8320 -26940
rect 8400 -27020 8940 -26940
rect 9020 -27020 9560 -26940
rect 9640 -27020 10160 -26940
rect 10240 -27020 10780 -26940
rect 10860 -27020 11400 -26940
rect 11480 -27020 12020 -26940
rect 12100 -27020 12620 -26940
rect 12700 -27020 13240 -26940
rect 13320 -27020 13860 -26940
rect 13940 -27020 14480 -26940
rect 14560 -27020 14880 -26940
rect 4200 -27060 14880 -27020
rect 4200 -27140 4620 -27060
rect 4700 -27140 5240 -27060
rect 5320 -27140 5860 -27060
rect 5940 -27140 6480 -27060
rect 6560 -27140 7080 -27060
rect 7160 -27140 7700 -27060
rect 7780 -27140 8320 -27060
rect 8400 -27140 8940 -27060
rect 9020 -27140 9560 -27060
rect 9640 -27140 10160 -27060
rect 10240 -27140 10780 -27060
rect 10860 -27140 11400 -27060
rect 11480 -27140 12020 -27060
rect 12100 -27140 12620 -27060
rect 12700 -27140 13240 -27060
rect 13320 -27140 13860 -27060
rect 13940 -27140 14480 -27060
rect 14560 -27140 14880 -27060
rect 4200 -27160 14880 -27140
rect 4619 -27374 4723 -27360
rect 1690 -27420 2710 -27402
rect 1690 -27482 1700 -27420
rect 1762 -27482 1818 -27420
rect 1880 -27422 2630 -27420
rect 1880 -27424 2506 -27422
rect 1880 -27482 2366 -27424
rect 1690 -27486 2366 -27482
rect 2428 -27484 2506 -27424
rect 2568 -27482 2630 -27422
rect 2692 -27482 2710 -27420
rect 2568 -27484 2710 -27482
rect 2428 -27486 2710 -27484
rect 1690 -27500 2710 -27486
rect 4619 -27469 4626 -27374
rect 4713 -27469 4723 -27374
rect 4619 -27517 4723 -27469
rect 2144 -27620 2257 -27596
rect 2144 -27697 2160 -27620
rect 2238 -27697 2257 -27620
rect 2144 -27740 2257 -27697
rect 2144 -27818 2160 -27740
rect 2239 -27817 2257 -27740
rect 4619 -27612 4626 -27517
rect 4713 -27612 4723 -27517
rect 4619 -27654 4723 -27612
rect 4619 -27749 4628 -27654
rect 4714 -27749 4723 -27654
rect 4619 -27761 4723 -27749
rect 2238 -27818 2257 -27817
rect 2144 -27826 2257 -27818
rect 1808 -28146 3199 -28139
rect 1200 -28280 1400 -28200
rect 1808 -28205 1929 -28146
rect 1988 -28205 2048 -28146
rect 2107 -28205 2368 -28146
rect 2427 -28205 2461 -28146
rect 2520 -28200 3199 -28146
rect 2520 -28205 3200 -28200
rect 1808 -28218 3200 -28205
rect 1200 -28287 2580 -28280
rect 1200 -28351 1846 -28287
rect 1908 -28351 1937 -28287
rect 1999 -28351 2390 -28287
rect 2452 -28351 2489 -28287
rect 2551 -28351 2580 -28287
rect 1200 -28360 2580 -28351
rect 1200 -32620 1400 -28360
rect 1200 -32680 1220 -32620
rect 1280 -32680 1320 -32620
rect 1380 -32680 1400 -32620
rect 1200 -32720 1400 -32680
rect 1200 -32780 1220 -32720
rect 1280 -32780 1320 -32720
rect 1380 -32780 1400 -32720
rect 1200 -32800 1400 -32780
rect 3000 -32620 3200 -28218
rect 14560 -28280 14880 -27160
rect 14560 -28360 14580 -28280
rect 14660 -28360 14780 -28280
rect 14860 -28360 14880 -28280
rect 14560 -28400 14880 -28360
rect 14560 -28480 14580 -28400
rect 14660 -28480 14780 -28400
rect 14860 -28480 14880 -28400
rect 14560 -28520 14880 -28480
rect 14560 -28600 14580 -28520
rect 14660 -28600 14780 -28520
rect 14860 -28600 14880 -28520
rect 14560 -28640 14880 -28600
rect 14560 -28720 14580 -28640
rect 14660 -28720 14780 -28640
rect 14860 -28720 14880 -28640
rect 14560 -29920 14880 -28720
rect 3000 -32680 3020 -32620
rect 3080 -32680 3120 -32620
rect 3180 -32680 3200 -32620
rect 3000 -32720 3200 -32680
rect 3000 -32780 3020 -32720
rect 3080 -32780 3120 -32720
rect 3180 -32780 3200 -32720
rect 3000 -32800 3200 -32780
rect 12500 -29980 14880 -29920
rect 12500 -30000 13200 -29980
rect 12500 -30080 12520 -30000
rect 12600 -30080 12640 -30000
rect 12720 -30080 12760 -30000
rect 12840 -30060 13200 -30000
rect 13280 -30060 13820 -29980
rect 13900 -30060 14440 -29980
rect 14520 -30060 14880 -29980
rect 12840 -30080 14880 -30060
rect 12500 -30100 14880 -30080
rect 12500 -30120 13200 -30100
rect 12500 -30200 12520 -30120
rect 12600 -30200 12640 -30120
rect 12720 -30200 12760 -30120
rect 12840 -30180 13200 -30120
rect 13280 -30180 13820 -30100
rect 13900 -30180 14440 -30100
rect 14520 -30180 14880 -30100
rect 12840 -30200 14880 -30180
rect 12500 -30220 14880 -30200
rect 12500 -30240 13200 -30220
rect 12500 -30320 12520 -30240
rect 12600 -30320 12640 -30240
rect 12720 -30320 12760 -30240
rect 12840 -30300 13200 -30240
rect 13280 -30300 13820 -30220
rect 13900 -30300 14440 -30220
rect 14520 -30300 14880 -30220
rect 12840 -30320 14880 -30300
rect 12500 -30360 12860 -30320
rect 12500 -30440 12520 -30360
rect 12600 -30440 12640 -30360
rect 12720 -30440 12760 -30360
rect 12840 -30440 12860 -30360
rect 12500 -34620 12860 -30440
rect 12500 -34700 12520 -34620
rect 12600 -34700 12640 -34620
rect 12720 -34700 12760 -34620
rect 12840 -34700 12860 -34620
rect 12500 -34720 12860 -34700
rect 12500 -34800 12520 -34720
rect 12600 -34800 12640 -34720
rect 12720 -34800 12760 -34720
rect 12840 -34800 12860 -34720
rect 12500 -34820 12860 -34800
rect 12500 -34900 12520 -34820
rect 12600 -34900 12640 -34820
rect 12720 -34900 12760 -34820
rect 12840 -34900 12860 -34820
rect 12500 -34920 12860 -34900
rect 12500 -35000 12520 -34920
rect 12600 -35000 12640 -34920
rect 12720 -35000 12760 -34920
rect 12840 -35000 12860 -34920
rect 12500 -35020 12860 -35000
<< via3 >>
rect 4626 -27469 4712 -27374
rect 4712 -27469 4713 -27374
rect 2160 -27697 2238 -27620
rect 2160 -27818 2238 -27740
rect 4627 -27612 4713 -27517
rect 4628 -27749 4714 -27654
rect 12520 -30080 12600 -30000
rect 12640 -30080 12720 -30000
rect 12760 -30080 12840 -30000
rect 12520 -30200 12600 -30120
rect 12640 -30200 12720 -30120
rect 12760 -30200 12840 -30120
rect 12520 -30320 12600 -30240
rect 12640 -30320 12720 -30240
rect 12760 -30320 12840 -30240
rect 12520 -30440 12600 -30360
rect 12640 -30440 12720 -30360
rect 12760 -30440 12840 -30360
rect 12520 -34700 12600 -34620
rect 12640 -34700 12720 -34620
rect 12760 -34700 12840 -34620
rect 12520 -34800 12600 -34720
rect 12640 -34800 12720 -34720
rect 12760 -34800 12840 -34720
rect 12520 -34900 12600 -34820
rect 12640 -34900 12720 -34820
rect 12760 -34900 12840 -34820
rect 12520 -35000 12600 -34920
rect 12640 -35000 12720 -34920
rect 12760 -35000 12840 -34920
<< metal4 >>
rect 4619 -27374 4723 -27360
rect 4619 -27469 4626 -27374
rect 4713 -27469 4723 -27374
rect 4619 -27517 4723 -27469
rect 2144 -27620 2257 -27597
rect 2144 -27697 2160 -27620
rect 2238 -27659 2257 -27620
rect 4619 -27612 4627 -27517
rect 4713 -27612 4723 -27517
rect 4619 -27654 4723 -27612
rect 4619 -27657 4628 -27654
rect 3209 -27659 4628 -27657
rect 2238 -27697 4628 -27659
rect 2144 -27740 4628 -27697
rect 2144 -27818 2160 -27740
rect 2238 -27749 4628 -27740
rect 4714 -27749 4723 -27654
rect 2238 -27760 4723 -27749
rect 2238 -27818 2257 -27760
rect 2144 -27825 2257 -27818
rect 3209 -27761 4723 -27760
rect 3209 -27762 4720 -27761
rect 3209 -27886 3325 -27762
rect 3208 -27975 3325 -27886
rect 3208 -27977 3663 -27975
rect 3208 -28080 12242 -27977
rect 3208 -28141 3325 -28080
rect 3208 -32587 3321 -28141
rect 12500 -30000 12860 -29920
rect 12500 -30080 12520 -30000
rect 12600 -30080 12640 -30000
rect 12720 -30080 12760 -30000
rect 12840 -30080 12860 -30000
rect 12500 -30120 12860 -30080
rect 12500 -30200 12520 -30120
rect 12600 -30200 12640 -30120
rect 12720 -30200 12760 -30120
rect 12840 -30200 12860 -30120
rect 12140 -30240 12860 -30200
rect 12140 -30320 12520 -30240
rect 12600 -30320 12640 -30240
rect 12720 -30320 12760 -30240
rect 12840 -30320 12860 -30240
rect 12140 -30360 12860 -30320
rect 12140 -30420 12520 -30360
rect 12500 -30440 12520 -30420
rect 12600 -30440 12640 -30360
rect 12720 -30440 12760 -30360
rect 12840 -30440 12860 -30360
rect 12500 -30460 12860 -30440
rect 3208 -32688 12244 -32587
rect 12500 -34620 12860 -34560
rect 12500 -34700 12520 -34620
rect 12600 -34700 12640 -34620
rect 12720 -34700 12760 -34620
rect 12840 -34700 12860 -34620
rect 12500 -34720 12860 -34700
rect 12500 -34800 12520 -34720
rect 12600 -34800 12640 -34720
rect 12720 -34800 12760 -34720
rect 12840 -34800 12860 -34720
rect 12160 -34820 12860 -34800
rect 12160 -34900 12520 -34820
rect 12600 -34900 12640 -34820
rect 12720 -34900 12760 -34820
rect 12840 -34900 12860 -34820
rect 12160 -34920 12860 -34900
rect 12160 -35000 12520 -34920
rect 12600 -35000 12640 -34920
rect 12720 -35000 12760 -34920
rect 12840 -35000 12860 -34920
rect 12160 -35020 12860 -35000
use sky130_fd_pr__cap_mim_m3_1_VUG9HY  sky130_fd_pr__cap_mim_m3_1_VUG9HY_0
timestamp 1769400417
transform 0 -1 7920 1 0 -32468
box -4492 -4320 4492 4320
use sky130_fd_pr__nfet_01v8_UBWUWY  sky130_fd_pr__nfet_01v8_UBWUWY_0
timestamp 1769402310
transform 1 0 2196 0 1 -28498
box -436 -182 436 182
use sky130_fd_pr__pfet_01v8_GRDUQF  sky130_fd_pr__pfet_01v8_GRDUQF_0
timestamp 1769402310
transform 1 0 -1303 0 1 -26866
box -1297 -334 1297 368
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_0
timestamp 1769400417
transform 0 1 -1840 -1 0 -30221
box -141 -740 141 740
use sky130_fd_pr__nfet_01v8_9SDSBW  XM3
timestamp 1769406237
transform 1 0 337 0 1 -30003
box -337 -397 337 397
use sky130_fd_pr__pfet_01v8_GRDUQF  XM5
timestamp 1769402310
transform 1 0 2297 0 1 -26866
box -1297 -334 1297 368
use sky130_fd_pr__nfet_01v8_BU786C  XM9
timestamp 1769402310
transform 1 0 2183 0 1 -30003
box -183 -397 183 397
use sky130_fd_pr__pfet_01v8_3HNK2A  XM11
timestamp 1769406237
transform 1 0 9593 0 1 -26992
box -4993 -408 4993 442
use sky130_fd_pr__nfet_01v8_CH4F5S  XM12
timestamp 1769406237
transform 1 0 13865 0 1 -30093
box -645 -307 645 307
use sky130_fd_pr__nfet_01v8_T8V4TE  XM14
timestamp 1769400417
transform 1 0 402 0 1 -28506
box -73 -142 73 142
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  XR1
timestamp 1769400417
transform 0 1 -1831 -1 0 -28595
box -141 -740 141 740
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  XR2
timestamp 1769400417
transform 0 1 -1840 -1 0 -29021
box -141 -740 141 740
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  XR3
timestamp 1769400417
transform 0 1 -1840 -1 0 -29421
box -141 -740 141 740
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  XR4
timestamp 1769400417
transform 0 1 -1840 -1 0 -29821
box -141 -740 141 740
<< labels >>
flabel metal1 -3200 -24800 -3000 -24600 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 -3200 -32400 -3000 -32200 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 1200 -32800 1400 -32600 0 FreeSans 256 0 0 0 VP
port 2 nsew
flabel metal1 3000 -32800 3200 -32600 0 FreeSans 256 0 0 0 VN
port 3 nsew
flabel metal1 15400 -28600 15600 -28540 0 FreeSans 256 0 0 0 OUT
port 4 nsew
<< end >>
