magic
tech sky130A
magscale 1 2
timestamp 1770083657
<< error_s >>
rect 1234 2340 7466 2366
rect 1234 -160 1240 2340
rect 1300 2274 7400 2300
rect 1300 -94 1306 2274
rect 7374 -94 7400 2274
rect 1300 -100 7400 -94
rect 7440 -160 7466 2340
rect 1234 -166 7466 -160
<< nwell >>
rect 1240 -160 7440 2340
<< mvnsubdiff >>
rect 1300 2267 7400 2300
rect 1300 2233 1443 2267
rect 1477 2233 1511 2267
rect 1545 2233 1579 2267
rect 1613 2233 1647 2267
rect 1681 2233 1715 2267
rect 1749 2233 1783 2267
rect 1817 2233 1851 2267
rect 1885 2233 1919 2267
rect 1953 2233 1987 2267
rect 2021 2233 2055 2267
rect 2089 2233 2123 2267
rect 2157 2233 2191 2267
rect 2225 2233 2259 2267
rect 2293 2233 2327 2267
rect 2361 2233 2395 2267
rect 2429 2233 2463 2267
rect 2497 2233 2531 2267
rect 2565 2233 2599 2267
rect 2633 2233 2667 2267
rect 2701 2233 2735 2267
rect 2769 2233 2803 2267
rect 2837 2233 2871 2267
rect 2905 2233 2939 2267
rect 2973 2233 3007 2267
rect 3041 2233 3075 2267
rect 3109 2233 3143 2267
rect 3177 2233 3211 2267
rect 3245 2233 3279 2267
rect 3313 2233 3347 2267
rect 3381 2233 3415 2267
rect 3449 2233 3483 2267
rect 3517 2233 3551 2267
rect 3585 2233 3619 2267
rect 3653 2233 3687 2267
rect 3721 2233 3755 2267
rect 3789 2233 3823 2267
rect 3857 2233 3891 2267
rect 3925 2233 3959 2267
rect 3993 2233 4027 2267
rect 4061 2233 4095 2267
rect 4129 2233 4163 2267
rect 4197 2233 4231 2267
rect 4265 2233 4299 2267
rect 4333 2233 4367 2267
rect 4401 2233 4435 2267
rect 4469 2233 4503 2267
rect 4537 2233 4571 2267
rect 4605 2233 4639 2267
rect 4673 2233 4707 2267
rect 4741 2233 4775 2267
rect 4809 2233 4843 2267
rect 4877 2233 4911 2267
rect 4945 2233 4979 2267
rect 5013 2233 5047 2267
rect 5081 2233 5115 2267
rect 5149 2233 5183 2267
rect 5217 2233 5251 2267
rect 5285 2233 5319 2267
rect 5353 2233 5387 2267
rect 5421 2233 5455 2267
rect 5489 2233 5523 2267
rect 5557 2233 5591 2267
rect 5625 2233 5659 2267
rect 5693 2233 5727 2267
rect 5761 2233 5795 2267
rect 5829 2233 5863 2267
rect 5897 2233 5931 2267
rect 5965 2233 5999 2267
rect 6033 2233 6067 2267
rect 6101 2233 6135 2267
rect 6169 2233 6203 2267
rect 6237 2233 6271 2267
rect 6305 2233 6339 2267
rect 6373 2233 6407 2267
rect 6441 2233 6475 2267
rect 6509 2233 6543 2267
rect 6577 2233 6611 2267
rect 6645 2233 6679 2267
rect 6713 2233 6747 2267
rect 6781 2233 6815 2267
rect 6849 2233 6883 2267
rect 6917 2233 6951 2267
rect 6985 2233 7019 2267
rect 7053 2233 7087 2267
rect 7121 2233 7155 2267
rect 7189 2233 7223 2267
rect 7257 2233 7400 2267
rect 1300 2200 7400 2233
rect 1300 2171 1400 2200
rect 1300 2137 1333 2171
rect 1367 2137 1400 2171
rect 1300 2103 1400 2137
rect 1300 2069 1333 2103
rect 1367 2069 1400 2103
rect 1300 2035 1400 2069
rect 1300 2001 1333 2035
rect 1367 2001 1400 2035
rect 1300 1967 1400 2001
rect 1300 1933 1333 1967
rect 1367 1933 1400 1967
rect 1300 1899 1400 1933
rect 1300 1865 1333 1899
rect 1367 1865 1400 1899
rect 1300 1831 1400 1865
rect 1300 1797 1333 1831
rect 1367 1797 1400 1831
rect 1300 1763 1400 1797
rect 1300 1729 1333 1763
rect 1367 1729 1400 1763
rect 1300 1695 1400 1729
rect 1300 1661 1333 1695
rect 1367 1661 1400 1695
rect 1300 1627 1400 1661
rect 1300 1593 1333 1627
rect 1367 1593 1400 1627
rect 1300 1559 1400 1593
rect 1300 1525 1333 1559
rect 1367 1525 1400 1559
rect 1300 1491 1400 1525
rect 1300 1457 1333 1491
rect 1367 1457 1400 1491
rect 1300 1423 1400 1457
rect 1300 1389 1333 1423
rect 1367 1389 1400 1423
rect 1300 1355 1400 1389
rect 1300 1321 1333 1355
rect 1367 1321 1400 1355
rect 1300 1287 1400 1321
rect 1300 1253 1333 1287
rect 1367 1253 1400 1287
rect 1300 1219 1400 1253
rect 1300 1185 1333 1219
rect 1367 1185 1400 1219
rect 1300 1151 1400 1185
rect 1300 1117 1333 1151
rect 1367 1117 1400 1151
rect 1300 1083 1400 1117
rect 1300 1049 1333 1083
rect 1367 1049 1400 1083
rect 1300 1015 1400 1049
rect 1300 981 1333 1015
rect 1367 981 1400 1015
rect 1300 947 1400 981
rect 1300 913 1333 947
rect 1367 913 1400 947
rect 1300 879 1400 913
rect 1300 845 1333 879
rect 1367 845 1400 879
rect 1300 811 1400 845
rect 1300 777 1333 811
rect 1367 777 1400 811
rect 1300 743 1400 777
rect 1300 709 1333 743
rect 1367 709 1400 743
rect 1300 675 1400 709
rect 1300 641 1333 675
rect 1367 641 1400 675
rect 1300 607 1400 641
rect 1300 573 1333 607
rect 1367 573 1400 607
rect 1300 539 1400 573
rect 1300 505 1333 539
rect 1367 505 1400 539
rect 1300 471 1400 505
rect 1300 437 1333 471
rect 1367 437 1400 471
rect 1300 403 1400 437
rect 1300 369 1333 403
rect 1367 369 1400 403
rect 1300 335 1400 369
rect 1300 301 1333 335
rect 1367 301 1400 335
rect 1300 267 1400 301
rect 1300 233 1333 267
rect 1367 233 1400 267
rect 1300 199 1400 233
rect 1300 165 1333 199
rect 1367 165 1400 199
rect 1300 131 1400 165
rect 1300 97 1333 131
rect 1367 97 1400 131
rect 1300 63 1400 97
rect 1300 29 1333 63
rect 1367 29 1400 63
rect 1300 0 1400 29
rect 7300 2171 7400 2200
rect 7300 2137 7333 2171
rect 7367 2137 7400 2171
rect 7300 2103 7400 2137
rect 7300 2069 7333 2103
rect 7367 2069 7400 2103
rect 7300 2035 7400 2069
rect 7300 2001 7333 2035
rect 7367 2001 7400 2035
rect 7300 1967 7400 2001
rect 7300 1933 7333 1967
rect 7367 1933 7400 1967
rect 7300 1899 7400 1933
rect 7300 1865 7333 1899
rect 7367 1865 7400 1899
rect 7300 1831 7400 1865
rect 7300 1797 7333 1831
rect 7367 1797 7400 1831
rect 7300 1763 7400 1797
rect 7300 1729 7333 1763
rect 7367 1729 7400 1763
rect 7300 1695 7400 1729
rect 7300 1661 7333 1695
rect 7367 1661 7400 1695
rect 7300 1627 7400 1661
rect 7300 1593 7333 1627
rect 7367 1593 7400 1627
rect 7300 1559 7400 1593
rect 7300 1525 7333 1559
rect 7367 1525 7400 1559
rect 7300 1491 7400 1525
rect 7300 1457 7333 1491
rect 7367 1457 7400 1491
rect 7300 1423 7400 1457
rect 7300 1389 7333 1423
rect 7367 1389 7400 1423
rect 7300 1355 7400 1389
rect 7300 1321 7333 1355
rect 7367 1321 7400 1355
rect 7300 1287 7400 1321
rect 7300 1253 7333 1287
rect 7367 1253 7400 1287
rect 7300 1219 7400 1253
rect 7300 1185 7333 1219
rect 7367 1185 7400 1219
rect 7300 1151 7400 1185
rect 7300 1117 7333 1151
rect 7367 1117 7400 1151
rect 7300 1083 7400 1117
rect 7300 1049 7333 1083
rect 7367 1049 7400 1083
rect 7300 1015 7400 1049
rect 7300 981 7333 1015
rect 7367 981 7400 1015
rect 7300 947 7400 981
rect 7300 913 7333 947
rect 7367 913 7400 947
rect 7300 879 7400 913
rect 7300 845 7333 879
rect 7367 845 7400 879
rect 7300 811 7400 845
rect 7300 777 7333 811
rect 7367 777 7400 811
rect 7300 743 7400 777
rect 7300 709 7333 743
rect 7367 709 7400 743
rect 7300 675 7400 709
rect 7300 641 7333 675
rect 7367 641 7400 675
rect 7300 607 7400 641
rect 7300 573 7333 607
rect 7367 573 7400 607
rect 7300 539 7400 573
rect 7300 505 7333 539
rect 7367 505 7400 539
rect 7300 471 7400 505
rect 7300 437 7333 471
rect 7367 437 7400 471
rect 7300 403 7400 437
rect 7300 369 7333 403
rect 7367 369 7400 403
rect 7300 335 7400 369
rect 7300 301 7333 335
rect 7367 301 7400 335
rect 7300 267 7400 301
rect 7300 233 7333 267
rect 7367 233 7400 267
rect 7300 199 7400 233
rect 7300 165 7333 199
rect 7367 165 7400 199
rect 7300 131 7400 165
rect 7300 97 7333 131
rect 7367 97 7400 131
rect 7300 63 7400 97
rect 7300 29 7333 63
rect 7367 29 7400 63
rect 7300 0 7400 29
rect 1300 -33 7400 0
rect 1300 -67 1443 -33
rect 1477 -67 1511 -33
rect 1545 -67 1579 -33
rect 1613 -67 1647 -33
rect 1681 -67 1715 -33
rect 1749 -67 1783 -33
rect 1817 -67 1851 -33
rect 1885 -67 1919 -33
rect 1953 -67 1987 -33
rect 2021 -67 2055 -33
rect 2089 -67 2123 -33
rect 2157 -67 2191 -33
rect 2225 -67 2259 -33
rect 2293 -67 2327 -33
rect 2361 -67 2395 -33
rect 2429 -67 2463 -33
rect 2497 -67 2531 -33
rect 2565 -67 2599 -33
rect 2633 -67 2667 -33
rect 2701 -67 2735 -33
rect 2769 -67 2803 -33
rect 2837 -67 2871 -33
rect 2905 -67 2939 -33
rect 2973 -67 3007 -33
rect 3041 -67 3075 -33
rect 3109 -67 3143 -33
rect 3177 -67 3211 -33
rect 3245 -67 3279 -33
rect 3313 -67 3347 -33
rect 3381 -67 3415 -33
rect 3449 -67 3483 -33
rect 3517 -67 3551 -33
rect 3585 -67 3619 -33
rect 3653 -67 3687 -33
rect 3721 -67 3755 -33
rect 3789 -67 3823 -33
rect 3857 -67 3891 -33
rect 3925 -67 3959 -33
rect 3993 -67 4027 -33
rect 4061 -67 4095 -33
rect 4129 -67 4163 -33
rect 4197 -67 4231 -33
rect 4265 -67 4299 -33
rect 4333 -67 4367 -33
rect 4401 -67 4435 -33
rect 4469 -67 4503 -33
rect 4537 -67 4571 -33
rect 4605 -67 4639 -33
rect 4673 -67 4707 -33
rect 4741 -67 4775 -33
rect 4809 -67 4843 -33
rect 4877 -67 4911 -33
rect 4945 -67 4979 -33
rect 5013 -67 5047 -33
rect 5081 -67 5115 -33
rect 5149 -67 5183 -33
rect 5217 -67 5251 -33
rect 5285 -67 5319 -33
rect 5353 -67 5387 -33
rect 5421 -67 5455 -33
rect 5489 -67 5523 -33
rect 5557 -67 5591 -33
rect 5625 -67 5659 -33
rect 5693 -67 5727 -33
rect 5761 -67 5795 -33
rect 5829 -67 5863 -33
rect 5897 -67 5931 -33
rect 5965 -67 5999 -33
rect 6033 -67 6067 -33
rect 6101 -67 6135 -33
rect 6169 -67 6203 -33
rect 6237 -67 6271 -33
rect 6305 -67 6339 -33
rect 6373 -67 6407 -33
rect 6441 -67 6475 -33
rect 6509 -67 6543 -33
rect 6577 -67 6611 -33
rect 6645 -67 6679 -33
rect 6713 -67 6747 -33
rect 6781 -67 6815 -33
rect 6849 -67 6883 -33
rect 6917 -67 6951 -33
rect 6985 -67 7019 -33
rect 7053 -67 7087 -33
rect 7121 -67 7155 -33
rect 7189 -67 7223 -33
rect 7257 -67 7400 -33
rect 1300 -100 7400 -67
<< mvnsubdiffcont >>
rect 1443 2233 1477 2267
rect 1511 2233 1545 2267
rect 1579 2233 1613 2267
rect 1647 2233 1681 2267
rect 1715 2233 1749 2267
rect 1783 2233 1817 2267
rect 1851 2233 1885 2267
rect 1919 2233 1953 2267
rect 1987 2233 2021 2267
rect 2055 2233 2089 2267
rect 2123 2233 2157 2267
rect 2191 2233 2225 2267
rect 2259 2233 2293 2267
rect 2327 2233 2361 2267
rect 2395 2233 2429 2267
rect 2463 2233 2497 2267
rect 2531 2233 2565 2267
rect 2599 2233 2633 2267
rect 2667 2233 2701 2267
rect 2735 2233 2769 2267
rect 2803 2233 2837 2267
rect 2871 2233 2905 2267
rect 2939 2233 2973 2267
rect 3007 2233 3041 2267
rect 3075 2233 3109 2267
rect 3143 2233 3177 2267
rect 3211 2233 3245 2267
rect 3279 2233 3313 2267
rect 3347 2233 3381 2267
rect 3415 2233 3449 2267
rect 3483 2233 3517 2267
rect 3551 2233 3585 2267
rect 3619 2233 3653 2267
rect 3687 2233 3721 2267
rect 3755 2233 3789 2267
rect 3823 2233 3857 2267
rect 3891 2233 3925 2267
rect 3959 2233 3993 2267
rect 4027 2233 4061 2267
rect 4095 2233 4129 2267
rect 4163 2233 4197 2267
rect 4231 2233 4265 2267
rect 4299 2233 4333 2267
rect 4367 2233 4401 2267
rect 4435 2233 4469 2267
rect 4503 2233 4537 2267
rect 4571 2233 4605 2267
rect 4639 2233 4673 2267
rect 4707 2233 4741 2267
rect 4775 2233 4809 2267
rect 4843 2233 4877 2267
rect 4911 2233 4945 2267
rect 4979 2233 5013 2267
rect 5047 2233 5081 2267
rect 5115 2233 5149 2267
rect 5183 2233 5217 2267
rect 5251 2233 5285 2267
rect 5319 2233 5353 2267
rect 5387 2233 5421 2267
rect 5455 2233 5489 2267
rect 5523 2233 5557 2267
rect 5591 2233 5625 2267
rect 5659 2233 5693 2267
rect 5727 2233 5761 2267
rect 5795 2233 5829 2267
rect 5863 2233 5897 2267
rect 5931 2233 5965 2267
rect 5999 2233 6033 2267
rect 6067 2233 6101 2267
rect 6135 2233 6169 2267
rect 6203 2233 6237 2267
rect 6271 2233 6305 2267
rect 6339 2233 6373 2267
rect 6407 2233 6441 2267
rect 6475 2233 6509 2267
rect 6543 2233 6577 2267
rect 6611 2233 6645 2267
rect 6679 2233 6713 2267
rect 6747 2233 6781 2267
rect 6815 2233 6849 2267
rect 6883 2233 6917 2267
rect 6951 2233 6985 2267
rect 7019 2233 7053 2267
rect 7087 2233 7121 2267
rect 7155 2233 7189 2267
rect 7223 2233 7257 2267
rect 1333 2137 1367 2171
rect 1333 2069 1367 2103
rect 1333 2001 1367 2035
rect 1333 1933 1367 1967
rect 1333 1865 1367 1899
rect 1333 1797 1367 1831
rect 1333 1729 1367 1763
rect 1333 1661 1367 1695
rect 1333 1593 1367 1627
rect 1333 1525 1367 1559
rect 1333 1457 1367 1491
rect 1333 1389 1367 1423
rect 1333 1321 1367 1355
rect 1333 1253 1367 1287
rect 1333 1185 1367 1219
rect 1333 1117 1367 1151
rect 1333 1049 1367 1083
rect 1333 981 1367 1015
rect 1333 913 1367 947
rect 1333 845 1367 879
rect 1333 777 1367 811
rect 1333 709 1367 743
rect 1333 641 1367 675
rect 1333 573 1367 607
rect 1333 505 1367 539
rect 1333 437 1367 471
rect 1333 369 1367 403
rect 1333 301 1367 335
rect 1333 233 1367 267
rect 1333 165 1367 199
rect 1333 97 1367 131
rect 1333 29 1367 63
rect 7333 2137 7367 2171
rect 7333 2069 7367 2103
rect 7333 2001 7367 2035
rect 7333 1933 7367 1967
rect 7333 1865 7367 1899
rect 7333 1797 7367 1831
rect 7333 1729 7367 1763
rect 7333 1661 7367 1695
rect 7333 1593 7367 1627
rect 7333 1525 7367 1559
rect 7333 1457 7367 1491
rect 7333 1389 7367 1423
rect 7333 1321 7367 1355
rect 7333 1253 7367 1287
rect 7333 1185 7367 1219
rect 7333 1117 7367 1151
rect 7333 1049 7367 1083
rect 7333 981 7367 1015
rect 7333 913 7367 947
rect 7333 845 7367 879
rect 7333 777 7367 811
rect 7333 709 7367 743
rect 7333 641 7367 675
rect 7333 573 7367 607
rect 7333 505 7367 539
rect 7333 437 7367 471
rect 7333 369 7367 403
rect 7333 301 7367 335
rect 7333 233 7367 267
rect 7333 165 7367 199
rect 7333 97 7367 131
rect 7333 29 7367 63
rect 1443 -67 1477 -33
rect 1511 -67 1545 -33
rect 1579 -67 1613 -33
rect 1647 -67 1681 -33
rect 1715 -67 1749 -33
rect 1783 -67 1817 -33
rect 1851 -67 1885 -33
rect 1919 -67 1953 -33
rect 1987 -67 2021 -33
rect 2055 -67 2089 -33
rect 2123 -67 2157 -33
rect 2191 -67 2225 -33
rect 2259 -67 2293 -33
rect 2327 -67 2361 -33
rect 2395 -67 2429 -33
rect 2463 -67 2497 -33
rect 2531 -67 2565 -33
rect 2599 -67 2633 -33
rect 2667 -67 2701 -33
rect 2735 -67 2769 -33
rect 2803 -67 2837 -33
rect 2871 -67 2905 -33
rect 2939 -67 2973 -33
rect 3007 -67 3041 -33
rect 3075 -67 3109 -33
rect 3143 -67 3177 -33
rect 3211 -67 3245 -33
rect 3279 -67 3313 -33
rect 3347 -67 3381 -33
rect 3415 -67 3449 -33
rect 3483 -67 3517 -33
rect 3551 -67 3585 -33
rect 3619 -67 3653 -33
rect 3687 -67 3721 -33
rect 3755 -67 3789 -33
rect 3823 -67 3857 -33
rect 3891 -67 3925 -33
rect 3959 -67 3993 -33
rect 4027 -67 4061 -33
rect 4095 -67 4129 -33
rect 4163 -67 4197 -33
rect 4231 -67 4265 -33
rect 4299 -67 4333 -33
rect 4367 -67 4401 -33
rect 4435 -67 4469 -33
rect 4503 -67 4537 -33
rect 4571 -67 4605 -33
rect 4639 -67 4673 -33
rect 4707 -67 4741 -33
rect 4775 -67 4809 -33
rect 4843 -67 4877 -33
rect 4911 -67 4945 -33
rect 4979 -67 5013 -33
rect 5047 -67 5081 -33
rect 5115 -67 5149 -33
rect 5183 -67 5217 -33
rect 5251 -67 5285 -33
rect 5319 -67 5353 -33
rect 5387 -67 5421 -33
rect 5455 -67 5489 -33
rect 5523 -67 5557 -33
rect 5591 -67 5625 -33
rect 5659 -67 5693 -33
rect 5727 -67 5761 -33
rect 5795 -67 5829 -33
rect 5863 -67 5897 -33
rect 5931 -67 5965 -33
rect 5999 -67 6033 -33
rect 6067 -67 6101 -33
rect 6135 -67 6169 -33
rect 6203 -67 6237 -33
rect 6271 -67 6305 -33
rect 6339 -67 6373 -33
rect 6407 -67 6441 -33
rect 6475 -67 6509 -33
rect 6543 -67 6577 -33
rect 6611 -67 6645 -33
rect 6679 -67 6713 -33
rect 6747 -67 6781 -33
rect 6815 -67 6849 -33
rect 6883 -67 6917 -33
rect 6951 -67 6985 -33
rect 7019 -67 7053 -33
rect 7087 -67 7121 -33
rect 7155 -67 7189 -33
rect 7223 -67 7257 -33
<< locali >>
rect 1300 2267 7400 2300
rect 1300 2233 1443 2267
rect 1477 2233 1511 2267
rect 1545 2233 1579 2267
rect 1613 2233 1647 2267
rect 1681 2233 1715 2267
rect 1749 2233 1783 2267
rect 1817 2233 1851 2267
rect 1885 2233 1919 2267
rect 1953 2233 1987 2267
rect 2021 2233 2055 2267
rect 2089 2233 2123 2267
rect 2157 2233 2191 2267
rect 2225 2233 2259 2267
rect 2293 2233 2327 2267
rect 2361 2233 2395 2267
rect 2429 2233 2463 2267
rect 2497 2233 2531 2267
rect 2565 2233 2599 2267
rect 2633 2233 2667 2267
rect 2701 2233 2735 2267
rect 2769 2233 2803 2267
rect 2837 2233 2871 2267
rect 2905 2233 2939 2267
rect 2973 2233 3007 2267
rect 3041 2233 3075 2267
rect 3109 2233 3143 2267
rect 3177 2233 3211 2267
rect 3245 2233 3279 2267
rect 3313 2233 3347 2267
rect 3381 2233 3415 2267
rect 3449 2233 3483 2267
rect 3517 2233 3551 2267
rect 3585 2233 3619 2267
rect 3653 2233 3687 2267
rect 3721 2233 3755 2267
rect 3789 2233 3823 2267
rect 3857 2233 3891 2267
rect 3925 2233 3959 2267
rect 3993 2233 4027 2267
rect 4061 2233 4095 2267
rect 4129 2233 4163 2267
rect 4197 2233 4231 2267
rect 4265 2233 4299 2267
rect 4333 2233 4367 2267
rect 4401 2233 4435 2267
rect 4469 2233 4503 2267
rect 4537 2233 4571 2267
rect 4605 2233 4639 2267
rect 4673 2233 4707 2267
rect 4741 2233 4775 2267
rect 4809 2233 4843 2267
rect 4877 2233 4911 2267
rect 4945 2233 4979 2267
rect 5013 2233 5047 2267
rect 5081 2233 5115 2267
rect 5149 2233 5183 2267
rect 5217 2233 5251 2267
rect 5285 2233 5319 2267
rect 5353 2233 5387 2267
rect 5421 2233 5455 2267
rect 5489 2233 5523 2267
rect 5557 2233 5591 2267
rect 5625 2233 5659 2267
rect 5693 2233 5727 2267
rect 5761 2233 5795 2267
rect 5829 2233 5863 2267
rect 5897 2233 5931 2267
rect 5965 2233 5999 2267
rect 6033 2233 6067 2267
rect 6101 2233 6135 2267
rect 6169 2233 6203 2267
rect 6237 2233 6271 2267
rect 6305 2233 6339 2267
rect 6373 2233 6407 2267
rect 6441 2233 6475 2267
rect 6509 2233 6543 2267
rect 6577 2233 6611 2267
rect 6645 2233 6679 2267
rect 6713 2233 6747 2267
rect 6781 2233 6815 2267
rect 6849 2233 6883 2267
rect 6917 2233 6951 2267
rect 6985 2233 7019 2267
rect 7053 2233 7087 2267
rect 7121 2233 7155 2267
rect 7189 2233 7223 2267
rect 7257 2233 7400 2267
rect 1300 2200 7400 2233
rect 1300 2171 1400 2200
rect 1300 2137 1333 2171
rect 1367 2137 1400 2171
rect 1300 2103 1400 2137
rect 1300 2069 1333 2103
rect 1367 2069 1400 2103
rect 1300 2035 1400 2069
rect 1300 2001 1333 2035
rect 1367 2001 1400 2035
rect 1300 1967 1400 2001
rect 1300 1933 1333 1967
rect 1367 1933 1400 1967
rect 1300 1899 1400 1933
rect 1300 1865 1333 1899
rect 1367 1865 1400 1899
rect 1300 1831 1400 1865
rect 1300 1797 1333 1831
rect 1367 1797 1400 1831
rect 1300 1763 1400 1797
rect 1300 1729 1333 1763
rect 1367 1729 1400 1763
rect 1300 1695 1400 1729
rect 1300 1661 1333 1695
rect 1367 1661 1400 1695
rect 1300 1627 1400 1661
rect 1300 1593 1333 1627
rect 1367 1593 1400 1627
rect 1300 1559 1400 1593
rect 1300 1525 1333 1559
rect 1367 1525 1400 1559
rect 1300 1491 1400 1525
rect 1300 1457 1333 1491
rect 1367 1457 1400 1491
rect 1300 1423 1400 1457
rect 1300 1389 1333 1423
rect 1367 1389 1400 1423
rect 1300 1355 1400 1389
rect 1300 1321 1333 1355
rect 1367 1321 1400 1355
rect 1300 1287 1400 1321
rect 1300 1253 1333 1287
rect 1367 1253 1400 1287
rect 1300 1219 1400 1253
rect 1300 1185 1333 1219
rect 1367 1185 1400 1219
rect 1300 1151 1400 1185
rect 1300 1117 1333 1151
rect 1367 1117 1400 1151
rect 1300 1083 1400 1117
rect 1300 1049 1333 1083
rect 1367 1049 1400 1083
rect 1300 1015 1400 1049
rect 1300 981 1333 1015
rect 1367 981 1400 1015
rect 1300 947 1400 981
rect 1300 913 1333 947
rect 1367 913 1400 947
rect 1300 879 1400 913
rect 1300 845 1333 879
rect 1367 845 1400 879
rect 1300 811 1400 845
rect 1300 777 1333 811
rect 1367 777 1400 811
rect 1300 743 1400 777
rect 1300 709 1333 743
rect 1367 709 1400 743
rect 1300 675 1400 709
rect 1300 641 1333 675
rect 1367 641 1400 675
rect 1300 607 1400 641
rect 1300 573 1333 607
rect 1367 573 1400 607
rect 1300 539 1400 573
rect 1300 505 1333 539
rect 1367 505 1400 539
rect 1300 471 1400 505
rect 1300 437 1333 471
rect 1367 437 1400 471
rect 1300 403 1400 437
rect 1300 369 1333 403
rect 1367 369 1400 403
rect 1300 335 1400 369
rect 1300 301 1333 335
rect 1367 301 1400 335
rect 1300 267 1400 301
rect 1300 233 1333 267
rect 1367 233 1400 267
rect 1300 199 1400 233
rect 1300 165 1333 199
rect 1367 165 1400 199
rect 1300 131 1400 165
rect 1300 97 1333 131
rect 1367 97 1400 131
rect 1300 63 1400 97
rect 1560 160 1860 2080
rect 2120 200 2240 2200
rect 2740 200 2860 2200
rect 3040 160 3160 2080
rect 3360 200 3480 2200
rect 3960 200 4080 2200
rect 4280 260 4400 2080
rect 4200 160 4500 260
rect 4580 200 4700 2200
rect 5200 200 5320 2200
rect 5500 160 5620 2080
rect 5820 200 5940 2200
rect 6440 200 6560 2200
rect 7300 2171 7400 2200
rect 7300 2137 7333 2171
rect 7367 2137 7400 2171
rect 7300 2103 7400 2137
rect 6800 160 7100 2080
rect 1560 117 7100 160
rect 1560 83 4323 117
rect 4357 83 7100 117
rect 1560 80 7100 83
rect 7300 2069 7333 2103
rect 7367 2069 7400 2103
rect 7300 2035 7400 2069
rect 7300 2001 7333 2035
rect 7367 2001 7400 2035
rect 7300 1967 7400 2001
rect 7300 1933 7333 1967
rect 7367 1933 7400 1967
rect 7300 1899 7400 1933
rect 7300 1865 7333 1899
rect 7367 1865 7400 1899
rect 7300 1831 7400 1865
rect 7300 1797 7333 1831
rect 7367 1797 7400 1831
rect 7300 1763 7400 1797
rect 7300 1729 7333 1763
rect 7367 1729 7400 1763
rect 7300 1695 7400 1729
rect 7300 1661 7333 1695
rect 7367 1661 7400 1695
rect 7300 1627 7400 1661
rect 7300 1593 7333 1627
rect 7367 1593 7400 1627
rect 7300 1559 7400 1593
rect 7300 1525 7333 1559
rect 7367 1525 7400 1559
rect 7300 1491 7400 1525
rect 7300 1457 7333 1491
rect 7367 1457 7400 1491
rect 7300 1423 7400 1457
rect 7300 1389 7333 1423
rect 7367 1389 7400 1423
rect 7300 1355 7400 1389
rect 7300 1321 7333 1355
rect 7367 1321 7400 1355
rect 7300 1287 7400 1321
rect 7300 1253 7333 1287
rect 7367 1253 7400 1287
rect 7300 1219 7400 1253
rect 7300 1185 7333 1219
rect 7367 1185 7400 1219
rect 7300 1151 7400 1185
rect 7300 1117 7333 1151
rect 7367 1117 7400 1151
rect 7300 1083 7400 1117
rect 7300 1049 7333 1083
rect 7367 1049 7400 1083
rect 7300 1015 7400 1049
rect 7300 981 7333 1015
rect 7367 981 7400 1015
rect 7300 947 7400 981
rect 7300 913 7333 947
rect 7367 913 7400 947
rect 7300 879 7400 913
rect 7300 845 7333 879
rect 7367 845 7400 879
rect 7300 811 7400 845
rect 7300 777 7333 811
rect 7367 777 7400 811
rect 7300 743 7400 777
rect 7300 709 7333 743
rect 7367 709 7400 743
rect 7300 675 7400 709
rect 7300 641 7333 675
rect 7367 641 7400 675
rect 7300 607 7400 641
rect 7300 573 7333 607
rect 7367 573 7400 607
rect 7300 539 7400 573
rect 7300 505 7333 539
rect 7367 505 7400 539
rect 7300 471 7400 505
rect 7300 437 7333 471
rect 7367 437 7400 471
rect 7300 403 7400 437
rect 7300 369 7333 403
rect 7367 369 7400 403
rect 7300 335 7400 369
rect 7300 301 7333 335
rect 7367 301 7400 335
rect 7300 267 7400 301
rect 7300 233 7333 267
rect 7367 233 7400 267
rect 7300 199 7400 233
rect 7300 165 7333 199
rect 7367 165 7400 199
rect 7300 131 7400 165
rect 7300 97 7333 131
rect 7367 97 7400 131
rect 1300 29 1333 63
rect 1367 29 1400 63
rect 4200 40 4500 80
rect 7300 63 7400 97
rect 1300 0 1400 29
rect 7300 29 7333 63
rect 7367 29 7400 63
rect 7300 0 7400 29
rect 1300 -33 7400 0
rect 1300 -67 1333 -33
rect 1367 -67 1443 -33
rect 1477 -67 1511 -33
rect 1545 -67 1579 -33
rect 1613 -67 1647 -33
rect 1681 -67 1715 -33
rect 1749 -67 1783 -33
rect 1817 -67 1851 -33
rect 1885 -67 1919 -33
rect 1953 -67 1987 -33
rect 2021 -67 2055 -33
rect 2089 -67 2123 -33
rect 2157 -67 2191 -33
rect 2225 -67 2259 -33
rect 2293 -67 2327 -33
rect 2361 -67 2395 -33
rect 2429 -67 2463 -33
rect 2497 -67 2531 -33
rect 2565 -67 2599 -33
rect 2633 -67 2667 -33
rect 2701 -67 2735 -33
rect 2769 -67 2803 -33
rect 2837 -67 2871 -33
rect 2905 -67 2939 -33
rect 2973 -67 3007 -33
rect 3041 -67 3075 -33
rect 3109 -67 3143 -33
rect 3177 -67 3211 -33
rect 3245 -67 3279 -33
rect 3313 -67 3347 -33
rect 3381 -67 3415 -33
rect 3449 -67 3483 -33
rect 3517 -67 3551 -33
rect 3585 -67 3619 -33
rect 3653 -67 3687 -33
rect 3721 -67 3755 -33
rect 3789 -67 3823 -33
rect 3857 -67 3891 -33
rect 3925 -67 3959 -33
rect 3993 -67 4027 -33
rect 4061 -67 4095 -33
rect 4129 -67 4163 -33
rect 4197 -67 4231 -33
rect 4265 -67 4299 -33
rect 4333 -67 4367 -33
rect 4401 -67 4435 -33
rect 4469 -67 4503 -33
rect 4537 -67 4571 -33
rect 4605 -67 4639 -33
rect 4673 -67 4707 -33
rect 4741 -67 4775 -33
rect 4809 -67 4843 -33
rect 4877 -67 4911 -33
rect 4945 -67 4979 -33
rect 5013 -67 5047 -33
rect 5081 -67 5115 -33
rect 5149 -67 5183 -33
rect 5217 -67 5251 -33
rect 5285 -67 5319 -33
rect 5353 -67 5387 -33
rect 5421 -67 5455 -33
rect 5489 -67 5523 -33
rect 5557 -67 5591 -33
rect 5625 -67 5659 -33
rect 5693 -67 5727 -33
rect 5761 -67 5795 -33
rect 5829 -67 5863 -33
rect 5897 -67 5931 -33
rect 5965 -67 5999 -33
rect 6033 -67 6067 -33
rect 6101 -67 6135 -33
rect 6169 -67 6203 -33
rect 6237 -67 6271 -33
rect 6305 -67 6339 -33
rect 6373 -67 6407 -33
rect 6441 -67 6475 -33
rect 6509 -67 6543 -33
rect 6577 -67 6611 -33
rect 6645 -67 6679 -33
rect 6713 -67 6747 -33
rect 6781 -67 6815 -33
rect 6849 -67 6883 -33
rect 6917 -67 6951 -33
rect 6985 -67 7019 -33
rect 7053 -67 7087 -33
rect 7121 -67 7155 -33
rect 7189 -67 7223 -33
rect 7257 -67 7400 -33
rect 1300 -100 7400 -67
rect 4200 -233 4500 -220
rect 4200 -267 4233 -233
rect 4267 -267 4333 -233
rect 4367 -267 4433 -233
rect 4467 -267 4500 -233
rect 4200 -333 4500 -267
rect 4200 -367 4233 -333
rect 4267 -367 4333 -333
rect 4367 -367 4433 -333
rect 4467 -367 4500 -333
rect 4200 -433 4500 -367
rect 4200 -467 4233 -433
rect 4267 -467 4333 -433
rect 4367 -467 4433 -433
rect 4467 -467 4500 -433
rect 4200 -500 4500 -467
<< viali >>
rect 4323 83 4357 117
rect 1333 -67 1367 -33
rect 4233 -267 4267 -233
rect 4333 -267 4367 -233
rect 4433 -267 4467 -233
rect 4233 -367 4267 -333
rect 4333 -367 4367 -333
rect 4433 -367 4467 -333
rect 4233 -467 4267 -433
rect 4333 -467 4367 -433
rect 4433 -467 4467 -433
<< metal1 >>
rect 900 1276 1200 1300
rect 900 1224 924 1276
rect 976 1224 1024 1276
rect 1076 1224 1124 1276
rect 1176 1224 1200 1276
rect 900 1176 1200 1224
rect 900 1124 924 1176
rect 976 1124 1024 1176
rect 1076 1124 1124 1176
rect 1176 1124 1200 1176
rect 900 1076 1200 1124
rect 900 1024 924 1076
rect 976 1024 1024 1076
rect 1076 1024 1124 1076
rect 1176 1024 1200 1076
rect 900 1000 1200 1024
rect 2400 1276 2600 1300
rect 2400 1224 2424 1276
rect 2476 1224 2524 1276
rect 2576 1224 2600 1276
rect 2400 1176 2600 1224
rect 2400 1124 2424 1176
rect 2476 1124 2524 1176
rect 2576 1124 2600 1176
rect 2400 1076 2600 1124
rect 2400 1024 2424 1076
rect 2476 1024 2524 1076
rect 2576 1024 2600 1076
rect 2400 1000 2600 1024
rect 3600 1276 3800 1300
rect 3600 1224 3624 1276
rect 3676 1224 3724 1276
rect 3776 1224 3800 1276
rect 3600 1176 3800 1224
rect 3600 1124 3624 1176
rect 3676 1124 3724 1176
rect 3776 1124 3800 1176
rect 3600 1076 3800 1124
rect 3600 1024 3624 1076
rect 3676 1024 3724 1076
rect 3776 1024 3800 1076
rect 3600 1000 3800 1024
rect 4860 1276 5060 1300
rect 4860 1224 4884 1276
rect 4936 1224 4984 1276
rect 5036 1224 5060 1276
rect 4860 1176 5060 1224
rect 4860 1124 4884 1176
rect 4936 1124 4984 1176
rect 5036 1124 5060 1176
rect 4860 1076 5060 1124
rect 4860 1024 4884 1076
rect 4936 1024 4984 1076
rect 5036 1024 5060 1076
rect 4860 1000 5060 1024
rect 6100 1276 6300 1300
rect 6100 1224 6124 1276
rect 6176 1224 6224 1276
rect 6276 1224 6300 1276
rect 6100 1176 6300 1224
rect 6100 1124 6124 1176
rect 6176 1124 6224 1176
rect 6276 1124 6300 1176
rect 6100 1076 6300 1124
rect 6100 1024 6124 1076
rect 6176 1024 6224 1076
rect 6276 1024 6300 1076
rect 6100 1000 6300 1024
rect 7500 1276 7800 1300
rect 7500 1224 7524 1276
rect 7576 1224 7624 1276
rect 7676 1224 7724 1276
rect 7776 1224 7800 1276
rect 7500 1176 7800 1224
rect 7500 1124 7524 1176
rect 7576 1124 7624 1176
rect 7676 1124 7724 1176
rect 7776 1124 7800 1176
rect 7500 1076 7800 1124
rect 7500 1024 7524 1076
rect 7576 1024 7624 1076
rect 7676 1024 7724 1076
rect 7776 1024 7800 1076
rect 7500 1000 7800 1024
rect 4200 117 4500 260
rect 4200 83 4323 117
rect 4357 83 4500 117
rect 1300 -33 1400 0
rect 1300 -67 1333 -33
rect 1367 -67 1400 -33
rect 1300 -100 1400 -67
rect 4200 -233 4500 83
rect 4200 -267 4233 -233
rect 4267 -267 4333 -233
rect 4367 -267 4433 -233
rect 4467 -267 4500 -233
rect 4200 -333 4500 -267
rect 4200 -367 4233 -333
rect 4267 -367 4333 -333
rect 4367 -367 4433 -333
rect 4467 -367 4500 -333
rect 4200 -433 4500 -367
rect 4200 -467 4233 -433
rect 4267 -467 4333 -433
rect 4367 -467 4433 -433
rect 4467 -467 4500 -433
rect 4200 -500 4500 -467
<< via1 >>
rect 924 1224 976 1276
rect 1024 1224 1076 1276
rect 1124 1224 1176 1276
rect 924 1124 976 1176
rect 1024 1124 1076 1176
rect 1124 1124 1176 1176
rect 924 1024 976 1076
rect 1024 1024 1076 1076
rect 1124 1024 1176 1076
rect 2424 1224 2476 1276
rect 2524 1224 2576 1276
rect 2424 1124 2476 1176
rect 2524 1124 2576 1176
rect 2424 1024 2476 1076
rect 2524 1024 2576 1076
rect 3624 1224 3676 1276
rect 3724 1224 3776 1276
rect 3624 1124 3676 1176
rect 3724 1124 3776 1176
rect 3624 1024 3676 1076
rect 3724 1024 3776 1076
rect 4884 1224 4936 1276
rect 4984 1224 5036 1276
rect 4884 1124 4936 1176
rect 4984 1124 5036 1176
rect 4884 1024 4936 1076
rect 4984 1024 5036 1076
rect 6124 1224 6176 1276
rect 6224 1224 6276 1276
rect 6124 1124 6176 1176
rect 6224 1124 6276 1176
rect 6124 1024 6176 1076
rect 6224 1024 6276 1076
rect 7524 1224 7576 1276
rect 7624 1224 7676 1276
rect 7724 1224 7776 1276
rect 7524 1124 7576 1176
rect 7624 1124 7676 1176
rect 7724 1124 7776 1176
rect 7524 1024 7576 1076
rect 7624 1024 7676 1076
rect 7724 1024 7776 1076
<< metal2 >>
rect 900 1276 7800 1300
rect 900 1224 924 1276
rect 976 1224 1024 1276
rect 1076 1224 1124 1276
rect 1176 1224 2424 1276
rect 2476 1224 2524 1276
rect 2576 1224 3624 1276
rect 3676 1224 3724 1276
rect 3776 1224 4884 1276
rect 4936 1224 4984 1276
rect 5036 1224 6124 1276
rect 6176 1224 6224 1276
rect 6276 1224 7524 1276
rect 7576 1224 7624 1276
rect 7676 1224 7724 1276
rect 7776 1224 7800 1276
rect 900 1176 7800 1224
rect 900 1124 924 1176
rect 976 1124 1024 1176
rect 1076 1124 1124 1176
rect 1176 1124 2424 1176
rect 2476 1124 2524 1176
rect 2576 1124 3624 1176
rect 3676 1124 3724 1176
rect 3776 1124 4884 1176
rect 4936 1124 4984 1176
rect 5036 1124 6124 1176
rect 6176 1124 6224 1176
rect 6276 1124 7524 1176
rect 7576 1124 7624 1176
rect 7676 1124 7724 1176
rect 7776 1124 7800 1176
rect 900 1076 7800 1124
rect 900 1024 924 1076
rect 976 1024 1024 1076
rect 1076 1024 1124 1076
rect 1176 1024 2424 1076
rect 2476 1024 2524 1076
rect 2576 1024 3624 1076
rect 3676 1024 3724 1076
rect 3776 1024 4884 1076
rect 4936 1024 4984 1076
rect 5036 1024 6124 1076
rect 6176 1024 6224 1076
rect 6276 1024 7524 1076
rect 7576 1024 7624 1076
rect 7676 1024 7724 1076
rect 7776 1024 7800 1076
rect 900 1000 7800 1024
use sky130_fd_pr__pfet_g5v0d10v5_ZPXM7F  XM2
timestamp 1770083657
transform 1 0 4337 0 1 1104
box -2867 -1004 2867 1042
<< labels >>
flabel metal1 s 1300 -100 1400 0 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal1 s 4300 -400 4400 -300 0 FreeSans 320 0 0 0 D1
port 2 nsew
flabel metal1 s 1000 1100 1100 1200 0 FreeSans 320 0 0 0 D2
port 3 nsew
<< end >>
