magic
tech sky130A
magscale 1 2
timestamp 1769616064
<< error_p >>
rect -496 -254 -428 -248
rect -188 -254 -120 -248
rect 120 -254 188 -248
rect 428 -254 496 -248
rect -496 -288 -484 -254
rect -188 -288 -176 -254
rect 120 -288 132 -254
rect 428 -288 440 -254
rect -496 -294 -428 -288
rect -188 -294 -120 -288
rect 120 -294 188 -288
rect 428 -294 496 -288
<< nwell >>
rect -845 -505 845 505
<< mvpmos >>
rect -587 -207 -337 279
rect -279 -207 -29 279
rect 29 -207 279 279
rect 337 -207 587 279
<< mvpdiff >>
rect -645 267 -587 279
rect -645 -195 -633 267
rect -599 -195 -587 267
rect -645 -207 -587 -195
rect -337 267 -279 279
rect -337 -195 -325 267
rect -291 -195 -279 267
rect -337 -207 -279 -195
rect -29 267 29 279
rect -29 -195 -17 267
rect 17 -195 29 267
rect -29 -207 29 -195
rect 279 267 337 279
rect 279 -195 291 267
rect 325 -195 337 267
rect 279 -207 337 -195
rect 587 267 645 279
rect 587 -195 599 267
rect 633 -195 645 267
rect 587 -207 645 -195
<< mvpdiffc >>
rect -633 -195 -599 267
rect -325 -195 -291 267
rect -17 -195 17 267
rect 291 -195 325 267
rect 599 -195 633 267
<< mvnsubdiff >>
rect -779 427 779 439
rect -779 393 -671 427
rect 671 393 779 427
rect -779 381 779 393
rect -779 -381 -721 381
rect 721 -381 779 381
rect -779 -439 779 -381
<< mvnsubdiffcont >>
rect -671 393 671 427
<< poly >>
rect -587 279 -337 305
rect -279 279 -29 305
rect 29 279 279 305
rect 337 279 587 305
rect -587 -254 -337 -207
rect -587 -271 -484 -254
rect -500 -288 -484 -271
rect -440 -271 -337 -254
rect -279 -254 -29 -207
rect -279 -271 -176 -254
rect -440 -288 -424 -271
rect -500 -304 -424 -288
rect -192 -288 -176 -271
rect -132 -271 -29 -254
rect 29 -254 279 -207
rect 29 -271 132 -254
rect -132 -288 -116 -271
rect -192 -304 -116 -288
rect 116 -288 132 -271
rect 176 -271 279 -254
rect 337 -254 587 -207
rect 337 -271 440 -254
rect 176 -288 192 -271
rect 116 -304 192 -288
rect 424 -288 440 -271
rect 484 -271 587 -254
rect 484 -288 500 -271
rect 424 -304 500 -288
<< polycont >>
rect -484 -288 -440 -254
rect -176 -288 -132 -254
rect 132 -288 176 -254
rect 440 -288 484 -254
<< locali >>
rect -687 393 -671 427
rect 671 393 687 427
rect -633 267 -599 283
rect -633 -211 -599 -195
rect -325 267 -291 283
rect -325 -211 -291 -195
rect -17 267 17 283
rect -17 -211 17 -195
rect 291 267 325 283
rect 291 -211 325 -195
rect 599 267 633 283
rect 599 -211 633 -195
rect -500 -288 -484 -254
rect -440 -288 -424 -254
rect -192 -288 -176 -254
rect -132 -288 -116 -254
rect 116 -288 132 -254
rect 176 -288 192 -254
rect 424 -288 440 -254
rect 484 -288 500 -254
<< viali >>
rect -633 -195 -599 267
rect -325 -195 -291 267
rect -17 -195 17 267
rect 291 -195 325 267
rect 599 -195 633 267
rect -484 -288 -440 -254
rect -176 -288 -132 -254
rect 132 -288 176 -254
rect 440 -288 484 -254
<< metal1 >>
rect -639 267 -593 279
rect -639 -195 -633 267
rect -599 -195 -593 267
rect -639 -207 -593 -195
rect -331 267 -285 279
rect -331 -195 -325 267
rect -291 -195 -285 267
rect -331 -207 -285 -195
rect -23 267 23 279
rect -23 -195 -17 267
rect 17 -195 23 267
rect -23 -207 23 -195
rect 285 267 331 279
rect 285 -195 291 267
rect 325 -195 331 267
rect 285 -207 331 -195
rect 593 267 639 279
rect 593 -195 599 267
rect 633 -195 639 267
rect 593 -207 639 -195
rect -496 -254 -428 -248
rect -496 -288 -484 -254
rect -440 -288 -428 -254
rect -496 -294 -428 -288
rect -188 -254 -120 -248
rect -188 -288 -176 -254
rect -132 -288 -120 -254
rect -188 -294 -120 -288
rect 120 -254 188 -248
rect 120 -288 132 -254
rect 176 -288 188 -254
rect 120 -294 188 -288
rect 428 -254 496 -248
rect 428 -288 440 -254
rect 484 -288 496 -254
rect 428 -294 496 -288
<< properties >>
string FIXED_BBOX -750 -410 750 410
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.425 l 1.25 m 1 nf 4 diffcov 100 polycov 20 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
