magic
tech sky130A
magscale 1 2
timestamp 1770112220
<< mvnmos >>
rect -129 -781 -29 719
rect 29 -781 129 719
<< mvndiff >>
rect -187 707 -129 719
rect -187 -769 -175 707
rect -141 -769 -129 707
rect -187 -781 -129 -769
rect -29 707 29 719
rect -29 -769 -17 707
rect 17 -769 29 707
rect -29 -781 29 -769
rect 129 707 187 719
rect 129 -769 141 707
rect 175 -769 187 707
rect 129 -781 187 -769
<< mvndiffc >>
rect -175 -769 -141 707
rect -17 -769 17 707
rect 141 -769 175 707
<< poly >>
rect -129 791 -29 807
rect -129 757 -113 791
rect -45 757 -29 791
rect -129 719 -29 757
rect 29 791 129 807
rect 29 757 45 791
rect 113 757 129 791
rect 29 719 129 757
rect -129 -807 -29 -781
rect 29 -807 129 -781
<< polycont >>
rect -113 757 -45 791
rect 45 757 113 791
<< locali >>
rect -129 757 -113 791
rect -45 757 -29 791
rect 29 757 45 791
rect 113 757 129 791
rect -175 707 -141 723
rect -175 -785 -141 -769
rect -17 707 17 723
rect -17 -785 17 -769
rect 141 707 175 723
rect 141 -785 175 -769
<< viali >>
rect -113 757 -45 791
rect 45 757 113 791
rect -175 -769 -141 707
rect -17 -769 17 707
rect 141 -769 175 707
<< metal1 >>
rect -125 791 -33 797
rect -125 757 -113 791
rect -45 757 -33 791
rect -125 751 -33 757
rect 33 791 125 797
rect 33 757 45 791
rect 113 757 125 791
rect 33 751 125 757
rect -181 707 -135 719
rect -181 -769 -175 707
rect -141 -769 -135 707
rect -181 -781 -135 -769
rect -23 707 23 719
rect -23 -769 -17 707
rect 17 -769 23 707
rect -23 -781 23 -769
rect 135 707 181 719
rect 135 -769 141 707
rect 175 -769 181 707
rect 135 -781 181 -769
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
