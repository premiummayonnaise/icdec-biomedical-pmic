magic
tech sky130A
magscale 1 2
timestamp 1769411983
<< error_p >>
rect -2559 1038 2559 1042
rect -2559 -970 -2529 1038
rect -2493 972 2493 976
rect -2493 -904 -2463 972
rect 2463 -904 2493 972
rect 2529 -970 2559 1038
<< nwell >>
rect -2529 -1004 2529 1038
<< mvpmos >>
rect -2435 -904 -2185 976
rect -2127 -904 -1877 976
rect -1819 -904 -1569 976
rect -1511 -904 -1261 976
rect -1203 -904 -953 976
rect -895 -904 -645 976
rect -587 -904 -337 976
rect -279 -904 -29 976
rect 29 -904 279 976
rect 337 -904 587 976
rect 645 -904 895 976
rect 953 -904 1203 976
rect 1261 -904 1511 976
rect 1569 -904 1819 976
rect 1877 -904 2127 976
rect 2185 -904 2435 976
<< mvpdiff >>
rect -2493 964 -2435 976
rect -2493 -892 -2481 964
rect -2447 -892 -2435 964
rect -2493 -904 -2435 -892
rect -2185 964 -2127 976
rect -2185 -892 -2173 964
rect -2139 -892 -2127 964
rect -2185 -904 -2127 -892
rect -1877 964 -1819 976
rect -1877 -892 -1865 964
rect -1831 -892 -1819 964
rect -1877 -904 -1819 -892
rect -1569 964 -1511 976
rect -1569 -892 -1557 964
rect -1523 -892 -1511 964
rect -1569 -904 -1511 -892
rect -1261 964 -1203 976
rect -1261 -892 -1249 964
rect -1215 -892 -1203 964
rect -1261 -904 -1203 -892
rect -953 964 -895 976
rect -953 -892 -941 964
rect -907 -892 -895 964
rect -953 -904 -895 -892
rect -645 964 -587 976
rect -645 -892 -633 964
rect -599 -892 -587 964
rect -645 -904 -587 -892
rect -337 964 -279 976
rect -337 -892 -325 964
rect -291 -892 -279 964
rect -337 -904 -279 -892
rect -29 964 29 976
rect -29 -892 -17 964
rect 17 -892 29 964
rect -29 -904 29 -892
rect 279 964 337 976
rect 279 -892 291 964
rect 325 -892 337 964
rect 279 -904 337 -892
rect 587 964 645 976
rect 587 -892 599 964
rect 633 -892 645 964
rect 587 -904 645 -892
rect 895 964 953 976
rect 895 -892 907 964
rect 941 -892 953 964
rect 895 -904 953 -892
rect 1203 964 1261 976
rect 1203 -892 1215 964
rect 1249 -892 1261 964
rect 1203 -904 1261 -892
rect 1511 964 1569 976
rect 1511 -892 1523 964
rect 1557 -892 1569 964
rect 1511 -904 1569 -892
rect 1819 964 1877 976
rect 1819 -892 1831 964
rect 1865 -892 1877 964
rect 1819 -904 1877 -892
rect 2127 964 2185 976
rect 2127 -892 2139 964
rect 2173 -892 2185 964
rect 2127 -904 2185 -892
rect 2435 964 2493 976
rect 2435 -892 2447 964
rect 2481 -892 2493 964
rect 2435 -904 2493 -892
<< mvpdiffc >>
rect -2481 -892 -2447 964
rect -2173 -892 -2139 964
rect -1865 -892 -1831 964
rect -1557 -892 -1523 964
rect -1249 -892 -1215 964
rect -941 -892 -907 964
rect -633 -892 -599 964
rect -325 -892 -291 964
rect -17 -892 17 964
rect 291 -892 325 964
rect 599 -892 633 964
rect 907 -892 941 964
rect 1215 -892 1249 964
rect 1523 -892 1557 964
rect 1831 -892 1865 964
rect 2139 -892 2173 964
rect 2447 -892 2481 964
<< poly >>
rect -2435 976 -2185 1002
rect -2127 976 -1877 1002
rect -1819 976 -1569 1002
rect -1511 976 -1261 1002
rect -1203 976 -953 1002
rect -895 976 -645 1002
rect -587 976 -337 1002
rect -279 976 -29 1002
rect 29 976 279 1002
rect 337 976 587 1002
rect 645 976 895 1002
rect 953 976 1203 1002
rect 1261 976 1511 1002
rect 1569 976 1819 1002
rect 1877 976 2127 1002
rect 2185 976 2435 1002
rect -2435 -951 -2185 -904
rect -2435 -985 -2419 -951
rect -2201 -985 -2185 -951
rect -2435 -1001 -2185 -985
rect -2127 -951 -1877 -904
rect -2127 -985 -2111 -951
rect -1893 -985 -1877 -951
rect -2127 -1001 -1877 -985
rect -1819 -951 -1569 -904
rect -1819 -985 -1803 -951
rect -1585 -985 -1569 -951
rect -1819 -1001 -1569 -985
rect -1511 -951 -1261 -904
rect -1511 -985 -1495 -951
rect -1277 -985 -1261 -951
rect -1511 -1001 -1261 -985
rect -1203 -951 -953 -904
rect -1203 -985 -1187 -951
rect -969 -985 -953 -951
rect -1203 -1001 -953 -985
rect -895 -951 -645 -904
rect -895 -985 -879 -951
rect -661 -985 -645 -951
rect -895 -1001 -645 -985
rect -587 -951 -337 -904
rect -587 -985 -571 -951
rect -353 -985 -337 -951
rect -587 -1001 -337 -985
rect -279 -951 -29 -904
rect -279 -985 -263 -951
rect -45 -985 -29 -951
rect -279 -1001 -29 -985
rect 29 -951 279 -904
rect 29 -985 45 -951
rect 263 -985 279 -951
rect 29 -1001 279 -985
rect 337 -951 587 -904
rect 337 -985 353 -951
rect 571 -985 587 -951
rect 337 -1001 587 -985
rect 645 -951 895 -904
rect 645 -985 661 -951
rect 879 -985 895 -951
rect 645 -1001 895 -985
rect 953 -951 1203 -904
rect 953 -985 969 -951
rect 1187 -985 1203 -951
rect 953 -1001 1203 -985
rect 1261 -951 1511 -904
rect 1261 -985 1277 -951
rect 1495 -985 1511 -951
rect 1261 -1001 1511 -985
rect 1569 -951 1819 -904
rect 1569 -985 1585 -951
rect 1803 -985 1819 -951
rect 1569 -1001 1819 -985
rect 1877 -951 2127 -904
rect 1877 -985 1893 -951
rect 2111 -985 2127 -951
rect 1877 -1001 2127 -985
rect 2185 -951 2435 -904
rect 2185 -985 2201 -951
rect 2419 -985 2435 -951
rect 2185 -1001 2435 -985
<< polycont >>
rect -2419 -985 -2201 -951
rect -2111 -985 -1893 -951
rect -1803 -985 -1585 -951
rect -1495 -985 -1277 -951
rect -1187 -985 -969 -951
rect -879 -985 -661 -951
rect -571 -985 -353 -951
rect -263 -985 -45 -951
rect 45 -985 263 -951
rect 353 -985 571 -951
rect 661 -985 879 -951
rect 969 -985 1187 -951
rect 1277 -985 1495 -951
rect 1585 -985 1803 -951
rect 1893 -985 2111 -951
rect 2201 -985 2419 -951
<< locali >>
rect -2481 964 -2447 980
rect -2481 -908 -2447 -892
rect -2173 964 -2139 980
rect -2173 -908 -2139 -892
rect -1865 964 -1831 980
rect -1865 -908 -1831 -892
rect -1557 964 -1523 980
rect -1557 -908 -1523 -892
rect -1249 964 -1215 980
rect -1249 -908 -1215 -892
rect -941 964 -907 980
rect -941 -908 -907 -892
rect -633 964 -599 980
rect -633 -908 -599 -892
rect -325 964 -291 980
rect -325 -908 -291 -892
rect -17 964 17 980
rect -17 -908 17 -892
rect 291 964 325 980
rect 291 -908 325 -892
rect 599 964 633 980
rect 599 -908 633 -892
rect 907 964 941 980
rect 907 -908 941 -892
rect 1215 964 1249 980
rect 1215 -908 1249 -892
rect 1523 964 1557 980
rect 1523 -908 1557 -892
rect 1831 964 1865 980
rect 1831 -908 1865 -892
rect 2139 964 2173 980
rect 2139 -908 2173 -892
rect 2447 964 2481 980
rect 2447 -908 2481 -892
rect -2435 -985 -2419 -951
rect -2201 -985 -2185 -951
rect -2127 -985 -2111 -951
rect -1893 -985 -1877 -951
rect -1819 -985 -1803 -951
rect -1585 -985 -1569 -951
rect -1511 -985 -1495 -951
rect -1277 -985 -1261 -951
rect -1203 -985 -1187 -951
rect -969 -985 -953 -951
rect -895 -985 -879 -951
rect -661 -985 -645 -951
rect -587 -985 -571 -951
rect -353 -985 -337 -951
rect -279 -985 -263 -951
rect -45 -985 -29 -951
rect 29 -985 45 -951
rect 263 -985 279 -951
rect 337 -985 353 -951
rect 571 -985 587 -951
rect 645 -985 661 -951
rect 879 -985 895 -951
rect 953 -985 969 -951
rect 1187 -985 1203 -951
rect 1261 -985 1277 -951
rect 1495 -985 1511 -951
rect 1569 -985 1585 -951
rect 1803 -985 1819 -951
rect 1877 -985 1893 -951
rect 2111 -985 2127 -951
rect 2185 -985 2201 -951
rect 2419 -985 2435 -951
<< viali >>
rect -2481 -892 -2447 964
rect -2173 -892 -2139 964
rect -1865 -892 -1831 964
rect -1557 -892 -1523 964
rect -1249 -892 -1215 964
rect -941 -892 -907 964
rect -633 -892 -599 964
rect -325 -892 -291 964
rect -17 -892 17 964
rect 291 -892 325 964
rect 599 -892 633 964
rect 907 -892 941 964
rect 1215 -892 1249 964
rect 1523 -892 1557 964
rect 1831 -892 1865 964
rect 2139 -892 2173 964
rect 2447 -892 2481 964
rect -2419 -985 -2201 -951
rect -2111 -985 -1893 -951
rect -1803 -985 -1585 -951
rect -1495 -985 -1277 -951
rect -1187 -985 -969 -951
rect -879 -985 -661 -951
rect -571 -985 -353 -951
rect -263 -985 -45 -951
rect 45 -985 263 -951
rect 353 -985 571 -951
rect 661 -985 879 -951
rect 969 -985 1187 -951
rect 1277 -985 1495 -951
rect 1585 -985 1803 -951
rect 1893 -985 2111 -951
rect 2201 -985 2419 -951
<< metal1 >>
rect -2487 964 -2441 976
rect -2487 -892 -2481 964
rect -2447 -892 -2441 964
rect -2487 -904 -2441 -892
rect -2179 964 -2133 976
rect -2179 -892 -2173 964
rect -2139 -892 -2133 964
rect -2179 -904 -2133 -892
rect -1871 964 -1825 976
rect -1871 -892 -1865 964
rect -1831 -892 -1825 964
rect -1871 -904 -1825 -892
rect -1563 964 -1517 976
rect -1563 -892 -1557 964
rect -1523 -892 -1517 964
rect -1563 -904 -1517 -892
rect -1255 964 -1209 976
rect -1255 -892 -1249 964
rect -1215 -892 -1209 964
rect -1255 -904 -1209 -892
rect -947 964 -901 976
rect -947 -892 -941 964
rect -907 -892 -901 964
rect -947 -904 -901 -892
rect -639 964 -593 976
rect -639 -892 -633 964
rect -599 -892 -593 964
rect -639 -904 -593 -892
rect -331 964 -285 976
rect -331 -892 -325 964
rect -291 -892 -285 964
rect -331 -904 -285 -892
rect -23 964 23 976
rect -23 -892 -17 964
rect 17 -892 23 964
rect -23 -904 23 -892
rect 285 964 331 976
rect 285 -892 291 964
rect 325 -892 331 964
rect 285 -904 331 -892
rect 593 964 639 976
rect 593 -892 599 964
rect 633 -892 639 964
rect 593 -904 639 -892
rect 901 964 947 976
rect 901 -892 907 964
rect 941 -892 947 964
rect 901 -904 947 -892
rect 1209 964 1255 976
rect 1209 -892 1215 964
rect 1249 -892 1255 964
rect 1209 -904 1255 -892
rect 1517 964 1563 976
rect 1517 -892 1523 964
rect 1557 -892 1563 964
rect 1517 -904 1563 -892
rect 1825 964 1871 976
rect 1825 -892 1831 964
rect 1865 -892 1871 964
rect 1825 -904 1871 -892
rect 2133 964 2179 976
rect 2133 -892 2139 964
rect 2173 -892 2179 964
rect 2133 -904 2179 -892
rect 2441 964 2487 976
rect 2441 -892 2447 964
rect 2481 -892 2487 964
rect 2441 -904 2487 -892
rect -2431 -951 -2189 -945
rect -2431 -985 -2419 -951
rect -2201 -985 -2189 -951
rect -2431 -991 -2189 -985
rect -2123 -951 -1881 -945
rect -2123 -985 -2111 -951
rect -1893 -985 -1881 -951
rect -2123 -991 -1881 -985
rect -1815 -951 -1573 -945
rect -1815 -985 -1803 -951
rect -1585 -985 -1573 -951
rect -1815 -991 -1573 -985
rect -1507 -951 -1265 -945
rect -1507 -985 -1495 -951
rect -1277 -985 -1265 -951
rect -1507 -991 -1265 -985
rect -1199 -951 -957 -945
rect -1199 -985 -1187 -951
rect -969 -985 -957 -951
rect -1199 -991 -957 -985
rect -891 -951 -649 -945
rect -891 -985 -879 -951
rect -661 -985 -649 -951
rect -891 -991 -649 -985
rect -583 -951 -341 -945
rect -583 -985 -571 -951
rect -353 -985 -341 -951
rect -583 -991 -341 -985
rect -275 -951 -33 -945
rect -275 -985 -263 -951
rect -45 -985 -33 -951
rect -275 -991 -33 -985
rect 33 -951 275 -945
rect 33 -985 45 -951
rect 263 -985 275 -951
rect 33 -991 275 -985
rect 341 -951 583 -945
rect 341 -985 353 -951
rect 571 -985 583 -951
rect 341 -991 583 -985
rect 649 -951 891 -945
rect 649 -985 661 -951
rect 879 -985 891 -951
rect 649 -991 891 -985
rect 957 -951 1199 -945
rect 957 -985 969 -951
rect 1187 -985 1199 -951
rect 957 -991 1199 -985
rect 1265 -951 1507 -945
rect 1265 -985 1277 -951
rect 1495 -985 1507 -951
rect 1265 -991 1507 -985
rect 1573 -951 1815 -945
rect 1573 -985 1585 -951
rect 1803 -985 1815 -951
rect 1573 -991 1815 -985
rect 1881 -951 2123 -945
rect 1881 -985 1893 -951
rect 2111 -985 2123 -951
rect 1881 -991 2123 -985
rect 2189 -951 2431 -945
rect 2189 -985 2201 -951
rect 2419 -985 2431 -951
rect 2189 -991 2431 -985
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9.4 l 1.25 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
