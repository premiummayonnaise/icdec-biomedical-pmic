magic
tech sky130A
magscale 1 2
timestamp 1770083437
<< nwell >>
rect 1200 2100 9200 5200
rect 1200 -4200 1800 2100
rect 8600 -4200 9200 2100
rect 1200 -4600 9200 -4200
<< pwell >>
rect 1800 -4200 8600 2000
<< psubdiff >>
rect 2400 -2200 2500 -1800
rect 7900 -2200 8000 -1800
<< nsubdiff >>
rect 1300 5060 9100 5100
rect 1300 4940 1500 5060
rect 2060 4940 8340 5060
rect 8900 4940 9100 5060
rect 1300 4900 9100 4940
rect 1300 4880 1500 4900
rect 1300 -4280 1340 4880
rect 1460 -4280 1500 4880
rect 2080 4760 8280 4900
rect 8900 4880 9100 4900
rect 1300 -4300 1500 -4280
rect 8900 -4280 8940 4880
rect 9060 -4280 9100 4880
rect 8900 -4300 9100 -4280
rect 1300 -4340 9100 -4300
rect 1300 -4460 1520 -4340
rect 8880 -4460 9100 -4340
rect 1300 -4500 9100 -4460
<< nsubdiffcont >>
rect 1500 4940 2060 5060
rect 8340 4940 8900 5060
rect 1340 -4280 1460 4880
rect 8940 -4280 9060 4880
rect 1520 -4460 8880 -4340
<< locali >>
rect 1300 5060 9100 5100
rect 1300 4940 1500 5060
rect 2060 5000 2100 5060
rect 2160 5000 2200 5060
rect 2260 5000 2300 5060
rect 2360 5000 2400 5060
rect 2460 5000 2500 5060
rect 2560 5000 2600 5060
rect 2660 5000 2700 5060
rect 2760 5000 2800 5060
rect 2860 5000 2900 5060
rect 2960 5000 3000 5060
rect 3060 5000 3100 5060
rect 3160 5000 3200 5060
rect 3260 5000 3300 5060
rect 3360 5000 3400 5060
rect 3460 5000 3500 5060
rect 3560 5000 3600 5060
rect 3660 5000 3700 5060
rect 3760 5000 3800 5060
rect 3860 5000 3900 5060
rect 3960 5000 4000 5060
rect 4060 5000 4100 5060
rect 4160 5000 4200 5060
rect 4260 5000 4300 5060
rect 4360 5000 4400 5060
rect 4460 5000 4500 5060
rect 4560 5000 4600 5060
rect 4660 5000 4700 5060
rect 4760 5000 4800 5060
rect 4860 5000 4900 5060
rect 4960 5000 5000 5060
rect 5060 5000 5100 5060
rect 5160 5000 5200 5060
rect 5260 5000 5300 5060
rect 5360 5000 5400 5060
rect 5460 5000 5500 5060
rect 5560 5000 5600 5060
rect 5660 5000 5700 5060
rect 5760 5000 5800 5060
rect 5860 5000 5900 5060
rect 5960 5000 6000 5060
rect 6060 5000 6100 5060
rect 6160 5000 6200 5060
rect 6260 5000 6300 5060
rect 6360 5000 6400 5060
rect 6460 5000 6500 5060
rect 6560 5000 6600 5060
rect 6660 5000 6700 5060
rect 6760 5000 6800 5060
rect 6860 5000 6900 5060
rect 6960 5000 7000 5060
rect 7060 5000 7100 5060
rect 7160 5000 7200 5060
rect 7260 5000 7300 5060
rect 7360 5000 7400 5060
rect 7460 5000 7500 5060
rect 7560 5000 7600 5060
rect 7660 5000 7700 5060
rect 7760 5000 7800 5060
rect 7860 5000 7900 5060
rect 7960 5000 8000 5060
rect 8060 5000 8100 5060
rect 8160 5000 8200 5060
rect 8260 5000 8340 5060
rect 2060 4960 8340 5000
rect 2060 4940 2100 4960
rect 1300 4900 2100 4940
rect 2160 4900 2200 4960
rect 2260 4900 2300 4960
rect 2360 4900 2400 4960
rect 2460 4900 2500 4960
rect 2560 4900 2600 4960
rect 2660 4900 2700 4960
rect 2760 4900 2800 4960
rect 2860 4900 2900 4960
rect 2960 4900 3000 4960
rect 3060 4900 3100 4960
rect 3160 4900 3200 4960
rect 3260 4900 3300 4960
rect 3360 4900 3400 4960
rect 3460 4900 3500 4960
rect 3560 4900 3600 4960
rect 3660 4900 3700 4960
rect 3760 4900 3800 4960
rect 3860 4900 3900 4960
rect 3960 4900 4000 4960
rect 4060 4900 4100 4960
rect 4160 4900 4200 4960
rect 4260 4900 4300 4960
rect 4360 4900 4400 4960
rect 4460 4900 4500 4960
rect 4560 4900 4600 4960
rect 4660 4900 4700 4960
rect 4760 4900 4800 4960
rect 4860 4900 4900 4960
rect 4960 4900 5000 4960
rect 5060 4900 5100 4960
rect 5160 4900 5200 4960
rect 5260 4900 5300 4960
rect 5360 4900 5400 4960
rect 5460 4900 5500 4960
rect 5560 4900 5600 4960
rect 5660 4900 5700 4960
rect 5760 4900 5800 4960
rect 5860 4900 5900 4960
rect 5960 4900 6000 4960
rect 6060 4900 6100 4960
rect 6160 4900 6200 4960
rect 6260 4900 6300 4960
rect 6360 4900 6400 4960
rect 6460 4900 6500 4960
rect 6560 4900 6600 4960
rect 6660 4900 6700 4960
rect 6760 4900 6800 4960
rect 6860 4900 6900 4960
rect 6960 4900 7000 4960
rect 7060 4900 7100 4960
rect 7160 4900 7200 4960
rect 7260 4900 7300 4960
rect 7360 4900 7400 4960
rect 7460 4900 7500 4960
rect 7560 4900 7600 4960
rect 7660 4900 7700 4960
rect 7760 4900 7800 4960
rect 7860 4900 7900 4960
rect 7960 4900 8000 4960
rect 8060 4900 8100 4960
rect 8160 4900 8200 4960
rect 8260 4940 8340 4960
rect 8900 4940 9100 5060
rect 8260 4900 9100 4940
rect 1300 4880 9100 4900
rect 1300 -4280 1340 4880
rect 1460 4860 8940 4880
rect 1460 4800 2100 4860
rect 2160 4800 2200 4860
rect 2260 4800 2300 4860
rect 2360 4800 2400 4860
rect 2460 4800 2500 4860
rect 2560 4800 2600 4860
rect 2660 4800 2700 4860
rect 2760 4800 2800 4860
rect 2860 4800 2900 4860
rect 2960 4800 3000 4860
rect 3060 4800 3100 4860
rect 3160 4800 3200 4860
rect 3260 4800 3300 4860
rect 3360 4800 3400 4860
rect 3460 4800 3500 4860
rect 3560 4800 3600 4860
rect 3660 4800 3700 4860
rect 3760 4800 3800 4860
rect 3860 4800 3900 4860
rect 3960 4800 4000 4860
rect 4060 4800 4100 4860
rect 4160 4800 4200 4860
rect 4260 4800 4300 4860
rect 4360 4800 4400 4860
rect 4460 4800 4500 4860
rect 4560 4800 4600 4860
rect 4660 4800 4700 4860
rect 4760 4800 4800 4860
rect 4860 4800 4900 4860
rect 4960 4800 5000 4860
rect 5060 4800 5100 4860
rect 5160 4800 5200 4860
rect 5260 4800 5300 4860
rect 5360 4800 5400 4860
rect 5460 4800 5500 4860
rect 5560 4800 5600 4860
rect 5660 4800 5700 4860
rect 5760 4800 5800 4860
rect 5860 4800 5900 4860
rect 5960 4800 6000 4860
rect 6060 4800 6100 4860
rect 6160 4800 6200 4860
rect 6260 4800 6300 4860
rect 6360 4800 6400 4860
rect 6460 4800 6500 4860
rect 6560 4800 6600 4860
rect 6660 4800 6700 4860
rect 6760 4800 6800 4860
rect 6860 4800 6900 4860
rect 6960 4800 7000 4860
rect 7060 4800 7100 4860
rect 7160 4800 7200 4860
rect 7260 4800 7300 4860
rect 7360 4800 7400 4860
rect 7460 4800 7500 4860
rect 7560 4800 7600 4860
rect 7660 4800 7700 4860
rect 7760 4800 7800 4860
rect 7860 4800 7900 4860
rect 7960 4800 8000 4860
rect 8060 4800 8100 4860
rect 8160 4800 8200 4860
rect 8260 4800 8940 4860
rect 1460 4760 8940 4800
rect 1460 2496 2176 4760
rect 8216 2496 8940 4760
rect 1460 2380 8940 2496
rect 1460 2098 4800 2380
rect 5000 2100 5400 2300
rect 5600 2100 8940 2380
rect 1460 -4280 1500 2098
rect 1560 -1800 2400 2000
rect 8000 -1800 8840 2000
rect 1560 -1860 4920 -1800
rect 1560 -1940 2540 -1860
rect 2620 -1940 2660 -1860
rect 2740 -1940 2780 -1860
rect 2860 -1940 2900 -1860
rect 2980 -1940 3020 -1860
rect 3100 -1940 3140 -1860
rect 3220 -1940 3260 -1860
rect 3340 -1940 3380 -1860
rect 3460 -1940 3500 -1860
rect 3580 -1940 3620 -1860
rect 3700 -1940 3740 -1860
rect 3820 -1940 3860 -1860
rect 3940 -1940 3980 -1860
rect 4060 -1940 4100 -1860
rect 4180 -1940 4220 -1860
rect 4300 -1940 4340 -1860
rect 4420 -1940 4460 -1860
rect 4540 -1940 4580 -1860
rect 4660 -1940 4700 -1860
rect 4780 -1940 4820 -1860
rect 4900 -1940 4920 -1860
rect 1560 -1980 4920 -1940
rect 1560 -2060 2420 -1980
rect 2500 -2060 2540 -1980
rect 2620 -2060 2660 -1980
rect 2740 -2060 2780 -1980
rect 2860 -2060 2900 -1980
rect 2980 -2060 3020 -1980
rect 3100 -2060 3140 -1980
rect 3220 -2060 3260 -1980
rect 3340 -2060 3380 -1980
rect 3460 -2060 3500 -1980
rect 3580 -2060 3620 -1980
rect 3700 -2060 3740 -1980
rect 3820 -2060 3860 -1980
rect 3940 -2060 3980 -1980
rect 4060 -2060 4100 -1980
rect 4180 -2060 4220 -1980
rect 4300 -2060 4340 -1980
rect 4420 -2060 4460 -1980
rect 4540 -2060 4580 -1980
rect 4660 -2060 4700 -1980
rect 4780 -2060 4820 -1980
rect 4900 -2060 4920 -1980
rect 1560 -2100 4920 -2060
rect 1560 -2140 2420 -2100
rect 1560 -4100 2225 -2140
rect 2400 -2180 2420 -2140
rect 2500 -2180 2540 -2100
rect 2620 -2180 2660 -2100
rect 2740 -2180 2780 -2100
rect 2860 -2180 2900 -2100
rect 2980 -2180 3020 -2100
rect 3100 -2180 3140 -2100
rect 3220 -2180 3260 -2100
rect 3340 -2180 3380 -2100
rect 3460 -2180 3500 -2100
rect 3580 -2180 3620 -2100
rect 3700 -2180 3740 -2100
rect 3820 -2180 3860 -2100
rect 3940 -2180 3980 -2100
rect 4060 -2180 4100 -2100
rect 4180 -2180 4220 -2100
rect 4300 -2180 4340 -2100
rect 4420 -2180 4460 -2100
rect 4540 -2180 4580 -2100
rect 4660 -2180 4700 -2100
rect 4780 -2180 4820 -2100
rect 4900 -2180 4920 -2100
rect 2400 -2200 4920 -2180
rect 5480 -1860 8840 -1800
rect 5480 -1940 5500 -1860
rect 5580 -1940 5620 -1860
rect 5700 -1940 5740 -1860
rect 5820 -1940 5860 -1860
rect 5940 -1940 5980 -1860
rect 6060 -1940 6100 -1860
rect 6180 -1940 6220 -1860
rect 6300 -1940 6340 -1860
rect 6420 -1940 6460 -1860
rect 6540 -1940 6580 -1860
rect 6660 -1940 6700 -1860
rect 6780 -1940 6820 -1860
rect 6900 -1940 6940 -1860
rect 7020 -1940 7060 -1860
rect 7140 -1940 7180 -1860
rect 7260 -1940 7300 -1860
rect 7380 -1940 7420 -1860
rect 7500 -1940 7540 -1860
rect 7620 -1940 7660 -1860
rect 7740 -1940 7780 -1860
rect 7860 -1940 7900 -1860
rect 7980 -1940 8840 -1860
rect 5480 -1980 8840 -1940
rect 5480 -2060 5500 -1980
rect 5580 -2060 5620 -1980
rect 5700 -2060 5740 -1980
rect 5820 -2060 5860 -1980
rect 5940 -2060 5980 -1980
rect 6060 -2060 6100 -1980
rect 6180 -2060 6220 -1980
rect 6300 -2060 6340 -1980
rect 6420 -2060 6460 -1980
rect 6540 -2060 6580 -1980
rect 6660 -2060 6700 -1980
rect 6780 -2060 6820 -1980
rect 6900 -2060 6940 -1980
rect 7020 -2060 7060 -1980
rect 7140 -2060 7180 -1980
rect 7260 -2060 7300 -1980
rect 7380 -2060 7420 -1980
rect 7500 -2060 7540 -1980
rect 7620 -2060 7660 -1980
rect 7740 -2060 7780 -1980
rect 7860 -2060 7900 -1980
rect 7980 -2060 8840 -1980
rect 5480 -2100 8840 -2060
rect 5480 -2180 5500 -2100
rect 5580 -2180 5620 -2100
rect 5700 -2180 5740 -2100
rect 5820 -2180 5860 -2100
rect 5940 -2180 5980 -2100
rect 6060 -2180 6100 -2100
rect 6180 -2180 6220 -2100
rect 6300 -2180 6340 -2100
rect 6420 -2180 6460 -2100
rect 6540 -2180 6580 -2100
rect 6660 -2180 6700 -2100
rect 6780 -2180 6820 -2100
rect 6900 -2180 6940 -2100
rect 7020 -2180 7060 -2100
rect 7140 -2180 7180 -2100
rect 7260 -2180 7300 -2100
rect 7380 -2180 7420 -2100
rect 7500 -2180 7540 -2100
rect 7620 -2180 7660 -2100
rect 7740 -2180 7780 -2100
rect 7860 -2180 7900 -2100
rect 7980 -2160 8840 -2100
rect 7980 -2180 8000 -2160
rect 5480 -2200 8000 -2180
rect 8200 -4100 8840 -2160
rect 1560 -4260 8840 -4100
rect 1300 -4300 1500 -4280
rect 8900 -4280 8940 2100
rect 9060 -4280 9100 4880
rect 8900 -4300 9100 -4280
rect 1300 -4340 9100 -4300
rect 1300 -4460 1520 -4340
rect 8880 -4460 9100 -4340
rect 1300 -4500 9100 -4460
<< viali >>
rect 2100 5000 2160 5060
rect 2200 5000 2260 5060
rect 2300 5000 2360 5060
rect 2400 5000 2460 5060
rect 2500 5000 2560 5060
rect 2600 5000 2660 5060
rect 2700 5000 2760 5060
rect 2800 5000 2860 5060
rect 2900 5000 2960 5060
rect 3000 5000 3060 5060
rect 3100 5000 3160 5060
rect 3200 5000 3260 5060
rect 3300 5000 3360 5060
rect 3400 5000 3460 5060
rect 3500 5000 3560 5060
rect 3600 5000 3660 5060
rect 3700 5000 3760 5060
rect 3800 5000 3860 5060
rect 3900 5000 3960 5060
rect 4000 5000 4060 5060
rect 4100 5000 4160 5060
rect 4200 5000 4260 5060
rect 4300 5000 4360 5060
rect 4400 5000 4460 5060
rect 4500 5000 4560 5060
rect 4600 5000 4660 5060
rect 4700 5000 4760 5060
rect 4800 5000 4860 5060
rect 4900 5000 4960 5060
rect 5000 5000 5060 5060
rect 5100 5000 5160 5060
rect 5200 5000 5260 5060
rect 5300 5000 5360 5060
rect 5400 5000 5460 5060
rect 5500 5000 5560 5060
rect 5600 5000 5660 5060
rect 5700 5000 5760 5060
rect 5800 5000 5860 5060
rect 5900 5000 5960 5060
rect 6000 5000 6060 5060
rect 6100 5000 6160 5060
rect 6200 5000 6260 5060
rect 6300 5000 6360 5060
rect 6400 5000 6460 5060
rect 6500 5000 6560 5060
rect 6600 5000 6660 5060
rect 6700 5000 6760 5060
rect 6800 5000 6860 5060
rect 6900 5000 6960 5060
rect 7000 5000 7060 5060
rect 7100 5000 7160 5060
rect 7200 5000 7260 5060
rect 7300 5000 7360 5060
rect 7400 5000 7460 5060
rect 7500 5000 7560 5060
rect 7600 5000 7660 5060
rect 7700 5000 7760 5060
rect 7800 5000 7860 5060
rect 7900 5000 7960 5060
rect 8000 5000 8060 5060
rect 8100 5000 8160 5060
rect 8200 5000 8260 5060
rect 2100 4900 2160 4960
rect 2200 4900 2260 4960
rect 2300 4900 2360 4960
rect 2400 4900 2460 4960
rect 2500 4900 2560 4960
rect 2600 4900 2660 4960
rect 2700 4900 2760 4960
rect 2800 4900 2860 4960
rect 2900 4900 2960 4960
rect 3000 4900 3060 4960
rect 3100 4900 3160 4960
rect 3200 4900 3260 4960
rect 3300 4900 3360 4960
rect 3400 4900 3460 4960
rect 3500 4900 3560 4960
rect 3600 4900 3660 4960
rect 3700 4900 3760 4960
rect 3800 4900 3860 4960
rect 3900 4900 3960 4960
rect 4000 4900 4060 4960
rect 4100 4900 4160 4960
rect 4200 4900 4260 4960
rect 4300 4900 4360 4960
rect 4400 4900 4460 4960
rect 4500 4900 4560 4960
rect 4600 4900 4660 4960
rect 4700 4900 4760 4960
rect 4800 4900 4860 4960
rect 4900 4900 4960 4960
rect 5000 4900 5060 4960
rect 5100 4900 5160 4960
rect 5200 4900 5260 4960
rect 5300 4900 5360 4960
rect 5400 4900 5460 4960
rect 5500 4900 5560 4960
rect 5600 4900 5660 4960
rect 5700 4900 5760 4960
rect 5800 4900 5860 4960
rect 5900 4900 5960 4960
rect 6000 4900 6060 4960
rect 6100 4900 6160 4960
rect 6200 4900 6260 4960
rect 6300 4900 6360 4960
rect 6400 4900 6460 4960
rect 6500 4900 6560 4960
rect 6600 4900 6660 4960
rect 6700 4900 6760 4960
rect 6800 4900 6860 4960
rect 6900 4900 6960 4960
rect 7000 4900 7060 4960
rect 7100 4900 7160 4960
rect 7200 4900 7260 4960
rect 7300 4900 7360 4960
rect 7400 4900 7460 4960
rect 7500 4900 7560 4960
rect 7600 4900 7660 4960
rect 7700 4900 7760 4960
rect 7800 4900 7860 4960
rect 7900 4900 7960 4960
rect 8000 4900 8060 4960
rect 8100 4900 8160 4960
rect 8200 4900 8260 4960
rect 2100 4800 2160 4860
rect 2200 4800 2260 4860
rect 2300 4800 2360 4860
rect 2400 4800 2460 4860
rect 2500 4800 2560 4860
rect 2600 4800 2660 4860
rect 2700 4800 2760 4860
rect 2800 4800 2860 4860
rect 2900 4800 2960 4860
rect 3000 4800 3060 4860
rect 3100 4800 3160 4860
rect 3200 4800 3260 4860
rect 3300 4800 3360 4860
rect 3400 4800 3460 4860
rect 3500 4800 3560 4860
rect 3600 4800 3660 4860
rect 3700 4800 3760 4860
rect 3800 4800 3860 4860
rect 3900 4800 3960 4860
rect 4000 4800 4060 4860
rect 4100 4800 4160 4860
rect 4200 4800 4260 4860
rect 4300 4800 4360 4860
rect 4400 4800 4460 4860
rect 4500 4800 4560 4860
rect 4600 4800 4660 4860
rect 4700 4800 4760 4860
rect 4800 4800 4860 4860
rect 4900 4800 4960 4860
rect 5000 4800 5060 4860
rect 5100 4800 5160 4860
rect 5200 4800 5260 4860
rect 5300 4800 5360 4860
rect 5400 4800 5460 4860
rect 5500 4800 5560 4860
rect 5600 4800 5660 4860
rect 5700 4800 5760 4860
rect 5800 4800 5860 4860
rect 5900 4800 5960 4860
rect 6000 4800 6060 4860
rect 6100 4800 6160 4860
rect 6200 4800 6260 4860
rect 6300 4800 6360 4860
rect 6400 4800 6460 4860
rect 6500 4800 6560 4860
rect 6600 4800 6660 4860
rect 6700 4800 6760 4860
rect 6800 4800 6860 4860
rect 6900 4800 6960 4860
rect 7000 4800 7060 4860
rect 7100 4800 7160 4860
rect 7200 4800 7260 4860
rect 7300 4800 7360 4860
rect 7400 4800 7460 4860
rect 7500 4800 7560 4860
rect 7600 4800 7660 4860
rect 7700 4800 7760 4860
rect 7800 4800 7860 4860
rect 7900 4800 7960 4860
rect 8000 4800 8060 4860
rect 8100 4800 8160 4860
rect 8200 4800 8260 4860
rect 2540 -1940 2620 -1860
rect 2660 -1940 2740 -1860
rect 2780 -1940 2860 -1860
rect 2900 -1940 2980 -1860
rect 3020 -1940 3100 -1860
rect 3140 -1940 3220 -1860
rect 3260 -1940 3340 -1860
rect 3380 -1940 3460 -1860
rect 3500 -1940 3580 -1860
rect 3620 -1940 3700 -1860
rect 3740 -1940 3820 -1860
rect 3860 -1940 3940 -1860
rect 3980 -1940 4060 -1860
rect 4100 -1940 4180 -1860
rect 4220 -1940 4300 -1860
rect 4340 -1940 4420 -1860
rect 4460 -1940 4540 -1860
rect 4580 -1940 4660 -1860
rect 4700 -1940 4780 -1860
rect 4820 -1940 4900 -1860
rect 2420 -2060 2500 -1980
rect 2540 -2060 2620 -1980
rect 2660 -2060 2740 -1980
rect 2780 -2060 2860 -1980
rect 2900 -2060 2980 -1980
rect 3020 -2060 3100 -1980
rect 3140 -2060 3220 -1980
rect 3260 -2060 3340 -1980
rect 3380 -2060 3460 -1980
rect 3500 -2060 3580 -1980
rect 3620 -2060 3700 -1980
rect 3740 -2060 3820 -1980
rect 3860 -2060 3940 -1980
rect 3980 -2060 4060 -1980
rect 4100 -2060 4180 -1980
rect 4220 -2060 4300 -1980
rect 4340 -2060 4420 -1980
rect 4460 -2060 4540 -1980
rect 4580 -2060 4660 -1980
rect 4700 -2060 4780 -1980
rect 4820 -2060 4900 -1980
rect 2420 -2180 2500 -2100
rect 2540 -2180 2620 -2100
rect 2660 -2180 2740 -2100
rect 2780 -2180 2860 -2100
rect 2900 -2180 2980 -2100
rect 3020 -2180 3100 -2100
rect 3140 -2180 3220 -2100
rect 3260 -2180 3340 -2100
rect 3380 -2180 3460 -2100
rect 3500 -2180 3580 -2100
rect 3620 -2180 3700 -2100
rect 3740 -2180 3820 -2100
rect 3860 -2180 3940 -2100
rect 3980 -2180 4060 -2100
rect 4100 -2180 4180 -2100
rect 4220 -2180 4300 -2100
rect 4340 -2180 4420 -2100
rect 4460 -2180 4540 -2100
rect 4580 -2180 4660 -2100
rect 4700 -2180 4780 -2100
rect 4820 -2180 4900 -2100
rect 5500 -1940 5580 -1860
rect 5620 -1940 5700 -1860
rect 5740 -1940 5820 -1860
rect 5860 -1940 5940 -1860
rect 5980 -1940 6060 -1860
rect 6100 -1940 6180 -1860
rect 6220 -1940 6300 -1860
rect 6340 -1940 6420 -1860
rect 6460 -1940 6540 -1860
rect 6580 -1940 6660 -1860
rect 6700 -1940 6780 -1860
rect 6820 -1940 6900 -1860
rect 6940 -1940 7020 -1860
rect 7060 -1940 7140 -1860
rect 7180 -1940 7260 -1860
rect 7300 -1940 7380 -1860
rect 7420 -1940 7500 -1860
rect 7540 -1940 7620 -1860
rect 7660 -1940 7740 -1860
rect 7780 -1940 7860 -1860
rect 7900 -1940 7980 -1860
rect 5500 -2060 5580 -1980
rect 5620 -2060 5700 -1980
rect 5740 -2060 5820 -1980
rect 5860 -2060 5940 -1980
rect 5980 -2060 6060 -1980
rect 6100 -2060 6180 -1980
rect 6220 -2060 6300 -1980
rect 6340 -2060 6420 -1980
rect 6460 -2060 6540 -1980
rect 6580 -2060 6660 -1980
rect 6700 -2060 6780 -1980
rect 6820 -2060 6900 -1980
rect 6940 -2060 7020 -1980
rect 7060 -2060 7140 -1980
rect 7180 -2060 7260 -1980
rect 7300 -2060 7380 -1980
rect 7420 -2060 7500 -1980
rect 7540 -2060 7620 -1980
rect 7660 -2060 7740 -1980
rect 7780 -2060 7860 -1980
rect 7900 -2060 7980 -1980
rect 5500 -2180 5580 -2100
rect 5620 -2180 5700 -2100
rect 5740 -2180 5820 -2100
rect 5860 -2180 5940 -2100
rect 5980 -2180 6060 -2100
rect 6100 -2180 6180 -2100
rect 6220 -2180 6300 -2100
rect 6340 -2180 6420 -2100
rect 6460 -2180 6540 -2100
rect 6580 -2180 6660 -2100
rect 6700 -2180 6780 -2100
rect 6820 -2180 6900 -2100
rect 6940 -2180 7020 -2100
rect 7060 -2180 7140 -2100
rect 7180 -2180 7260 -2100
rect 7300 -2180 7380 -2100
rect 7420 -2180 7500 -2100
rect 7540 -2180 7620 -2100
rect 7660 -2180 7740 -2100
rect 7780 -2180 7860 -2100
rect 7900 -2180 7980 -2100
<< metal1 >>
rect 2080 5060 8280 5100
rect 2080 5000 2100 5060
rect 2160 5000 2200 5060
rect 2260 5000 2300 5060
rect 2360 5000 2400 5060
rect 2460 5000 2500 5060
rect 2560 5000 2600 5060
rect 2660 5000 2700 5060
rect 2760 5000 2800 5060
rect 2860 5000 2900 5060
rect 2960 5000 3000 5060
rect 3060 5000 3100 5060
rect 3160 5000 3200 5060
rect 3260 5000 3300 5060
rect 3360 5000 3400 5060
rect 3460 5000 3500 5060
rect 3560 5000 3600 5060
rect 3660 5000 3700 5060
rect 3760 5000 3800 5060
rect 3860 5000 3900 5060
rect 3960 5000 4000 5060
rect 4060 5000 4100 5060
rect 4160 5000 4200 5060
rect 4260 5000 4300 5060
rect 4360 5000 4400 5060
rect 4460 5000 4500 5060
rect 4560 5000 4600 5060
rect 4660 5000 4700 5060
rect 4760 5000 4800 5060
rect 4860 5000 4900 5060
rect 4960 5000 5000 5060
rect 5060 5000 5100 5060
rect 5160 5000 5200 5060
rect 5260 5000 5300 5060
rect 5360 5000 5400 5060
rect 5460 5000 5500 5060
rect 5560 5000 5600 5060
rect 5660 5000 5700 5060
rect 5760 5000 5800 5060
rect 5860 5000 5900 5060
rect 5960 5000 6000 5060
rect 6060 5000 6100 5060
rect 6160 5000 6200 5060
rect 6260 5000 6300 5060
rect 6360 5000 6400 5060
rect 6460 5000 6500 5060
rect 6560 5000 6600 5060
rect 6660 5000 6700 5060
rect 6760 5000 6800 5060
rect 6860 5000 6900 5060
rect 6960 5000 7000 5060
rect 7060 5000 7100 5060
rect 7160 5000 7200 5060
rect 7260 5000 7300 5060
rect 7360 5000 7400 5060
rect 7460 5000 7500 5060
rect 7560 5000 7600 5060
rect 7660 5000 7700 5060
rect 7760 5000 7800 5060
rect 7860 5000 7900 5060
rect 7960 5000 8000 5060
rect 8060 5000 8100 5060
rect 8160 5000 8200 5060
rect 8260 5000 8280 5060
rect 2080 4960 8280 5000
rect 2080 4900 2100 4960
rect 2160 4900 2200 4960
rect 2260 4900 2300 4960
rect 2360 4900 2400 4960
rect 2460 4900 2500 4960
rect 2560 4900 2600 4960
rect 2660 4900 2700 4960
rect 2760 4900 2800 4960
rect 2860 4900 2900 4960
rect 2960 4900 3000 4960
rect 3060 4900 3100 4960
rect 3160 4900 3200 4960
rect 3260 4900 3300 4960
rect 3360 4900 3400 4960
rect 3460 4900 3500 4960
rect 3560 4900 3600 4960
rect 3660 4900 3700 4960
rect 3760 4900 3800 4960
rect 3860 4900 3900 4960
rect 3960 4900 4000 4960
rect 4060 4900 4100 4960
rect 4160 4900 4200 4960
rect 4260 4900 4300 4960
rect 4360 4900 4400 4960
rect 4460 4900 4500 4960
rect 4560 4900 4600 4960
rect 4660 4900 4700 4960
rect 4760 4900 4800 4960
rect 4860 4900 4900 4960
rect 4960 4900 5000 4960
rect 5060 4900 5100 4960
rect 5160 4900 5200 4960
rect 5260 4900 5300 4960
rect 5360 4900 5400 4960
rect 5460 4900 5500 4960
rect 5560 4900 5600 4960
rect 5660 4900 5700 4960
rect 5760 4900 5800 4960
rect 5860 4900 5900 4960
rect 5960 4900 6000 4960
rect 6060 4900 6100 4960
rect 6160 4900 6200 4960
rect 6260 4900 6300 4960
rect 6360 4900 6400 4960
rect 6460 4900 6500 4960
rect 6560 4900 6600 4960
rect 6660 4900 6700 4960
rect 6760 4900 6800 4960
rect 6860 4900 6900 4960
rect 6960 4900 7000 4960
rect 7060 4900 7100 4960
rect 7160 4900 7200 4960
rect 7260 4900 7300 4960
rect 7360 4900 7400 4960
rect 7460 4900 7500 4960
rect 7560 4900 7600 4960
rect 7660 4900 7700 4960
rect 7760 4900 7800 4960
rect 7860 4900 7900 4960
rect 7960 4900 8000 4960
rect 8060 4900 8100 4960
rect 8160 4900 8200 4960
rect 8260 4900 8280 4960
rect 2080 4860 8280 4900
rect 2080 4800 2100 4860
rect 2160 4800 2200 4860
rect 2260 4800 2300 4860
rect 2360 4800 2400 4860
rect 2460 4800 2500 4860
rect 2560 4800 2600 4860
rect 2660 4800 2700 4860
rect 2760 4800 2800 4860
rect 2860 4800 2900 4860
rect 2960 4800 3000 4860
rect 3060 4800 3100 4860
rect 3160 4800 3200 4860
rect 3260 4800 3300 4860
rect 3360 4800 3400 4860
rect 3460 4800 3500 4860
rect 3560 4800 3600 4860
rect 3660 4800 3700 4860
rect 3760 4800 3800 4860
rect 3860 4800 3900 4860
rect 3960 4800 4000 4860
rect 4060 4800 4100 4860
rect 4160 4800 4200 4860
rect 4260 4800 4300 4860
rect 4360 4800 4400 4860
rect 4460 4800 4500 4860
rect 4560 4800 4600 4860
rect 4660 4800 4700 4860
rect 4760 4800 4800 4860
rect 4860 4800 4900 4860
rect 4960 4800 5000 4860
rect 5060 4800 5100 4860
rect 5160 4800 5200 4860
rect 5260 4800 5300 4860
rect 5360 4800 5400 4860
rect 5460 4800 5500 4860
rect 5560 4800 5600 4860
rect 5660 4800 5700 4860
rect 5760 4800 5800 4860
rect 5860 4800 5900 4860
rect 5960 4800 6000 4860
rect 6060 4800 6100 4860
rect 6160 4800 6200 4860
rect 6260 4800 6300 4860
rect 6360 4800 6400 4860
rect 6460 4800 6500 4860
rect 6560 4800 6600 4860
rect 6660 4800 6700 4860
rect 6760 4800 6800 4860
rect 6860 4800 6900 4860
rect 6960 4800 7000 4860
rect 7060 4800 7100 4860
rect 7160 4800 7200 4860
rect 7260 4800 7300 4860
rect 7360 4800 7400 4860
rect 7460 4800 7500 4860
rect 7560 4800 7600 4860
rect 7660 4800 7700 4860
rect 7760 4800 7800 4860
rect 7860 4800 7900 4860
rect 7960 4800 8000 4860
rect 8060 4800 8100 4860
rect 8160 4800 8200 4860
rect 8260 4800 8280 4860
rect 2080 4760 8280 4800
rect 5000 2280 5400 2300
rect 5000 2220 5020 2280
rect 5080 2220 5100 2280
rect 5160 2220 5240 2280
rect 5300 2220 5320 2280
rect 5380 2220 5400 2280
rect 5000 2180 5400 2220
rect 5000 2120 5020 2180
rect 5080 2120 5100 2180
rect 5160 2120 5240 2180
rect 5300 2120 5320 2180
rect 5380 2120 5400 2180
rect 5000 2100 5400 2120
rect 2400 -1860 4920 -1800
rect 2400 -1940 2540 -1860
rect 2620 -1940 2660 -1860
rect 2740 -1940 2780 -1860
rect 2860 -1940 2900 -1860
rect 2980 -1940 3020 -1860
rect 3100 -1940 3140 -1860
rect 3220 -1940 3260 -1860
rect 3340 -1940 3380 -1860
rect 3460 -1940 3500 -1860
rect 3580 -1940 3620 -1860
rect 3700 -1940 3740 -1860
rect 3820 -1940 3860 -1860
rect 3940 -1940 3980 -1860
rect 4060 -1940 4100 -1860
rect 4180 -1940 4220 -1860
rect 4300 -1940 4340 -1860
rect 4420 -1940 4460 -1860
rect 4540 -1940 4580 -1860
rect 4660 -1940 4700 -1860
rect 4780 -1940 4820 -1860
rect 4900 -1940 4920 -1860
rect 2400 -1980 4920 -1940
rect 2400 -2060 2420 -1980
rect 2500 -2060 2540 -1980
rect 2620 -2060 2660 -1980
rect 2740 -2060 2780 -1980
rect 2860 -2060 2900 -1980
rect 2980 -2060 3020 -1980
rect 3100 -2060 3140 -1980
rect 3220 -2060 3260 -1980
rect 3340 -2060 3380 -1980
rect 3460 -2060 3500 -1980
rect 3580 -2060 3620 -1980
rect 3700 -2060 3740 -1980
rect 3820 -2060 3860 -1980
rect 3940 -2060 3980 -1980
rect 4060 -2060 4100 -1980
rect 4180 -2060 4220 -1980
rect 4300 -2060 4340 -1980
rect 4420 -2060 4460 -1980
rect 4540 -2060 4580 -1980
rect 4660 -2060 4700 -1980
rect 4780 -2060 4820 -1980
rect 4900 -2060 4920 -1980
rect 2400 -2100 4920 -2060
rect 2400 -2180 2420 -2100
rect 2500 -2180 2540 -2100
rect 2620 -2180 2660 -2100
rect 2740 -2180 2780 -2100
rect 2860 -2180 2900 -2100
rect 2980 -2180 3020 -2100
rect 3100 -2180 3140 -2100
rect 3220 -2180 3260 -2100
rect 3340 -2180 3380 -2100
rect 3460 -2180 3500 -2100
rect 3580 -2180 3620 -2100
rect 3700 -2180 3740 -2100
rect 3820 -2180 3860 -2100
rect 3940 -2180 3980 -2100
rect 4060 -2180 4100 -2100
rect 4180 -2180 4220 -2100
rect 4300 -2180 4340 -2100
rect 4420 -2180 4460 -2100
rect 4540 -2180 4580 -2100
rect 4660 -2180 4700 -2100
rect 4780 -2180 4820 -2100
rect 4900 -2180 4920 -2100
rect 2400 -2200 4920 -2180
rect 5480 -1860 8000 -1800
rect 5480 -1940 5500 -1860
rect 5580 -1940 5620 -1860
rect 5700 -1940 5740 -1860
rect 5820 -1940 5860 -1860
rect 5940 -1940 5980 -1860
rect 6060 -1940 6100 -1860
rect 6180 -1940 6220 -1860
rect 6300 -1940 6340 -1860
rect 6420 -1940 6460 -1860
rect 6540 -1940 6580 -1860
rect 6660 -1940 6700 -1860
rect 6780 -1940 6820 -1860
rect 6900 -1940 6940 -1860
rect 7020 -1940 7060 -1860
rect 7140 -1940 7180 -1860
rect 7260 -1940 7300 -1860
rect 7380 -1940 7420 -1860
rect 7500 -1940 7540 -1860
rect 7620 -1940 7660 -1860
rect 7740 -1940 7780 -1860
rect 7860 -1940 7900 -1860
rect 7980 -1940 8000 -1860
rect 5480 -1980 8000 -1940
rect 5480 -2060 5500 -1980
rect 5580 -2060 5620 -1980
rect 5700 -2060 5740 -1980
rect 5820 -2060 5860 -1980
rect 5940 -2060 5980 -1980
rect 6060 -2060 6100 -1980
rect 6180 -2060 6220 -1980
rect 6300 -2060 6340 -1980
rect 6420 -2060 6460 -1980
rect 6540 -2060 6580 -1980
rect 6660 -2060 6700 -1980
rect 6780 -2060 6820 -1980
rect 6900 -2060 6940 -1980
rect 7020 -2060 7060 -1980
rect 7140 -2060 7180 -1980
rect 7260 -2060 7300 -1980
rect 7380 -2060 7420 -1980
rect 7500 -2060 7540 -1980
rect 7620 -2060 7660 -1980
rect 7740 -2060 7780 -1980
rect 7860 -2060 7900 -1980
rect 7980 -2060 8000 -1980
rect 5480 -2100 8000 -2060
rect 5480 -2180 5500 -2100
rect 5580 -2180 5620 -2100
rect 5700 -2180 5740 -2100
rect 5820 -2180 5860 -2100
rect 5940 -2180 5980 -2100
rect 6060 -2180 6100 -2100
rect 6180 -2180 6220 -2100
rect 6300 -2180 6340 -2100
rect 6420 -2180 6460 -2100
rect 6540 -2180 6580 -2100
rect 6660 -2180 6700 -2100
rect 6780 -2180 6820 -2100
rect 6900 -2180 6940 -2100
rect 7020 -2180 7060 -2100
rect 7140 -2180 7180 -2100
rect 7260 -2180 7300 -2100
rect 7380 -2180 7420 -2100
rect 7500 -2180 7540 -2100
rect 7620 -2180 7660 -2100
rect 7740 -2180 7780 -2100
rect 7860 -2180 7900 -2100
rect 7980 -2180 8000 -2100
rect 5480 -2200 8000 -2180
<< via1 >>
rect 5020 2220 5080 2280
rect 5100 2220 5160 2280
rect 5240 2220 5300 2280
rect 5320 2220 5380 2280
rect 5020 2120 5080 2180
rect 5100 2120 5160 2180
rect 5240 2120 5300 2180
rect 5320 2120 5380 2180
<< metal2 >>
rect 1400 3500 2000 3900
rect 8400 3500 9000 3900
rect 1400 1800 1600 3500
rect 1700 2280 8700 2300
rect 1700 2220 5020 2280
rect 5080 2220 5100 2280
rect 5160 2220 5240 2280
rect 5300 2220 5320 2280
rect 5380 2220 8700 2280
rect 1700 2180 8700 2220
rect 1700 2120 5020 2180
rect 5080 2120 5100 2180
rect 5160 2120 5240 2180
rect 5300 2120 5320 2180
rect 5380 2120 8700 2180
rect 1700 2100 8700 2120
rect 1700 1800 1900 2100
rect 8500 1800 8700 2100
rect 8800 1800 9000 3500
rect 5100 -3320 5300 -1900
use differential-pair  differential-pair_0
timestamp 1769952370
transform 1 0 1100 0 1 -1600
box 300 -500 7900 3600
use mirror-load  mirror-load_0
timestamp 1770000594
transform 1 0 840 0 1 2540
box 900 -500 7800 2340
use y  y_0
timestamp 1770003475
transform 1 0 104 0 1 -3222
box 1800 -1800 8400 1100
<< end >>
