magic
tech sky130A
magscale 1 2
timestamp 1769436194
<< nwell >>
rect 1200 5779 8120 5800
rect 1200 5774 31295 5779
rect 1200 2869 37920 5774
rect 1200 2417 37925 2869
rect 1200 2400 7629 2417
rect 31026 83 37925 2417
<< pwell >>
rect 7629 2400 30971 2417
rect 1200 73 30971 2400
rect 32438 73 37935 77
rect 1200 -2436 37935 73
rect 1200 -2800 8120 -2436
rect 31040 -2826 37935 -2436
rect 32438 -2999 37935 -2826
<< psubdiff >>
rect 2600 1560 6000 1600
rect 2600 1440 2800 1560
rect 5800 1440 6000 1560
rect 2600 1400 6000 1440
rect 2600 0 2640 1400
rect 2760 0 2800 1400
rect 5800 0 5840 1400
rect 5960 0 6000 1400
rect 1400 -40 7200 0
rect 1400 -160 1600 -40
rect 7000 -160 7200 -40
rect 1400 -200 7200 -160
rect 1400 -2480 1440 -200
rect 1560 -2480 1600 -200
rect 7000 -2480 7040 -200
rect 7160 -2480 7200 -200
rect 1400 -2520 7200 -2480
rect 1400 -2620 1600 -2520
rect 7000 -2620 7200 -2520
rect 1400 -2660 7200 -2620
rect 33000 -240 36400 -200
rect 33000 -360 33200 -240
rect 36200 -360 36400 -240
rect 33000 -400 36400 -360
rect 33000 -2460 33040 -400
rect 33160 -2460 33200 -400
rect 36200 -2460 36240 -400
rect 36360 -2460 36400 -400
rect 33000 -2500 36400 -2460
rect 33000 -2600 33200 -2500
rect 36200 -2600 36400 -2500
rect 33000 -2640 36400 -2600
rect 36200 -2660 36400 -2640
<< nsubdiff >>
rect 1400 5640 7400 5680
rect 1400 5540 1600 5640
rect 7200 5540 7400 5640
rect 1400 5500 7400 5540
rect 1400 3000 1440 5500
rect 1560 3000 1600 5500
rect 7200 3000 7240 5500
rect 7360 3000 7400 5500
rect 1400 2960 7400 3000
rect 1400 2840 1600 2960
rect 7200 2840 7400 2960
rect 1400 2800 7400 2840
rect 31720 5660 37720 5700
rect 31720 5560 31920 5660
rect 37520 5560 37720 5660
rect 31720 5540 37720 5560
rect 31720 5520 37560 5540
rect 31720 2760 31760 5520
rect 31880 2774 31920 5520
rect 37520 2780 37560 5520
rect 37680 2780 37720 5540
rect 37520 2774 37720 2780
rect 31880 2760 37720 2774
rect 31720 2740 37720 2760
rect 31720 2620 31920 2740
rect 37520 2620 37720 2740
rect 31720 2574 37720 2620
rect 33600 2560 33800 2574
rect 33600 800 33640 2560
rect 33760 800 33800 2560
rect 35300 2560 35500 2574
rect 37520 2560 37720 2574
rect 35300 800 35340 2560
rect 35460 800 35500 2560
rect 33600 760 35500 800
rect 33600 640 33800 760
rect 35300 640 35500 760
rect 33600 600 35500 640
<< psubdiffcont >>
rect 2800 1440 5800 1560
rect 2640 0 2760 1400
rect 5840 0 5960 1400
rect 1600 -160 7000 -40
rect 1440 -2480 1560 -200
rect 7040 -2480 7160 -200
rect 1600 -2620 7000 -2520
rect 33200 -360 36200 -240
rect 33040 -2460 33160 -400
rect 36240 -2460 36360 -400
rect 33200 -2600 36200 -2500
<< nsubdiffcont >>
rect 1600 5540 7200 5640
rect 1440 3000 1560 5500
rect 7240 3000 7360 5500
rect 1600 2840 7200 2960
rect 31920 5560 37520 5660
rect 31760 2760 31880 5520
rect 37560 2780 37680 5540
rect 31920 2620 37520 2740
rect 33640 800 33760 2560
rect 35340 800 35460 2560
rect 33800 640 35300 760
<< locali >>
rect 1000 7000 38000 7200
rect 1000 6800 1200 7000
rect 1018 6400 1200 6800
rect 2400 6400 2600 7000
rect 3800 6400 4000 7000
rect 5200 6400 5400 7000
rect 6600 6400 6800 7000
rect 8000 6400 8200 7000
rect 9400 6400 9600 7000
rect 10800 6400 11000 7000
rect 12200 6400 12400 7000
rect 13600 6400 13800 7000
rect 15000 6400 15200 7000
rect 16400 6400 16600 7000
rect 17800 6400 18000 7000
rect 19200 6400 19400 7000
rect 20600 6400 20800 7000
rect 22000 6400 22200 7000
rect 23400 6400 23600 7000
rect 24800 6400 25000 7000
rect 26200 6400 26400 7000
rect 27600 6400 27800 7000
rect 29000 6400 29200 7000
rect 30400 6400 30600 7000
rect 31800 6400 32000 7000
rect 33200 6400 33400 7000
rect 34600 6400 34800 7000
rect 36000 6400 36200 7000
rect 37400 6800 38000 7000
rect 37400 6400 37936 6800
rect 1018 6200 37936 6400
rect 1018 5600 1200 6200
rect 2400 5640 2600 6200
rect 3800 5640 4000 6200
rect 5200 5640 5400 6200
rect 6600 5640 6800 6200
rect 8000 5600 8200 6200
rect 9400 5600 9600 6200
rect 10800 5600 11000 6200
rect 12200 5600 12400 6200
rect 13600 5600 13800 6200
rect 15000 5600 15200 6200
rect 16400 5600 16600 6200
rect 17800 5600 18000 6200
rect 19200 5600 19400 6200
rect 20600 5600 20800 6200
rect 22000 5600 22200 6200
rect 23400 5600 23600 6200
rect 24800 5600 25000 6200
rect 26200 5600 26400 6200
rect 27600 5600 27800 6200
rect 29000 5600 29200 6200
rect 30400 5600 30600 6200
rect 31800 5660 32000 6200
rect 33200 5660 33400 6200
rect 34600 5660 34800 6200
rect 36000 5660 36200 6200
rect 37400 5660 37936 6200
rect 31800 5600 31920 5660
rect 1018 5540 1600 5600
rect 7200 5560 31920 5600
rect 37520 5560 37936 5660
rect 7200 5540 37936 5560
rect 1018 5520 37560 5540
rect 1018 5500 31760 5520
rect 1018 5390 1440 5500
rect 1400 3000 1440 5390
rect 1560 5390 7240 5500
rect 1560 3000 1600 5390
rect 2106 3304 2245 5390
rect 2716 3309 2855 5390
rect 3332 3309 3471 5390
rect 3952 3304 4091 5390
rect 4567 3309 4706 5390
rect 5187 3304 5326 5390
rect 5798 3304 5937 5390
rect 6413 3304 6552 5390
rect 7200 3000 7240 5390
rect 7360 5390 31760 5500
rect 7360 3000 7400 5390
rect 31040 5374 31760 5390
rect 1400 2960 7400 3000
rect 1400 2840 1600 2960
rect 7200 2840 7400 2960
rect 1400 2800 7400 2840
rect 31720 2760 31760 5374
rect 31880 5374 37560 5520
rect 31880 2774 31920 5374
rect 32400 3100 32600 5374
rect 33000 3100 33200 5374
rect 33600 3100 33800 5374
rect 34200 3100 34400 5374
rect 34900 3100 35100 5374
rect 35500 3100 35700 5374
rect 36100 3100 36300 5374
rect 36700 3100 36900 5374
rect 37520 2780 37560 5374
rect 37680 5390 37936 5540
rect 37680 5374 37920 5390
rect 37680 2780 37720 5374
rect 37520 2774 37720 2780
rect 31880 2760 37720 2774
rect 31720 2740 37720 2760
rect 31720 2620 31920 2740
rect 37520 2620 37720 2740
rect 31720 2574 37720 2620
rect 33600 2560 33800 2574
rect 2600 1560 6000 1600
rect 2600 1440 2800 1560
rect 5800 1440 6000 1560
rect 2600 1400 6000 1440
rect 2600 0 2640 1400
rect 2760 0 2800 1400
rect 3083 0 5480 1
rect 5800 0 5840 1400
rect 5960 0 6000 1400
rect 33600 800 33640 2560
rect 33760 800 33800 2560
rect 35300 2560 35500 2574
rect 35300 800 35340 2560
rect 35460 800 35500 2560
rect 33600 760 35500 800
rect 33600 640 33800 760
rect 35300 640 35500 760
rect 33600 600 35500 640
rect 1400 -40 7200 0
rect 1400 -160 1600 -40
rect 7000 -160 7200 -40
rect 1400 -200 7200 -160
rect 1400 -2382 1440 -200
rect 1018 -2400 1440 -2382
rect 1560 -2382 1600 -200
rect 1944 -619 6809 -528
rect 2083 -2382 2191 -668
rect 2704 -2382 2798 -668
rect 3316 -2382 3412 -668
rect 3931 -2382 4027 -669
rect 4550 -2382 4646 -669
rect 5163 -2382 5259 -669
rect 5785 -2382 5881 -672
rect 6401 -2382 6497 -669
rect 7000 -2382 7040 -200
rect 1560 -2400 7040 -2382
rect 7160 -2382 7200 -200
rect 33005 -240 36396 -194
rect 33005 -360 33200 -240
rect 36200 -360 36396 -240
rect 33005 -394 36396 -360
rect 33005 -400 33205 -394
rect 33005 -2361 33040 -400
rect 32438 -2382 33040 -2361
rect 7160 -2400 33040 -2382
rect 1018 -3000 1200 -2400
rect 2400 -2520 2600 -2400
rect 3800 -2520 4000 -2400
rect 5200 -2520 5400 -2400
rect 6600 -2520 6800 -2400
rect 2400 -3000 2600 -2620
rect 3800 -3000 4000 -2620
rect 5200 -3000 5400 -2620
rect 6600 -3000 6800 -2620
rect 8000 -3000 8200 -2400
rect 10600 -3000 10800 -2400
rect 12000 -3000 12200 -2400
rect 13400 -3000 13600 -2400
rect 14800 -3000 15000 -2400
rect 16200 -3000 16400 -2400
rect 17600 -3000 17800 -2400
rect 19000 -3000 19200 -2400
rect 20400 -3000 20600 -2400
rect 21800 -3000 22000 -2400
rect 23200 -3000 23400 -2400
rect 24600 -3000 24800 -2400
rect 26000 -3000 26200 -2400
rect 27400 -3000 27600 -2400
rect 28800 -3000 29000 -2400
rect 30200 -3000 30400 -2400
rect 31600 -3000 31800 -2400
rect 33000 -2460 33040 -2400
rect 33160 -2361 33205 -400
rect 36205 -400 36396 -394
rect 33686 -2361 33787 -673
rect 34306 -2361 34407 -665
rect 34920 -2361 35021 -668
rect 35536 -2361 35637 -665
rect 36205 -2361 36240 -400
rect 33160 -2400 36240 -2361
rect 36360 -2361 36396 -400
rect 36360 -2382 37935 -2361
rect 36360 -2400 37936 -2382
rect 33160 -2460 33200 -2400
rect 33000 -3000 33200 -2460
rect 34400 -2500 34600 -2400
rect 35800 -2500 36000 -2400
rect 34400 -3000 34600 -2600
rect 35800 -3000 36000 -2600
rect 37200 -3000 38000 -2400
rect 1018 -3200 38000 -3000
rect 1018 -3600 1200 -3200
rect 1000 -3800 1200 -3600
rect 2400 -3800 2600 -3200
rect 3800 -3800 4000 -3200
rect 5200 -3800 5400 -3200
rect 6600 -3800 6800 -3200
rect 8000 -3800 8200 -3200
rect 10600 -3800 10800 -3200
rect 12000 -3800 12200 -3200
rect 13400 -3800 13600 -3200
rect 14800 -3800 15000 -3200
rect 16200 -3800 16400 -3200
rect 17600 -3800 17800 -3200
rect 19000 -3800 19200 -3200
rect 20400 -3800 20600 -3200
rect 21800 -3800 22000 -3200
rect 23200 -3800 23400 -3200
rect 24600 -3800 24800 -3200
rect 26000 -3800 26200 -3200
rect 27400 -3800 27600 -3200
rect 28800 -3800 29000 -3200
rect 30200 -3800 30400 -3200
rect 31600 -3800 31800 -3200
rect 33000 -3800 33200 -3200
rect 34400 -3800 34600 -3200
rect 35800 -3800 36000 -3200
rect 37200 -3800 38000 -3200
rect 1000 -4200 38000 -3800
<< viali >>
rect 1200 6400 2400 7000
rect 2600 6400 3800 7000
rect 4000 6400 5200 7000
rect 5400 6400 6600 7000
rect 6800 6400 8000 7000
rect 8200 6400 9400 7000
rect 9600 6400 10800 7000
rect 11000 6400 12200 7000
rect 12400 6400 13600 7000
rect 13800 6400 15000 7000
rect 15200 6400 16400 7000
rect 16600 6400 17800 7000
rect 18000 6400 19200 7000
rect 19400 6400 20600 7000
rect 20800 6400 22000 7000
rect 22200 6400 23400 7000
rect 23600 6400 24800 7000
rect 25000 6400 26200 7000
rect 26400 6400 27600 7000
rect 27800 6400 29000 7000
rect 29200 6400 30400 7000
rect 30600 6400 31800 7000
rect 32000 6400 33200 7000
rect 33400 6400 34600 7000
rect 34800 6400 36000 7000
rect 36200 6400 37400 7000
rect 1200 5640 2400 6200
rect 2600 5640 3800 6200
rect 4000 5640 5200 6200
rect 5400 5640 6600 6200
rect 6800 5640 8000 6200
rect 1200 5600 1600 5640
rect 1600 5600 2400 5640
rect 2600 5600 3800 5640
rect 4000 5600 5200 5640
rect 5400 5600 6600 5640
rect 6800 5600 7200 5640
rect 7200 5600 8000 5640
rect 8200 5600 9400 6200
rect 9600 5600 10800 6200
rect 11000 5600 12200 6200
rect 12400 5600 13600 6200
rect 13800 5600 15000 6200
rect 15200 5600 16400 6200
rect 16600 5600 17800 6200
rect 18000 5600 19200 6200
rect 19400 5600 20600 6200
rect 20800 5600 22000 6200
rect 22200 5600 23400 6200
rect 23600 5600 24800 6200
rect 25000 5600 26200 6200
rect 26400 5600 27600 6200
rect 27800 5600 29000 6200
rect 29200 5600 30400 6200
rect 30600 5600 31800 6200
rect 32000 5660 33200 6200
rect 33400 5660 34600 6200
rect 34800 5660 36000 6200
rect 36200 5660 37400 6200
rect 32000 5600 33200 5660
rect 33400 5600 34600 5660
rect 34800 5600 36000 5660
rect 36200 5600 37400 5660
rect 1200 -2480 1440 -2400
rect 1440 -2480 1560 -2400
rect 1560 -2480 2400 -2400
rect 1200 -2520 2400 -2480
rect 2600 -2520 3800 -2400
rect 4000 -2520 5200 -2400
rect 5400 -2520 6600 -2400
rect 6800 -2480 7040 -2400
rect 7040 -2480 7160 -2400
rect 7160 -2480 8000 -2400
rect 6800 -2520 8000 -2480
rect 1200 -2620 1600 -2520
rect 1600 -2620 2400 -2520
rect 2600 -2620 3800 -2520
rect 4000 -2620 5200 -2520
rect 5400 -2620 6600 -2520
rect 6800 -2620 7000 -2520
rect 7000 -2620 8000 -2520
rect 1200 -3000 2400 -2620
rect 2600 -3000 3800 -2620
rect 4000 -3000 5200 -2620
rect 5400 -3000 6600 -2620
rect 6800 -3000 8000 -2620
rect 8200 -3000 10600 -2400
rect 10800 -3000 12000 -2400
rect 12200 -3000 13400 -2400
rect 13600 -3000 14800 -2400
rect 15000 -3000 16200 -2400
rect 16400 -3000 17600 -2400
rect 17800 -3000 19000 -2400
rect 19200 -3000 20400 -2400
rect 20600 -3000 21800 -2400
rect 22000 -3000 23200 -2400
rect 23400 -3000 24600 -2400
rect 24800 -3000 26000 -2400
rect 26200 -3000 27400 -2400
rect 27600 -3000 28800 -2400
rect 29000 -3000 30200 -2400
rect 30400 -3000 31600 -2400
rect 31800 -3000 33000 -2400
rect 33200 -2500 34400 -2400
rect 34600 -2500 35800 -2400
rect 36000 -2460 36240 -2400
rect 36240 -2460 36360 -2400
rect 36360 -2460 37200 -2400
rect 36000 -2500 37200 -2460
rect 33200 -2600 34400 -2500
rect 34600 -2600 35800 -2500
rect 36000 -2600 36200 -2500
rect 36200 -2600 37200 -2500
rect 33200 -3000 34400 -2600
rect 34600 -3000 35800 -2600
rect 36000 -3000 37200 -2600
rect 1200 -3800 2400 -3200
rect 2600 -3800 3800 -3200
rect 4000 -3800 5200 -3200
rect 5400 -3800 6600 -3200
rect 6800 -3800 8000 -3200
rect 8200 -3800 10600 -3200
rect 10800 -3800 12000 -3200
rect 12200 -3800 13400 -3200
rect 13600 -3800 14800 -3200
rect 15000 -3800 16200 -3200
rect 16400 -3800 17600 -3200
rect 17800 -3800 19000 -3200
rect 19200 -3800 20400 -3200
rect 20600 -3800 21800 -3200
rect 22000 -3800 23200 -3200
rect 23400 -3800 24600 -3200
rect 24800 -3800 26000 -3200
rect 26200 -3800 27400 -3200
rect 27600 -3800 28800 -3200
rect 29000 -3800 30200 -3200
rect 30400 -3800 31600 -3200
rect 31800 -3800 33000 -3200
rect 33200 -3800 34400 -3200
rect 34600 -3800 35800 -3200
rect 36000 -3800 37200 -3200
<< metal1 >>
rect 1000 7000 38000 7200
rect 1000 6800 1200 7000
rect 1020 6700 1200 6800
rect 1018 6400 1200 6700
rect 2400 6400 2600 7000
rect 3800 6400 4000 7000
rect 5200 6400 5400 7000
rect 6600 6400 6800 7000
rect 8000 6400 8200 7000
rect 9400 6400 9600 7000
rect 10800 6400 11000 7000
rect 12200 6400 12400 7000
rect 13600 6400 13800 7000
rect 15000 6400 15200 7000
rect 16400 6400 16600 7000
rect 17800 6400 18000 7000
rect 19200 6400 19400 7000
rect 20600 6400 20800 7000
rect 22000 6400 22200 7000
rect 23400 6400 23600 7000
rect 24800 6400 25000 7000
rect 26200 6400 26400 7000
rect 27600 6400 27800 7000
rect 29000 6400 29200 7000
rect 30400 6400 30600 7000
rect 31800 6400 32000 7000
rect 33200 6400 33400 7000
rect 34600 6400 34800 7000
rect 36000 6400 36200 7000
rect 37400 6800 38000 7000
rect 37400 6400 37936 6800
rect 1018 6200 37936 6400
rect 1018 5600 1200 6200
rect 2400 5600 2600 6200
rect 3800 5600 4000 6200
rect 5200 5600 5400 6200
rect 6600 5600 6800 6200
rect 8000 5600 8200 6200
rect 9400 5600 9600 6200
rect 10800 5600 11000 6200
rect 12200 5600 12400 6200
rect 13600 5600 13800 6200
rect 15000 5600 15200 6200
rect 16400 5600 16600 6200
rect 17800 5600 18000 6200
rect 19200 5600 19400 6200
rect 20600 5600 20800 6200
rect 22000 5600 22200 6200
rect 23400 5600 23600 6200
rect 24800 5600 25000 6200
rect 26200 5600 26400 6200
rect 27600 5600 27800 6200
rect 29000 5600 29200 6200
rect 30400 5600 30600 6200
rect 31800 5600 32000 6200
rect 33200 5600 33400 6200
rect 34600 5600 34800 6200
rect 36000 5600 36200 6200
rect 37400 5600 37936 6200
rect 1018 5390 37936 5600
rect 31040 5374 37920 5390
rect 1759 3240 1900 5220
rect 3026 3240 3167 5222
rect 4256 3240 4397 5218
rect 5493 3240 5634 5218
rect 6751 3240 6892 5214
rect 32100 4460 32300 4500
rect 32100 4300 32120 4460
rect 32280 4300 32300 4460
rect 32100 4220 32300 4300
rect 32100 4060 32120 4220
rect 32280 4060 32300 4220
rect 32100 3980 32300 4060
rect 32100 3820 32120 3980
rect 32280 3820 32300 3980
rect 32100 3800 32300 3820
rect 32700 4460 32900 4500
rect 32700 4300 32720 4460
rect 32880 4300 32900 4460
rect 32700 4220 32900 4300
rect 32700 4060 32720 4220
rect 32880 4060 32900 4220
rect 32700 3980 32900 4060
rect 32700 3820 32720 3980
rect 32880 3820 32900 3980
rect 32700 3800 32900 3820
rect 33300 4460 33500 4500
rect 33300 4300 33320 4460
rect 33480 4300 33500 4460
rect 33300 4220 33500 4300
rect 33300 4060 33320 4220
rect 33480 4060 33500 4220
rect 33300 3980 33500 4060
rect 33300 3820 33320 3980
rect 33480 3820 33500 3980
rect 33300 3800 33500 3820
rect 33900 4460 34100 4500
rect 33900 4300 33920 4460
rect 34080 4300 34100 4460
rect 33900 4220 34100 4300
rect 33900 4060 33920 4220
rect 34080 4060 34100 4220
rect 33900 3980 34100 4060
rect 33900 3820 33920 3980
rect 34080 3820 34100 3980
rect 33900 3800 34100 3820
rect 34600 4460 34800 4500
rect 34600 4300 34620 4460
rect 34780 4300 34800 4460
rect 34600 4220 34800 4300
rect 34600 4060 34620 4220
rect 34780 4060 34800 4220
rect 34600 3980 34800 4060
rect 34600 3820 34620 3980
rect 34780 3820 34800 3980
rect 34600 3800 34800 3820
rect 35200 4460 35400 4500
rect 35200 4300 35220 4460
rect 35380 4300 35400 4460
rect 35200 4220 35400 4300
rect 35200 4060 35220 4220
rect 35380 4060 35400 4220
rect 35200 3980 35400 4060
rect 35200 3820 35220 3980
rect 35380 3820 35400 3980
rect 35200 3800 35400 3820
rect 35800 4460 36000 4500
rect 35800 4300 35820 4460
rect 35980 4300 36000 4460
rect 35800 4220 36000 4300
rect 35800 4060 35820 4220
rect 35980 4060 36000 4220
rect 35800 3980 36000 4060
rect 35800 3820 35820 3980
rect 35980 3820 36000 3980
rect 35800 3800 36000 3820
rect 36400 4440 36600 4500
rect 36400 4280 36420 4440
rect 36580 4280 36600 4440
rect 36400 4220 36600 4280
rect 36400 4060 36420 4220
rect 36580 4060 36600 4220
rect 36400 3980 36600 4060
rect 36400 3820 36420 3980
rect 36580 3820 36600 3980
rect 36400 3800 36600 3820
rect 37000 4440 37200 4500
rect 37000 4280 37020 4440
rect 37180 4280 37200 4440
rect 37000 4220 37200 4280
rect 37000 4060 37020 4220
rect 37180 4060 37200 4220
rect 37000 3980 37200 4060
rect 37000 3820 37020 3980
rect 37180 3820 37200 3980
rect 37000 3800 37200 3820
rect 1759 3139 6894 3240
rect -320 2280 -120 2300
rect -320 2220 -300 2280
rect -240 2220 -200 2280
rect -140 2220 -120 2280
rect -320 2180 -120 2220
rect -320 2120 -300 2180
rect -240 2120 -200 2180
rect -140 2120 -120 2180
rect -320 2100 -120 2120
rect -320 1880 -120 1900
rect -320 1820 -300 1880
rect -240 1820 -200 1880
rect -140 1820 -120 1880
rect -320 1780 -120 1820
rect -320 1720 -300 1780
rect -240 1720 -200 1780
rect -140 1720 -120 1780
rect -320 1700 -120 1720
rect 2940 1440 3100 3139
rect 3580 1440 3740 3139
rect 4200 1440 4360 3139
rect 4840 1440 5000 3139
rect 5480 1440 5640 3139
rect 30449 3043 30881 3595
rect 30378 2941 36997 3043
rect 30449 2325 30881 2941
rect 34260 1700 34400 1720
rect 34260 1600 34280 1700
rect 34380 1600 34400 1700
rect 34260 1540 34400 1600
rect 34260 1440 34280 1540
rect 34380 1440 34400 1540
rect 3012 201 3040 1440
rect 3076 1362 3612 1363
rect 3076 1345 3614 1362
rect 3076 1292 3078 1345
rect 3134 1299 3614 1345
rect 3134 1292 3141 1299
rect 3076 1263 3141 1292
rect 3076 1210 3079 1263
rect 3135 1210 3141 1263
rect 3076 1201 3141 1210
rect 3231 1199 3460 1261
rect 3549 1202 3614 1299
rect 3140 -325 3234 1151
rect 3452 -325 3546 1156
rect 3645 196 3673 1440
rect 3706 1343 4247 1361
rect 3706 1341 3714 1343
rect 3705 1290 3714 1341
rect 3770 1298 4247 1343
rect 3770 1290 3776 1298
rect 3705 1263 3776 1290
rect 3705 1210 3716 1263
rect 3772 1210 3776 1263
rect 3705 1202 3776 1210
rect 3862 1196 4092 1260
rect 4179 1207 4247 1298
rect 3770 -325 3864 1161
rect 4088 -325 4182 1159
rect 4275 201 4303 1440
rect 4339 1362 4403 1363
rect 4339 1345 4881 1362
rect 4339 1308 4820 1345
rect 4339 1203 4403 1308
rect 4817 1292 4820 1308
rect 4876 1292 4881 1345
rect 4494 1200 4724 1264
rect 4817 1260 4881 1292
rect 4817 1207 4820 1260
rect 4876 1207 4883 1260
rect 4817 1202 4883 1207
rect 4872 1200 4883 1202
rect 4405 -325 4499 1159
rect 4722 -325 4816 1163
rect 4912 197 4940 1440
rect 4972 1345 5514 1362
rect 4972 1308 5450 1345
rect 4972 1202 5054 1308
rect 5431 1292 5450 1308
rect 5506 1308 5514 1345
rect 5506 1292 5513 1308
rect 5111 1259 5360 1265
rect 5431 1262 5513 1292
rect 5111 1202 5362 1259
rect 5431 1209 5450 1262
rect 5506 1209 5513 1262
rect 5431 1203 5513 1209
rect 5111 1200 5360 1202
rect 5033 -325 5127 1156
rect 5353 -325 5447 1163
rect 5545 199 5573 1440
rect 34260 1380 34400 1440
rect 34260 1280 34280 1380
rect 34380 1280 34400 1380
rect 34260 1240 34400 1280
rect 34740 1700 34880 1720
rect 34740 1600 34760 1700
rect 34860 1600 34880 1700
rect 34740 1540 34880 1600
rect 34740 1440 34760 1540
rect 34860 1440 34880 1540
rect 34740 1380 34880 1440
rect 38100 1580 38300 1600
rect 38100 1520 38120 1580
rect 38180 1520 38220 1580
rect 38280 1520 38300 1580
rect 38100 1480 38300 1520
rect 38100 1420 38120 1480
rect 38180 1420 38220 1480
rect 38280 1420 38300 1480
rect 38100 1400 38300 1420
rect 34740 1280 34760 1380
rect 34860 1280 34880 1380
rect 34740 1240 34880 1280
rect 34020 940 36400 1160
rect 2403 -326 6191 -325
rect 2403 -328 6193 -326
rect 2399 -412 6193 -328
rect -320 -460 -120 -440
rect -320 -520 -300 -460
rect -240 -520 -200 -460
rect -140 -520 -120 -460
rect 1759 -480 2331 -458
rect 1759 -497 1760 -480
rect -320 -560 -120 -520
rect -320 -620 -300 -560
rect -240 -620 -200 -560
rect -140 -620 -120 -560
rect 1757 -561 1760 -497
rect -320 -640 -120 -620
rect 1756 -600 1760 -561
rect 1880 -600 1980 -480
rect 2100 -600 2200 -480
rect 2320 -600 2331 -480
rect 2399 -497 2489 -412
rect 2539 -480 3569 -463
rect 1756 -641 2331 -600
rect 1756 -645 2330 -641
rect 1757 -2202 1852 -645
rect 1760 -2235 1847 -2202
rect 2397 -2204 2493 -497
rect 2539 -555 2560 -480
rect 2535 -600 2560 -555
rect 2680 -600 2780 -480
rect 2920 -600 3000 -480
rect 3120 -600 3200 -480
rect 3340 -600 3420 -480
rect 3540 -551 3569 -480
rect 3631 -497 3721 -412
rect 3793 -480 4791 -461
rect 3629 -498 3725 -497
rect 3540 -600 3571 -551
rect 2535 -639 3571 -600
rect 3012 -640 3571 -639
rect 3012 -2050 3108 -640
rect 3627 -670 3725 -498
rect 3793 -600 3820 -480
rect 3940 -600 4020 -480
rect 4140 -600 4220 -480
rect 4340 -600 4440 -480
rect 4560 -600 4640 -480
rect 4760 -551 4791 -480
rect 4859 -497 4949 -412
rect 5021 -480 6019 -459
rect 4760 -600 4792 -551
rect 3793 -641 4792 -600
rect 3012 -2204 3110 -2050
rect 3629 -2201 3725 -670
rect 4244 -2195 4340 -641
rect 3013 -2235 3110 -2204
rect 4251 -2235 4335 -2195
rect 4859 -2198 4955 -497
rect 5021 -600 5040 -480
rect 5160 -600 5240 -480
rect 5360 -600 5460 -480
rect 5580 -600 5680 -480
rect 5800 -600 5880 -480
rect 6000 -551 6019 -480
rect 6103 -497 6193 -412
rect 6740 -459 35800 -320
rect 6000 -600 6023 -551
rect 5021 -639 6023 -600
rect 5024 -641 6023 -639
rect 5476 -2048 5572 -641
rect 6094 -648 6193 -497
rect 6259 -480 35800 -459
rect 6259 -555 6280 -480
rect 6255 -600 6280 -555
rect 6400 -600 6480 -480
rect 6600 -600 6680 -480
rect 6800 -600 35800 -480
rect 6255 -620 35800 -600
rect 6255 -637 6813 -620
rect 6255 -641 6811 -637
rect 5475 -2235 5575 -2048
rect 6094 -2192 6190 -648
rect 6715 -2061 6811 -641
rect 33300 -1140 33500 -1100
rect 33300 -1300 33320 -1140
rect 33480 -1300 33500 -1140
rect 33300 -1380 33500 -1300
rect 33300 -1540 33320 -1380
rect 33480 -1540 33500 -1380
rect 33300 -1620 33500 -1540
rect 33300 -1780 33320 -1620
rect 33480 -1780 33500 -1620
rect 33300 -1800 33500 -1780
rect 34000 -1140 34200 -1100
rect 34000 -1300 34020 -1140
rect 34180 -1300 34200 -1140
rect 34000 -1380 34200 -1300
rect 34000 -1540 34020 -1380
rect 34180 -1540 34200 -1380
rect 34000 -1620 34200 -1540
rect 34000 -1780 34020 -1620
rect 34180 -1780 34200 -1620
rect 34000 -1800 34200 -1780
rect 34600 -1140 34800 -1100
rect 34600 -1300 34620 -1140
rect 34780 -1300 34800 -1140
rect 34600 -1380 34800 -1300
rect 34600 -1540 34620 -1380
rect 34780 -1540 34800 -1380
rect 34600 -1620 34800 -1540
rect 34600 -1780 34620 -1620
rect 34780 -1780 34800 -1620
rect 34600 -1800 34800 -1780
rect 35200 -1140 35400 -1100
rect 35200 -1300 35220 -1140
rect 35380 -1300 35400 -1140
rect 35200 -1380 35400 -1300
rect 35200 -1540 35220 -1380
rect 35380 -1540 35400 -1380
rect 35200 -1620 35400 -1540
rect 35200 -1780 35220 -1620
rect 35380 -1780 35400 -1620
rect 35200 -1800 35400 -1780
rect 35800 -1140 36000 -1100
rect 35800 -1300 35820 -1140
rect 35980 -1300 36000 -1140
rect 35800 -1380 36000 -1300
rect 35800 -1540 35820 -1380
rect 35980 -1540 36000 -1380
rect 35800 -1620 36000 -1540
rect 35800 -1780 35820 -1620
rect 35980 -1780 36000 -1620
rect 35800 -1800 36000 -1780
rect 6715 -2198 6816 -2061
rect 6716 -2235 6816 -2198
rect 1760 -2298 6816 -2235
rect 1762 -2313 6816 -2298
rect 1762 -2314 6811 -2313
rect 36160 -2361 36400 940
rect 32438 -2382 37935 -2361
rect 1018 -2400 37936 -2382
rect 1018 -2480 1200 -2400
rect 1020 -2680 1200 -2480
rect 1018 -3000 1200 -2680
rect 2400 -3000 2600 -2400
rect 3800 -3000 4000 -2400
rect 5200 -3000 5400 -2400
rect 6600 -3000 6800 -2400
rect 8000 -3000 8200 -2400
rect 10600 -3000 10800 -2400
rect 12000 -3000 12200 -2400
rect 13400 -3000 13600 -2400
rect 14800 -3000 15000 -2400
rect 16200 -3000 16400 -2400
rect 17600 -3000 17800 -2400
rect 19000 -3000 19200 -2400
rect 20400 -3000 20600 -2400
rect 21800 -3000 22000 -2400
rect 23200 -3000 23400 -2400
rect 24600 -3000 24800 -2400
rect 26000 -3000 26200 -2400
rect 27400 -3000 27600 -2400
rect 28800 -3000 29000 -2400
rect 30200 -3000 30400 -2400
rect 31600 -3000 31800 -2400
rect 33000 -3000 33200 -2400
rect 34400 -3000 34600 -2400
rect 35800 -3000 36000 -2400
rect 37200 -3000 38000 -2400
rect 1018 -3200 38000 -3000
rect 1018 -3600 1200 -3200
rect 1000 -3800 1200 -3600
rect 2400 -3800 2600 -3200
rect 3800 -3800 4000 -3200
rect 5200 -3800 5400 -3200
rect 6600 -3800 6800 -3200
rect 8000 -3800 8200 -3200
rect 10600 -3800 10800 -3200
rect 12000 -3800 12200 -3200
rect 13400 -3800 13600 -3200
rect 14800 -3800 15000 -3200
rect 16200 -3800 16400 -3200
rect 17600 -3800 17800 -3200
rect 19000 -3800 19200 -3200
rect 20400 -3800 20600 -3200
rect 21800 -3800 22000 -3200
rect 23200 -3800 23400 -3200
rect 24600 -3800 24800 -3200
rect 26000 -3800 26200 -3200
rect 27400 -3800 27600 -3200
rect 28800 -3800 29000 -3200
rect 30200 -3800 30400 -3200
rect 31600 -3800 31800 -3200
rect 33000 -3800 33200 -3200
rect 34400 -3800 34600 -3200
rect 35800 -3800 36000 -3200
rect 37200 -3800 38000 -3200
rect 1000 -4200 38000 -3800
<< via1 >>
rect 32120 4300 32280 4460
rect 32120 4060 32280 4220
rect 32120 3820 32280 3980
rect 32720 4300 32880 4460
rect 32720 4060 32880 4220
rect 32720 3820 32880 3980
rect 33320 4300 33480 4460
rect 33320 4060 33480 4220
rect 33320 3820 33480 3980
rect 33920 4300 34080 4460
rect 33920 4060 34080 4220
rect 33920 3820 34080 3980
rect 34620 4300 34780 4460
rect 34620 4060 34780 4220
rect 34620 3820 34780 3980
rect 35220 4300 35380 4460
rect 35220 4060 35380 4220
rect 35220 3820 35380 3980
rect 35820 4300 35980 4460
rect 35820 4060 35980 4220
rect 35820 3820 35980 3980
rect 36420 4280 36580 4440
rect 36420 4060 36580 4220
rect 36420 3820 36580 3980
rect 37020 4280 37180 4440
rect 37020 4060 37180 4220
rect 37020 3820 37180 3980
rect -300 2220 -240 2280
rect -200 2220 -140 2280
rect -300 2120 -240 2180
rect -200 2120 -140 2180
rect -300 1820 -240 1880
rect -200 1820 -140 1880
rect -300 1720 -240 1780
rect -200 1720 -140 1780
rect 34280 1600 34380 1700
rect 34280 1440 34380 1540
rect 3078 1292 3134 1345
rect 3079 1210 3135 1263
rect 3714 1290 3770 1343
rect 3716 1210 3772 1263
rect 4820 1292 4876 1345
rect 4820 1207 4876 1260
rect 5450 1292 5506 1345
rect 5450 1209 5506 1262
rect 34280 1280 34380 1380
rect 34760 1600 34860 1700
rect 34760 1440 34860 1540
rect 38120 1520 38180 1580
rect 38220 1520 38280 1580
rect 38120 1420 38180 1480
rect 38220 1420 38280 1480
rect 34760 1280 34860 1380
rect -300 -520 -240 -460
rect -200 -520 -140 -460
rect -300 -620 -240 -560
rect -200 -620 -140 -560
rect 1760 -600 1880 -480
rect 1980 -600 2100 -480
rect 2200 -600 2320 -480
rect 2560 -600 2680 -480
rect 2780 -600 2920 -480
rect 3000 -600 3120 -480
rect 3200 -600 3340 -480
rect 3420 -600 3540 -480
rect 3820 -600 3940 -480
rect 4020 -600 4140 -480
rect 4220 -600 4340 -480
rect 4440 -600 4560 -480
rect 4640 -600 4760 -480
rect 5040 -600 5160 -480
rect 5240 -600 5360 -480
rect 5460 -600 5580 -480
rect 5680 -600 5800 -480
rect 5880 -600 6000 -480
rect 6280 -600 6400 -480
rect 6480 -600 6600 -480
rect 6680 -600 6800 -480
rect 33320 -1300 33480 -1140
rect 33320 -1540 33480 -1380
rect 33320 -1780 33480 -1620
rect 34020 -1300 34180 -1140
rect 34020 -1540 34180 -1380
rect 34020 -1780 34180 -1620
rect 34620 -1300 34780 -1140
rect 34620 -1540 34780 -1380
rect 34620 -1780 34780 -1620
rect 35220 -1300 35380 -1140
rect 35220 -1540 35380 -1380
rect 35220 -1780 35380 -1620
rect 35820 -1300 35980 -1140
rect 35820 -1540 35980 -1380
rect 35820 -1780 35980 -1620
<< metal2 >>
rect 2360 4540 2600 4560
rect 2360 4380 2400 4540
rect 2560 4380 2600 4540
rect 2360 4300 2600 4380
rect 2360 4120 2400 4300
rect 2560 4120 2600 4300
rect 2360 4040 2600 4120
rect 2360 3880 2400 4040
rect 2560 3880 2600 4040
rect 2360 3860 2600 3880
rect 3600 4540 3840 4560
rect 3600 4380 3640 4540
rect 3800 4380 3840 4540
rect 3600 4300 3840 4380
rect 3600 4120 3640 4300
rect 3800 4120 3840 4300
rect 3600 4040 3840 4120
rect 3600 3880 3640 4040
rect 3800 3880 3840 4040
rect 3600 3860 3840 3880
rect 4820 4540 5060 4560
rect 4820 4380 4860 4540
rect 5020 4380 5060 4540
rect 4820 4300 5060 4380
rect 4820 4120 4860 4300
rect 5020 4120 5060 4300
rect 4820 4040 5060 4120
rect 4820 3880 4860 4040
rect 5020 3880 5060 4040
rect 4820 3860 5060 3880
rect 6060 4540 6300 4560
rect 6060 4380 6100 4540
rect 6260 4380 6300 4540
rect 6060 4300 6300 4380
rect 6060 4120 6100 4300
rect 6260 4120 6300 4300
rect 6060 4040 6300 4120
rect 6060 3880 6100 4040
rect 6260 3880 6300 4040
rect 6060 3860 6300 3880
rect 32000 4460 37800 4500
rect 32000 4300 32120 4460
rect 32280 4300 32720 4460
rect 32880 4300 33320 4460
rect 33480 4300 33920 4460
rect 34080 4300 34620 4460
rect 34780 4300 35220 4460
rect 35380 4300 35820 4460
rect 35980 4440 37800 4460
rect 35980 4300 36420 4440
rect 32000 4280 36420 4300
rect 36580 4280 37020 4440
rect 37180 4280 37800 4440
rect 32000 4220 37800 4280
rect 32000 4060 32120 4220
rect 32280 4060 32720 4220
rect 32880 4060 33320 4220
rect 33480 4060 33920 4220
rect 34080 4060 34620 4220
rect 34780 4060 35220 4220
rect 35380 4060 35820 4220
rect 35980 4060 36420 4220
rect 36580 4060 37020 4220
rect 37180 4060 37800 4220
rect 32000 3980 37800 4060
rect 32000 3820 32120 3980
rect 32280 3820 32720 3980
rect 32880 3820 33320 3980
rect 33480 3820 33920 3980
rect 34080 3820 34620 3980
rect 34780 3820 35220 3980
rect 35380 3820 35820 3980
rect 35980 3820 36420 3980
rect 36580 3820 37020 3980
rect 37180 3820 37800 3980
rect 32000 3800 37800 3820
rect 30449 2325 30881 3595
rect -320 2280 6820 2300
rect -320 2220 -300 2280
rect -240 2220 -200 2280
rect -140 2220 3280 2280
rect -320 2180 3280 2220
rect -320 2120 -300 2180
rect -240 2120 -200 2180
rect -140 2120 3280 2180
rect 3440 2120 3480 2280
rect 3640 2120 3680 2280
rect 3840 2120 3880 2280
rect 4040 2120 4080 2280
rect 4240 2120 4280 2280
rect 4440 2120 4480 2280
rect 4640 2120 4680 2280
rect 4840 2120 4880 2280
rect 5040 2120 5080 2280
rect 5240 2120 6820 2280
rect -320 2100 6820 2120
rect 34020 2240 34160 2260
rect 34020 2140 34040 2240
rect 34140 2140 34160 2240
rect 34020 2060 34160 2140
rect 34020 1960 34040 2060
rect 34140 1960 34160 2060
rect 3076 1900 3142 1902
rect 34020 1900 34160 1960
rect -320 1880 6820 1900
rect -320 1820 -300 1880
rect -240 1820 -200 1880
rect -140 1820 6820 1880
rect -320 1780 6820 1820
rect 34020 1800 34040 1900
rect 34140 1800 34160 1900
rect 34020 1780 34160 1800
rect 34500 2240 34640 2260
rect 34500 2140 34520 2240
rect 34620 2140 34640 2240
rect 34500 2060 34640 2140
rect 34500 1960 34520 2060
rect 34620 1960 34640 2060
rect 34500 1900 34640 1960
rect 34500 1800 34520 1900
rect 34620 1800 34640 1900
rect 34500 1780 34640 1800
rect 34980 2240 35120 2260
rect 34980 2140 35000 2240
rect 35100 2140 35120 2240
rect 34980 2060 35120 2140
rect 34980 1960 35000 2060
rect 35100 1960 35120 2060
rect 34980 1900 35120 1960
rect 34980 1800 35000 1900
rect 35100 1800 35120 1900
rect 34980 1780 35120 1800
rect -320 1720 -300 1780
rect -240 1720 -200 1780
rect -140 1720 6820 1780
rect 37100 1720 37800 3800
rect -320 1700 6820 1720
rect 34040 1700 38300 1720
rect 3076 1362 3142 1700
rect 3707 1362 3773 1700
rect 3074 1345 3144 1362
rect 3074 1292 3078 1345
rect 3134 1292 3144 1345
rect 3074 1263 3144 1292
rect 3706 1343 3778 1362
rect 4815 1361 4880 1700
rect 5448 1363 5513 1700
rect 3706 1290 3714 1343
rect 3770 1290 3778 1343
rect 3228 1263 3460 1267
rect 3074 1210 3079 1263
rect 3135 1210 3144 1263
rect 3074 1200 3144 1210
rect 3227 1256 3460 1263
rect 3227 1255 3388 1256
rect 3227 1195 3236 1255
rect 3299 1196 3388 1255
rect 3451 1196 3460 1256
rect 3706 1263 3778 1290
rect 4814 1345 4883 1361
rect 4814 1292 4820 1345
rect 4876 1292 4883 1345
rect 3706 1210 3716 1263
rect 3772 1210 3778 1263
rect 4494 1261 4724 1264
rect 3706 1205 3778 1210
rect 3860 1255 4093 1260
rect 3860 1254 4021 1255
rect 3299 1195 3460 1196
rect 3227 1189 3460 1195
rect 3860 1194 3872 1254
rect 3935 1195 4021 1254
rect 4084 1195 4093 1255
rect 3935 1194 4093 1195
rect 3860 1186 4093 1194
rect 4493 1255 4726 1261
rect 4493 1254 4653 1255
rect 4493 1194 4503 1254
rect 4566 1195 4653 1254
rect 4716 1195 4726 1255
rect 4814 1260 4883 1292
rect 5444 1345 5513 1363
rect 5444 1292 5450 1345
rect 5506 1292 5513 1345
rect 4814 1207 4820 1260
rect 4876 1207 4883 1260
rect 4814 1200 4883 1207
rect 5111 1256 5360 1265
rect 5111 1255 5284 1256
rect 4566 1194 4726 1195
rect 4493 1187 4726 1194
rect 5111 1195 5125 1255
rect 5188 1196 5284 1255
rect 5347 1196 5360 1256
rect 5444 1262 5513 1292
rect 5444 1209 5450 1262
rect 5506 1209 5513 1262
rect 34040 1600 34280 1700
rect 34380 1600 34760 1700
rect 34860 1600 38300 1700
rect 34040 1580 38300 1600
rect 34040 1540 38120 1580
rect 34040 1440 34280 1540
rect 34380 1440 34760 1540
rect 34860 1520 38120 1540
rect 38180 1520 38220 1580
rect 38280 1520 38300 1580
rect 34860 1480 38300 1520
rect 34860 1440 38120 1480
rect 34040 1420 38120 1440
rect 38180 1420 38220 1480
rect 38280 1420 38300 1480
rect 34040 1380 38300 1420
rect 34040 1280 34280 1380
rect 34380 1280 34760 1380
rect 34860 1280 38300 1380
rect 34040 1260 38300 1280
rect 5444 1202 5513 1209
rect 5188 1195 5360 1196
rect 5111 1188 5360 1195
rect 3220 1040 3460 1060
rect 3220 880 3260 1040
rect 3420 880 3460 1040
rect 3220 820 3460 880
rect 3220 620 3260 820
rect 3420 620 3460 820
rect 3220 540 3460 620
rect 3220 380 3260 540
rect 3420 380 3460 540
rect 3220 360 3460 380
rect 3860 1040 4100 1060
rect 3860 880 3920 1040
rect 4080 880 4100 1040
rect 3860 820 4100 880
rect 3860 620 3920 820
rect 4080 620 4100 820
rect 3860 540 4100 620
rect 3860 380 3920 540
rect 4080 380 4100 540
rect 3860 360 4100 380
rect 4480 1040 4720 1060
rect 4480 880 4520 1040
rect 4680 880 4720 1040
rect 4480 820 4720 880
rect 4480 620 4520 820
rect 4680 620 4720 820
rect 4480 540 4720 620
rect 4480 380 4520 540
rect 4680 380 4720 540
rect 4480 360 4720 380
rect 5120 1040 5360 1060
rect 5120 880 5160 1040
rect 5320 880 5360 1040
rect 5120 820 5360 880
rect 5120 620 5160 820
rect 5320 620 5360 820
rect 5120 540 5360 620
rect 5120 380 5160 540
rect 5320 380 5360 540
rect 5120 360 5360 380
rect -320 -460 6820 -440
rect -320 -520 -300 -460
rect -240 -520 -200 -460
rect -140 -480 6820 -460
rect -140 -520 1760 -480
rect -320 -560 1760 -520
rect -320 -620 -300 -560
rect -240 -620 -200 -560
rect -140 -600 1760 -560
rect 1880 -600 1980 -480
rect 2100 -600 2200 -480
rect 2320 -600 2560 -480
rect 2680 -600 2780 -480
rect 2920 -600 3000 -480
rect 3120 -600 3200 -480
rect 3340 -600 3420 -480
rect 3540 -600 3820 -480
rect 3940 -600 4020 -480
rect 4140 -600 4220 -480
rect 4340 -600 4440 -480
rect 4560 -600 4640 -480
rect 4760 -600 5040 -480
rect 5160 -600 5240 -480
rect 5360 -600 5460 -480
rect 5580 -600 5680 -480
rect 5800 -600 5880 -480
rect 6000 -600 6280 -480
rect 6400 -600 6480 -480
rect 6600 -600 6680 -480
rect 6800 -600 6820 -480
rect -140 -620 6820 -600
rect -320 -640 6820 -620
rect 37100 -1100 37800 1260
rect 32400 -1140 37800 -1100
rect 32400 -1300 33320 -1140
rect 33480 -1300 34020 -1140
rect 34180 -1300 34620 -1140
rect 34780 -1300 35220 -1140
rect 35380 -1300 35820 -1140
rect 35980 -1300 37800 -1140
rect 32400 -1380 37800 -1300
rect 32400 -1540 33320 -1380
rect 33480 -1540 34020 -1380
rect 34180 -1540 34620 -1380
rect 34780 -1540 35220 -1380
rect 35380 -1540 35820 -1380
rect 35980 -1540 37800 -1380
rect 32400 -1620 37800 -1540
rect 32400 -1780 33320 -1620
rect 33480 -1780 34020 -1620
rect 34180 -1780 34620 -1620
rect 34780 -1780 35220 -1620
rect 35380 -1780 35820 -1620
rect 35980 -1780 37800 -1620
rect 32400 -1800 37800 -1780
<< via2 >>
rect 2400 4380 2560 4540
rect 2400 4120 2560 4300
rect 2400 3880 2560 4040
rect 3640 4380 3800 4540
rect 3640 4120 3800 4300
rect 3640 3880 3800 4040
rect 4860 4380 5020 4540
rect 4860 4120 5020 4300
rect 4860 3880 5020 4040
rect 6100 4380 6260 4540
rect 6100 4120 6260 4300
rect 6100 3880 6260 4040
rect 3280 2120 3440 2280
rect 3480 2120 3640 2280
rect 3680 2120 3840 2280
rect 3880 2120 4040 2280
rect 4080 2120 4240 2280
rect 4280 2120 4440 2280
rect 4480 2120 4640 2280
rect 4680 2120 4840 2280
rect 4880 2120 5040 2280
rect 5080 2120 5240 2280
rect 34040 2140 34140 2240
rect 34040 1960 34140 2060
rect 34040 1800 34140 1900
rect 34520 2140 34620 2240
rect 34520 1960 34620 2060
rect 34520 1800 34620 1900
rect 35000 2140 35100 2240
rect 35000 1960 35100 2060
rect 35000 1800 35100 1900
rect 3236 1195 3299 1255
rect 3388 1196 3451 1256
rect 3872 1194 3935 1254
rect 4021 1195 4084 1255
rect 4503 1194 4566 1254
rect 4653 1195 4716 1255
rect 5125 1195 5188 1255
rect 5284 1196 5347 1256
rect 3260 880 3420 1040
rect 3260 620 3420 820
rect 3260 380 3420 540
rect 3920 880 4080 1040
rect 3920 620 4080 820
rect 3920 380 4080 540
rect 4520 880 4680 1040
rect 4520 620 4680 820
rect 4520 380 4680 540
rect 5160 880 5320 1040
rect 5160 620 5320 820
rect 5160 380 5320 540
<< metal3 >>
rect 30004 4682 30407 4685
rect 30987 4682 31916 5378
rect 30004 4674 31916 4682
rect 1200 4540 8660 4560
rect 1200 4380 2400 4540
rect 2560 4380 3640 4540
rect 3800 4380 4860 4540
rect 5020 4380 6100 4540
rect 6260 4460 8660 4540
rect 6260 4380 7540 4460
rect 1200 4300 7540 4380
rect 1200 4120 2400 4300
rect 2560 4120 3640 4300
rect 3800 4120 4860 4300
rect 5020 4120 6100 4300
rect 6260 4120 7540 4300
rect 1200 4040 7540 4120
rect 1200 3880 2400 4040
rect 2560 3880 3640 4040
rect 3800 3880 4860 4040
rect 5020 3880 6100 4040
rect 6260 3880 7540 4040
rect 1200 3860 7540 3880
rect 7500 3480 7540 3860
rect 8620 3480 8660 4460
rect 8982 3711 31916 4674
rect 8982 3703 30331 3711
rect 7500 3440 8660 3480
rect 7500 2460 7540 3440
rect 8620 2460 8660 3440
rect 7500 2420 8660 2460
rect 3260 2280 5320 2300
rect 3260 2120 3280 2280
rect 3440 2120 3480 2280
rect 3640 2120 3680 2280
rect 3840 2120 3880 2280
rect 4040 2120 4080 2280
rect 4240 2120 4280 2280
rect 4440 2120 4480 2280
rect 4640 2120 4680 2280
rect 4840 2120 4880 2280
rect 5040 2120 5080 2280
rect 5240 2120 5320 2280
rect 3260 2100 5320 2120
rect 3308 1267 3379 2100
rect 3228 1263 3460 1267
rect 3227 1256 3460 1263
rect 3945 1261 4016 2100
rect 4572 1264 4643 2100
rect 5203 1265 5274 2100
rect 7500 1440 7540 2420
rect 8620 1440 8660 2420
rect 30449 3520 30881 3595
rect 30449 3440 30480 3520
rect 30560 3440 30620 3520
rect 30720 3440 30780 3520
rect 30860 3440 30881 3520
rect 30449 3400 30881 3440
rect 30449 3320 30480 3400
rect 30560 3320 30620 3400
rect 30720 3320 30780 3400
rect 30860 3320 30881 3400
rect 30449 3280 30881 3320
rect 30449 3200 30480 3280
rect 30560 3200 30620 3280
rect 30720 3200 30780 3280
rect 30860 3200 30881 3280
rect 30449 3160 30881 3200
rect 30449 3080 30480 3160
rect 30560 3080 30620 3160
rect 30720 3080 30780 3160
rect 30860 3080 30881 3160
rect 30449 3040 30881 3080
rect 30449 2960 30480 3040
rect 30560 2960 30620 3040
rect 30720 2960 30780 3040
rect 30860 2960 30881 3040
rect 30449 2920 30881 2960
rect 30449 2840 30480 2920
rect 30560 2840 30620 2920
rect 30720 2840 30780 2920
rect 30860 2840 30881 2920
rect 30449 2800 30881 2840
rect 30449 2720 30480 2800
rect 30560 2720 30620 2800
rect 30720 2720 30780 2800
rect 30860 2720 30881 2800
rect 30449 2680 30881 2720
rect 30449 2600 30480 2680
rect 30560 2600 30620 2680
rect 30720 2600 30780 2680
rect 30860 2600 30881 2680
rect 30449 2560 30881 2600
rect 30449 2480 30480 2560
rect 30560 2480 30620 2560
rect 30720 2480 30780 2560
rect 30860 2480 30881 2560
rect 30449 2440 30881 2480
rect 30449 2360 30480 2440
rect 30560 2360 30620 2440
rect 30720 2360 30780 2440
rect 30860 2360 30881 2440
rect 30449 2325 30881 2360
rect 7500 1380 8660 1440
rect 4494 1261 4724 1264
rect 3862 1260 4092 1261
rect 3227 1255 3388 1256
rect 3227 1195 3236 1255
rect 3299 1196 3388 1255
rect 3451 1196 3460 1256
rect 3299 1195 3460 1196
rect 3227 1189 3460 1195
rect 3860 1255 4093 1260
rect 3860 1254 4021 1255
rect 3860 1194 3872 1254
rect 3935 1195 4021 1254
rect 4084 1195 4093 1255
rect 3935 1194 4093 1195
rect 3860 1186 4093 1194
rect 4493 1255 4726 1261
rect 4493 1254 4653 1255
rect 4493 1194 4503 1254
rect 4566 1195 4653 1254
rect 4716 1195 4726 1255
rect 4566 1194 4726 1195
rect 4493 1187 4726 1194
rect 5111 1256 5360 1265
rect 5111 1255 5284 1256
rect 5111 1195 5125 1255
rect 5188 1196 5284 1255
rect 5347 1196 5360 1256
rect 5188 1195 5360 1196
rect 5111 1188 5360 1195
rect 7500 1060 7540 1380
rect 1200 1040 7540 1060
rect 1200 880 3260 1040
rect 3420 880 3920 1040
rect 4080 880 4520 1040
rect 4680 880 5160 1040
rect 5320 880 7540 1040
rect 1200 820 7540 880
rect 1200 620 3260 820
rect 3420 620 3920 820
rect 4080 620 4520 820
rect 4680 620 5160 820
rect 5320 620 7540 820
rect 1200 540 7540 620
rect 1200 380 3260 540
rect 3420 380 3920 540
rect 4080 380 4520 540
rect 4680 380 5160 540
rect 5320 400 7540 540
rect 8620 400 8660 1380
rect 5320 380 8660 400
rect 1200 360 8660 380
rect 30987 2260 31916 3711
rect 30987 2240 35520 2260
rect 30987 2140 34040 2240
rect 34140 2140 34520 2240
rect 34620 2140 35000 2240
rect 35100 2140 35520 2240
rect 30987 2060 35520 2140
rect 30987 1960 34040 2060
rect 34140 1960 34520 2060
rect 34620 1960 35000 2060
rect 35100 1960 35520 2060
rect 30987 1900 35520 1960
rect 30987 1800 34040 1900
rect 34140 1800 34520 1900
rect 34620 1800 35000 1900
rect 35100 1800 35520 1900
rect 30987 1780 35520 1800
rect 30050 -941 30357 -939
rect 30987 -941 31916 1780
rect 30050 -944 31916 -941
rect 8982 -1912 31916 -944
rect 8982 -1915 30331 -1912
rect 30987 -2322 31916 -1912
<< via3 >>
rect 7540 3480 8620 4460
rect 7540 2460 8620 3440
rect 7540 1440 8620 2420
rect 30480 3440 30560 3520
rect 30620 3440 30720 3520
rect 30780 3440 30860 3520
rect 30480 3320 30560 3400
rect 30620 3320 30720 3400
rect 30780 3320 30860 3400
rect 30480 3200 30560 3280
rect 30620 3200 30720 3280
rect 30780 3200 30860 3280
rect 30480 3080 30560 3160
rect 30620 3080 30720 3160
rect 30780 3080 30860 3160
rect 30480 2960 30560 3040
rect 30620 2960 30720 3040
rect 30780 2960 30860 3040
rect 30480 2840 30560 2920
rect 30620 2840 30720 2920
rect 30780 2840 30860 2920
rect 30480 2720 30560 2800
rect 30620 2720 30720 2800
rect 30780 2720 30860 2800
rect 30480 2600 30560 2680
rect 30620 2600 30720 2680
rect 30780 2600 30860 2680
rect 30480 2480 30560 2560
rect 30620 2480 30720 2560
rect 30780 2480 30860 2560
rect 30480 2360 30560 2440
rect 30620 2360 30720 2440
rect 30780 2360 30860 2440
rect 7540 400 8620 1380
<< metal4 >>
rect 7485 6993 8668 7002
rect 7477 6892 30309 6993
rect 7485 4460 8668 6892
rect 7485 3480 7540 4460
rect 8620 4216 8668 4460
rect 8620 4111 9298 4216
rect 8620 3480 8668 4111
rect 30234 4107 30744 4218
rect 30651 3600 30744 4107
rect 7485 3440 8668 3480
rect 7485 2460 7540 3440
rect 8620 2460 8668 3440
rect 7485 2420 8668 2460
rect 7485 1440 7540 2420
rect 8620 1440 8668 2420
rect 7485 1381 8668 1440
rect 30440 3595 30880 3600
rect 30440 3520 30881 3595
rect 30440 3440 30480 3520
rect 30560 3440 30620 3520
rect 30720 3440 30780 3520
rect 30860 3440 30881 3520
rect 30440 3400 30881 3440
rect 30440 3320 30480 3400
rect 30560 3320 30620 3400
rect 30720 3320 30780 3400
rect 30860 3320 30881 3400
rect 30440 3280 30881 3320
rect 30440 3200 30480 3280
rect 30560 3200 30620 3280
rect 30720 3200 30780 3280
rect 30860 3200 30881 3280
rect 30440 3160 30881 3200
rect 30440 3080 30480 3160
rect 30560 3080 30620 3160
rect 30720 3080 30780 3160
rect 30860 3080 30881 3160
rect 30440 3040 30881 3080
rect 30440 2960 30480 3040
rect 30560 2960 30620 3040
rect 30720 2960 30780 3040
rect 30860 2960 30881 3040
rect 30440 2920 30881 2960
rect 30440 2840 30480 2920
rect 30560 2840 30620 2920
rect 30720 2840 30780 2920
rect 30860 2840 30881 2920
rect 30440 2800 30881 2840
rect 30440 2720 30480 2800
rect 30560 2720 30620 2800
rect 30720 2720 30780 2800
rect 30860 2720 30881 2800
rect 30440 2680 30881 2720
rect 30440 2600 30480 2680
rect 30560 2600 30620 2680
rect 30720 2600 30780 2680
rect 30860 2600 30881 2680
rect 30440 2560 30881 2600
rect 30440 2480 30480 2560
rect 30560 2480 30620 2560
rect 30720 2480 30780 2560
rect 30860 2480 30881 2560
rect 30440 2440 30881 2480
rect 30440 2360 30480 2440
rect 30560 2360 30620 2440
rect 30720 2360 30780 2440
rect 30860 2360 30881 2440
rect 30440 2325 30881 2360
rect 7485 1380 30320 1381
rect 7485 400 7540 1380
rect 8620 1281 30320 1380
rect 8620 400 8668 1281
rect 7485 -1401 8668 400
rect 30440 -1220 30880 2325
rect 7485 -1506 9367 -1401
rect 30654 -1403 30743 -1220
rect 30186 -1498 30748 -1403
rect 7485 -3876 8668 -1506
use sky130_fd_pr__cap_mim_m3_1_RF494X  XC1
timestamp 1769436194
transform 0 -1 19666 1 0 1500
box -5492 -10640 5492 10640
use sky130_fd_pr__pfet_g5v0d10v5_4KVG5X  XM1
timestamp 1769412267
transform 1 0 4329 0 1 4204
box -2559 -1004 2559 1042
use sky130_fd_pr__nfet_g5v0d10v5_EP6D69  XM3
timestamp 1769412267
transform 1 0 4293 0 1 728
box -1293 -528 1293 528
use sky130_fd_pr__nfet_g5v0d10v5_H6999P  XM5
timestamp 1769412267
transform 1 0 4293 0 1 -1393
box -2493 -807 2493 807
use sky130_fd_pr__pfet_g5v0d10v5_ZC39X7  XM7
timestamp 1769412267
transform 1 0 34649 0 1 4038
box -2559 -1064 2559 1102
use sky130_fd_pr__nfet_g5v0d10v5_BYSCSD  XM8
timestamp 1769412267
transform 1 0 34666 0 1 -1387
box -1261 -807 1261 807
use sky130_fd_pr__pfet_g5v0d10v5_AKJWHE  XM9
timestamp 1769417084
transform 1 0 34571 0 1 1664
box -571 -564 571 602
<< labels >>
flabel metal1 1080 6720 1280 6920 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1180 -2700 1380 -2500 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 -320 -640 -120 -440 0 FreeSans 256 0 0 0 IBIAS
port 4 nsew
flabel metal1 -320 2100 -120 2300 0 FreeSans 256 0 0 0 VN
port 3 nsew
flabel metal1 -320 1700 -120 1900 0 FreeSans 256 0 0 0 VP
port 2 nsew
flabel metal1 38100 1400 38300 1600 0 FreeSans 256 0 0 0 OUT
port 1 nsew
<< end >>
