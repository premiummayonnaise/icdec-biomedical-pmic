magic
tech sky130A
magscale 1 2
timestamp 1770083657
<< error_p >>
rect -2867 1038 2867 1042
rect -2867 -970 -2837 1038
rect -2801 972 2801 976
rect -2801 -904 -2771 972
rect 2771 -904 2801 972
rect 2837 -970 2867 1038
<< nwell >>
rect -2837 -1004 2837 1038
<< mvpmos >>
rect -2743 -904 -2493 976
rect -2435 -904 -2185 976
rect -2127 -904 -1877 976
rect -1819 -904 -1569 976
rect -1511 -904 -1261 976
rect -1203 -904 -953 976
rect -895 -904 -645 976
rect -587 -904 -337 976
rect -279 -904 -29 976
rect 29 -904 279 976
rect 337 -904 587 976
rect 645 -904 895 976
rect 953 -904 1203 976
rect 1261 -904 1511 976
rect 1569 -904 1819 976
rect 1877 -904 2127 976
rect 2185 -904 2435 976
rect 2493 -904 2743 976
<< mvpdiff >>
rect -2801 937 -2743 976
rect -2801 903 -2789 937
rect -2755 903 -2743 937
rect -2801 869 -2743 903
rect -2801 835 -2789 869
rect -2755 835 -2743 869
rect -2801 801 -2743 835
rect -2801 767 -2789 801
rect -2755 767 -2743 801
rect -2801 733 -2743 767
rect -2801 699 -2789 733
rect -2755 699 -2743 733
rect -2801 665 -2743 699
rect -2801 631 -2789 665
rect -2755 631 -2743 665
rect -2801 597 -2743 631
rect -2801 563 -2789 597
rect -2755 563 -2743 597
rect -2801 529 -2743 563
rect -2801 495 -2789 529
rect -2755 495 -2743 529
rect -2801 461 -2743 495
rect -2801 427 -2789 461
rect -2755 427 -2743 461
rect -2801 393 -2743 427
rect -2801 359 -2789 393
rect -2755 359 -2743 393
rect -2801 325 -2743 359
rect -2801 291 -2789 325
rect -2755 291 -2743 325
rect -2801 257 -2743 291
rect -2801 223 -2789 257
rect -2755 223 -2743 257
rect -2801 189 -2743 223
rect -2801 155 -2789 189
rect -2755 155 -2743 189
rect -2801 121 -2743 155
rect -2801 87 -2789 121
rect -2755 87 -2743 121
rect -2801 53 -2743 87
rect -2801 19 -2789 53
rect -2755 19 -2743 53
rect -2801 -15 -2743 19
rect -2801 -49 -2789 -15
rect -2755 -49 -2743 -15
rect -2801 -83 -2743 -49
rect -2801 -117 -2789 -83
rect -2755 -117 -2743 -83
rect -2801 -151 -2743 -117
rect -2801 -185 -2789 -151
rect -2755 -185 -2743 -151
rect -2801 -219 -2743 -185
rect -2801 -253 -2789 -219
rect -2755 -253 -2743 -219
rect -2801 -287 -2743 -253
rect -2801 -321 -2789 -287
rect -2755 -321 -2743 -287
rect -2801 -355 -2743 -321
rect -2801 -389 -2789 -355
rect -2755 -389 -2743 -355
rect -2801 -423 -2743 -389
rect -2801 -457 -2789 -423
rect -2755 -457 -2743 -423
rect -2801 -491 -2743 -457
rect -2801 -525 -2789 -491
rect -2755 -525 -2743 -491
rect -2801 -559 -2743 -525
rect -2801 -593 -2789 -559
rect -2755 -593 -2743 -559
rect -2801 -627 -2743 -593
rect -2801 -661 -2789 -627
rect -2755 -661 -2743 -627
rect -2801 -695 -2743 -661
rect -2801 -729 -2789 -695
rect -2755 -729 -2743 -695
rect -2801 -763 -2743 -729
rect -2801 -797 -2789 -763
rect -2755 -797 -2743 -763
rect -2801 -831 -2743 -797
rect -2801 -865 -2789 -831
rect -2755 -865 -2743 -831
rect -2801 -904 -2743 -865
rect -2493 937 -2435 976
rect -2493 903 -2481 937
rect -2447 903 -2435 937
rect -2493 869 -2435 903
rect -2493 835 -2481 869
rect -2447 835 -2435 869
rect -2493 801 -2435 835
rect -2493 767 -2481 801
rect -2447 767 -2435 801
rect -2493 733 -2435 767
rect -2493 699 -2481 733
rect -2447 699 -2435 733
rect -2493 665 -2435 699
rect -2493 631 -2481 665
rect -2447 631 -2435 665
rect -2493 597 -2435 631
rect -2493 563 -2481 597
rect -2447 563 -2435 597
rect -2493 529 -2435 563
rect -2493 495 -2481 529
rect -2447 495 -2435 529
rect -2493 461 -2435 495
rect -2493 427 -2481 461
rect -2447 427 -2435 461
rect -2493 393 -2435 427
rect -2493 359 -2481 393
rect -2447 359 -2435 393
rect -2493 325 -2435 359
rect -2493 291 -2481 325
rect -2447 291 -2435 325
rect -2493 257 -2435 291
rect -2493 223 -2481 257
rect -2447 223 -2435 257
rect -2493 189 -2435 223
rect -2493 155 -2481 189
rect -2447 155 -2435 189
rect -2493 121 -2435 155
rect -2493 87 -2481 121
rect -2447 87 -2435 121
rect -2493 53 -2435 87
rect -2493 19 -2481 53
rect -2447 19 -2435 53
rect -2493 -15 -2435 19
rect -2493 -49 -2481 -15
rect -2447 -49 -2435 -15
rect -2493 -83 -2435 -49
rect -2493 -117 -2481 -83
rect -2447 -117 -2435 -83
rect -2493 -151 -2435 -117
rect -2493 -185 -2481 -151
rect -2447 -185 -2435 -151
rect -2493 -219 -2435 -185
rect -2493 -253 -2481 -219
rect -2447 -253 -2435 -219
rect -2493 -287 -2435 -253
rect -2493 -321 -2481 -287
rect -2447 -321 -2435 -287
rect -2493 -355 -2435 -321
rect -2493 -389 -2481 -355
rect -2447 -389 -2435 -355
rect -2493 -423 -2435 -389
rect -2493 -457 -2481 -423
rect -2447 -457 -2435 -423
rect -2493 -491 -2435 -457
rect -2493 -525 -2481 -491
rect -2447 -525 -2435 -491
rect -2493 -559 -2435 -525
rect -2493 -593 -2481 -559
rect -2447 -593 -2435 -559
rect -2493 -627 -2435 -593
rect -2493 -661 -2481 -627
rect -2447 -661 -2435 -627
rect -2493 -695 -2435 -661
rect -2493 -729 -2481 -695
rect -2447 -729 -2435 -695
rect -2493 -763 -2435 -729
rect -2493 -797 -2481 -763
rect -2447 -797 -2435 -763
rect -2493 -831 -2435 -797
rect -2493 -865 -2481 -831
rect -2447 -865 -2435 -831
rect -2493 -904 -2435 -865
rect -2185 937 -2127 976
rect -2185 903 -2173 937
rect -2139 903 -2127 937
rect -2185 869 -2127 903
rect -2185 835 -2173 869
rect -2139 835 -2127 869
rect -2185 801 -2127 835
rect -2185 767 -2173 801
rect -2139 767 -2127 801
rect -2185 733 -2127 767
rect -2185 699 -2173 733
rect -2139 699 -2127 733
rect -2185 665 -2127 699
rect -2185 631 -2173 665
rect -2139 631 -2127 665
rect -2185 597 -2127 631
rect -2185 563 -2173 597
rect -2139 563 -2127 597
rect -2185 529 -2127 563
rect -2185 495 -2173 529
rect -2139 495 -2127 529
rect -2185 461 -2127 495
rect -2185 427 -2173 461
rect -2139 427 -2127 461
rect -2185 393 -2127 427
rect -2185 359 -2173 393
rect -2139 359 -2127 393
rect -2185 325 -2127 359
rect -2185 291 -2173 325
rect -2139 291 -2127 325
rect -2185 257 -2127 291
rect -2185 223 -2173 257
rect -2139 223 -2127 257
rect -2185 189 -2127 223
rect -2185 155 -2173 189
rect -2139 155 -2127 189
rect -2185 121 -2127 155
rect -2185 87 -2173 121
rect -2139 87 -2127 121
rect -2185 53 -2127 87
rect -2185 19 -2173 53
rect -2139 19 -2127 53
rect -2185 -15 -2127 19
rect -2185 -49 -2173 -15
rect -2139 -49 -2127 -15
rect -2185 -83 -2127 -49
rect -2185 -117 -2173 -83
rect -2139 -117 -2127 -83
rect -2185 -151 -2127 -117
rect -2185 -185 -2173 -151
rect -2139 -185 -2127 -151
rect -2185 -219 -2127 -185
rect -2185 -253 -2173 -219
rect -2139 -253 -2127 -219
rect -2185 -287 -2127 -253
rect -2185 -321 -2173 -287
rect -2139 -321 -2127 -287
rect -2185 -355 -2127 -321
rect -2185 -389 -2173 -355
rect -2139 -389 -2127 -355
rect -2185 -423 -2127 -389
rect -2185 -457 -2173 -423
rect -2139 -457 -2127 -423
rect -2185 -491 -2127 -457
rect -2185 -525 -2173 -491
rect -2139 -525 -2127 -491
rect -2185 -559 -2127 -525
rect -2185 -593 -2173 -559
rect -2139 -593 -2127 -559
rect -2185 -627 -2127 -593
rect -2185 -661 -2173 -627
rect -2139 -661 -2127 -627
rect -2185 -695 -2127 -661
rect -2185 -729 -2173 -695
rect -2139 -729 -2127 -695
rect -2185 -763 -2127 -729
rect -2185 -797 -2173 -763
rect -2139 -797 -2127 -763
rect -2185 -831 -2127 -797
rect -2185 -865 -2173 -831
rect -2139 -865 -2127 -831
rect -2185 -904 -2127 -865
rect -1877 937 -1819 976
rect -1877 903 -1865 937
rect -1831 903 -1819 937
rect -1877 869 -1819 903
rect -1877 835 -1865 869
rect -1831 835 -1819 869
rect -1877 801 -1819 835
rect -1877 767 -1865 801
rect -1831 767 -1819 801
rect -1877 733 -1819 767
rect -1877 699 -1865 733
rect -1831 699 -1819 733
rect -1877 665 -1819 699
rect -1877 631 -1865 665
rect -1831 631 -1819 665
rect -1877 597 -1819 631
rect -1877 563 -1865 597
rect -1831 563 -1819 597
rect -1877 529 -1819 563
rect -1877 495 -1865 529
rect -1831 495 -1819 529
rect -1877 461 -1819 495
rect -1877 427 -1865 461
rect -1831 427 -1819 461
rect -1877 393 -1819 427
rect -1877 359 -1865 393
rect -1831 359 -1819 393
rect -1877 325 -1819 359
rect -1877 291 -1865 325
rect -1831 291 -1819 325
rect -1877 257 -1819 291
rect -1877 223 -1865 257
rect -1831 223 -1819 257
rect -1877 189 -1819 223
rect -1877 155 -1865 189
rect -1831 155 -1819 189
rect -1877 121 -1819 155
rect -1877 87 -1865 121
rect -1831 87 -1819 121
rect -1877 53 -1819 87
rect -1877 19 -1865 53
rect -1831 19 -1819 53
rect -1877 -15 -1819 19
rect -1877 -49 -1865 -15
rect -1831 -49 -1819 -15
rect -1877 -83 -1819 -49
rect -1877 -117 -1865 -83
rect -1831 -117 -1819 -83
rect -1877 -151 -1819 -117
rect -1877 -185 -1865 -151
rect -1831 -185 -1819 -151
rect -1877 -219 -1819 -185
rect -1877 -253 -1865 -219
rect -1831 -253 -1819 -219
rect -1877 -287 -1819 -253
rect -1877 -321 -1865 -287
rect -1831 -321 -1819 -287
rect -1877 -355 -1819 -321
rect -1877 -389 -1865 -355
rect -1831 -389 -1819 -355
rect -1877 -423 -1819 -389
rect -1877 -457 -1865 -423
rect -1831 -457 -1819 -423
rect -1877 -491 -1819 -457
rect -1877 -525 -1865 -491
rect -1831 -525 -1819 -491
rect -1877 -559 -1819 -525
rect -1877 -593 -1865 -559
rect -1831 -593 -1819 -559
rect -1877 -627 -1819 -593
rect -1877 -661 -1865 -627
rect -1831 -661 -1819 -627
rect -1877 -695 -1819 -661
rect -1877 -729 -1865 -695
rect -1831 -729 -1819 -695
rect -1877 -763 -1819 -729
rect -1877 -797 -1865 -763
rect -1831 -797 -1819 -763
rect -1877 -831 -1819 -797
rect -1877 -865 -1865 -831
rect -1831 -865 -1819 -831
rect -1877 -904 -1819 -865
rect -1569 937 -1511 976
rect -1569 903 -1557 937
rect -1523 903 -1511 937
rect -1569 869 -1511 903
rect -1569 835 -1557 869
rect -1523 835 -1511 869
rect -1569 801 -1511 835
rect -1569 767 -1557 801
rect -1523 767 -1511 801
rect -1569 733 -1511 767
rect -1569 699 -1557 733
rect -1523 699 -1511 733
rect -1569 665 -1511 699
rect -1569 631 -1557 665
rect -1523 631 -1511 665
rect -1569 597 -1511 631
rect -1569 563 -1557 597
rect -1523 563 -1511 597
rect -1569 529 -1511 563
rect -1569 495 -1557 529
rect -1523 495 -1511 529
rect -1569 461 -1511 495
rect -1569 427 -1557 461
rect -1523 427 -1511 461
rect -1569 393 -1511 427
rect -1569 359 -1557 393
rect -1523 359 -1511 393
rect -1569 325 -1511 359
rect -1569 291 -1557 325
rect -1523 291 -1511 325
rect -1569 257 -1511 291
rect -1569 223 -1557 257
rect -1523 223 -1511 257
rect -1569 189 -1511 223
rect -1569 155 -1557 189
rect -1523 155 -1511 189
rect -1569 121 -1511 155
rect -1569 87 -1557 121
rect -1523 87 -1511 121
rect -1569 53 -1511 87
rect -1569 19 -1557 53
rect -1523 19 -1511 53
rect -1569 -15 -1511 19
rect -1569 -49 -1557 -15
rect -1523 -49 -1511 -15
rect -1569 -83 -1511 -49
rect -1569 -117 -1557 -83
rect -1523 -117 -1511 -83
rect -1569 -151 -1511 -117
rect -1569 -185 -1557 -151
rect -1523 -185 -1511 -151
rect -1569 -219 -1511 -185
rect -1569 -253 -1557 -219
rect -1523 -253 -1511 -219
rect -1569 -287 -1511 -253
rect -1569 -321 -1557 -287
rect -1523 -321 -1511 -287
rect -1569 -355 -1511 -321
rect -1569 -389 -1557 -355
rect -1523 -389 -1511 -355
rect -1569 -423 -1511 -389
rect -1569 -457 -1557 -423
rect -1523 -457 -1511 -423
rect -1569 -491 -1511 -457
rect -1569 -525 -1557 -491
rect -1523 -525 -1511 -491
rect -1569 -559 -1511 -525
rect -1569 -593 -1557 -559
rect -1523 -593 -1511 -559
rect -1569 -627 -1511 -593
rect -1569 -661 -1557 -627
rect -1523 -661 -1511 -627
rect -1569 -695 -1511 -661
rect -1569 -729 -1557 -695
rect -1523 -729 -1511 -695
rect -1569 -763 -1511 -729
rect -1569 -797 -1557 -763
rect -1523 -797 -1511 -763
rect -1569 -831 -1511 -797
rect -1569 -865 -1557 -831
rect -1523 -865 -1511 -831
rect -1569 -904 -1511 -865
rect -1261 937 -1203 976
rect -1261 903 -1249 937
rect -1215 903 -1203 937
rect -1261 869 -1203 903
rect -1261 835 -1249 869
rect -1215 835 -1203 869
rect -1261 801 -1203 835
rect -1261 767 -1249 801
rect -1215 767 -1203 801
rect -1261 733 -1203 767
rect -1261 699 -1249 733
rect -1215 699 -1203 733
rect -1261 665 -1203 699
rect -1261 631 -1249 665
rect -1215 631 -1203 665
rect -1261 597 -1203 631
rect -1261 563 -1249 597
rect -1215 563 -1203 597
rect -1261 529 -1203 563
rect -1261 495 -1249 529
rect -1215 495 -1203 529
rect -1261 461 -1203 495
rect -1261 427 -1249 461
rect -1215 427 -1203 461
rect -1261 393 -1203 427
rect -1261 359 -1249 393
rect -1215 359 -1203 393
rect -1261 325 -1203 359
rect -1261 291 -1249 325
rect -1215 291 -1203 325
rect -1261 257 -1203 291
rect -1261 223 -1249 257
rect -1215 223 -1203 257
rect -1261 189 -1203 223
rect -1261 155 -1249 189
rect -1215 155 -1203 189
rect -1261 121 -1203 155
rect -1261 87 -1249 121
rect -1215 87 -1203 121
rect -1261 53 -1203 87
rect -1261 19 -1249 53
rect -1215 19 -1203 53
rect -1261 -15 -1203 19
rect -1261 -49 -1249 -15
rect -1215 -49 -1203 -15
rect -1261 -83 -1203 -49
rect -1261 -117 -1249 -83
rect -1215 -117 -1203 -83
rect -1261 -151 -1203 -117
rect -1261 -185 -1249 -151
rect -1215 -185 -1203 -151
rect -1261 -219 -1203 -185
rect -1261 -253 -1249 -219
rect -1215 -253 -1203 -219
rect -1261 -287 -1203 -253
rect -1261 -321 -1249 -287
rect -1215 -321 -1203 -287
rect -1261 -355 -1203 -321
rect -1261 -389 -1249 -355
rect -1215 -389 -1203 -355
rect -1261 -423 -1203 -389
rect -1261 -457 -1249 -423
rect -1215 -457 -1203 -423
rect -1261 -491 -1203 -457
rect -1261 -525 -1249 -491
rect -1215 -525 -1203 -491
rect -1261 -559 -1203 -525
rect -1261 -593 -1249 -559
rect -1215 -593 -1203 -559
rect -1261 -627 -1203 -593
rect -1261 -661 -1249 -627
rect -1215 -661 -1203 -627
rect -1261 -695 -1203 -661
rect -1261 -729 -1249 -695
rect -1215 -729 -1203 -695
rect -1261 -763 -1203 -729
rect -1261 -797 -1249 -763
rect -1215 -797 -1203 -763
rect -1261 -831 -1203 -797
rect -1261 -865 -1249 -831
rect -1215 -865 -1203 -831
rect -1261 -904 -1203 -865
rect -953 937 -895 976
rect -953 903 -941 937
rect -907 903 -895 937
rect -953 869 -895 903
rect -953 835 -941 869
rect -907 835 -895 869
rect -953 801 -895 835
rect -953 767 -941 801
rect -907 767 -895 801
rect -953 733 -895 767
rect -953 699 -941 733
rect -907 699 -895 733
rect -953 665 -895 699
rect -953 631 -941 665
rect -907 631 -895 665
rect -953 597 -895 631
rect -953 563 -941 597
rect -907 563 -895 597
rect -953 529 -895 563
rect -953 495 -941 529
rect -907 495 -895 529
rect -953 461 -895 495
rect -953 427 -941 461
rect -907 427 -895 461
rect -953 393 -895 427
rect -953 359 -941 393
rect -907 359 -895 393
rect -953 325 -895 359
rect -953 291 -941 325
rect -907 291 -895 325
rect -953 257 -895 291
rect -953 223 -941 257
rect -907 223 -895 257
rect -953 189 -895 223
rect -953 155 -941 189
rect -907 155 -895 189
rect -953 121 -895 155
rect -953 87 -941 121
rect -907 87 -895 121
rect -953 53 -895 87
rect -953 19 -941 53
rect -907 19 -895 53
rect -953 -15 -895 19
rect -953 -49 -941 -15
rect -907 -49 -895 -15
rect -953 -83 -895 -49
rect -953 -117 -941 -83
rect -907 -117 -895 -83
rect -953 -151 -895 -117
rect -953 -185 -941 -151
rect -907 -185 -895 -151
rect -953 -219 -895 -185
rect -953 -253 -941 -219
rect -907 -253 -895 -219
rect -953 -287 -895 -253
rect -953 -321 -941 -287
rect -907 -321 -895 -287
rect -953 -355 -895 -321
rect -953 -389 -941 -355
rect -907 -389 -895 -355
rect -953 -423 -895 -389
rect -953 -457 -941 -423
rect -907 -457 -895 -423
rect -953 -491 -895 -457
rect -953 -525 -941 -491
rect -907 -525 -895 -491
rect -953 -559 -895 -525
rect -953 -593 -941 -559
rect -907 -593 -895 -559
rect -953 -627 -895 -593
rect -953 -661 -941 -627
rect -907 -661 -895 -627
rect -953 -695 -895 -661
rect -953 -729 -941 -695
rect -907 -729 -895 -695
rect -953 -763 -895 -729
rect -953 -797 -941 -763
rect -907 -797 -895 -763
rect -953 -831 -895 -797
rect -953 -865 -941 -831
rect -907 -865 -895 -831
rect -953 -904 -895 -865
rect -645 937 -587 976
rect -645 903 -633 937
rect -599 903 -587 937
rect -645 869 -587 903
rect -645 835 -633 869
rect -599 835 -587 869
rect -645 801 -587 835
rect -645 767 -633 801
rect -599 767 -587 801
rect -645 733 -587 767
rect -645 699 -633 733
rect -599 699 -587 733
rect -645 665 -587 699
rect -645 631 -633 665
rect -599 631 -587 665
rect -645 597 -587 631
rect -645 563 -633 597
rect -599 563 -587 597
rect -645 529 -587 563
rect -645 495 -633 529
rect -599 495 -587 529
rect -645 461 -587 495
rect -645 427 -633 461
rect -599 427 -587 461
rect -645 393 -587 427
rect -645 359 -633 393
rect -599 359 -587 393
rect -645 325 -587 359
rect -645 291 -633 325
rect -599 291 -587 325
rect -645 257 -587 291
rect -645 223 -633 257
rect -599 223 -587 257
rect -645 189 -587 223
rect -645 155 -633 189
rect -599 155 -587 189
rect -645 121 -587 155
rect -645 87 -633 121
rect -599 87 -587 121
rect -645 53 -587 87
rect -645 19 -633 53
rect -599 19 -587 53
rect -645 -15 -587 19
rect -645 -49 -633 -15
rect -599 -49 -587 -15
rect -645 -83 -587 -49
rect -645 -117 -633 -83
rect -599 -117 -587 -83
rect -645 -151 -587 -117
rect -645 -185 -633 -151
rect -599 -185 -587 -151
rect -645 -219 -587 -185
rect -645 -253 -633 -219
rect -599 -253 -587 -219
rect -645 -287 -587 -253
rect -645 -321 -633 -287
rect -599 -321 -587 -287
rect -645 -355 -587 -321
rect -645 -389 -633 -355
rect -599 -389 -587 -355
rect -645 -423 -587 -389
rect -645 -457 -633 -423
rect -599 -457 -587 -423
rect -645 -491 -587 -457
rect -645 -525 -633 -491
rect -599 -525 -587 -491
rect -645 -559 -587 -525
rect -645 -593 -633 -559
rect -599 -593 -587 -559
rect -645 -627 -587 -593
rect -645 -661 -633 -627
rect -599 -661 -587 -627
rect -645 -695 -587 -661
rect -645 -729 -633 -695
rect -599 -729 -587 -695
rect -645 -763 -587 -729
rect -645 -797 -633 -763
rect -599 -797 -587 -763
rect -645 -831 -587 -797
rect -645 -865 -633 -831
rect -599 -865 -587 -831
rect -645 -904 -587 -865
rect -337 937 -279 976
rect -337 903 -325 937
rect -291 903 -279 937
rect -337 869 -279 903
rect -337 835 -325 869
rect -291 835 -279 869
rect -337 801 -279 835
rect -337 767 -325 801
rect -291 767 -279 801
rect -337 733 -279 767
rect -337 699 -325 733
rect -291 699 -279 733
rect -337 665 -279 699
rect -337 631 -325 665
rect -291 631 -279 665
rect -337 597 -279 631
rect -337 563 -325 597
rect -291 563 -279 597
rect -337 529 -279 563
rect -337 495 -325 529
rect -291 495 -279 529
rect -337 461 -279 495
rect -337 427 -325 461
rect -291 427 -279 461
rect -337 393 -279 427
rect -337 359 -325 393
rect -291 359 -279 393
rect -337 325 -279 359
rect -337 291 -325 325
rect -291 291 -279 325
rect -337 257 -279 291
rect -337 223 -325 257
rect -291 223 -279 257
rect -337 189 -279 223
rect -337 155 -325 189
rect -291 155 -279 189
rect -337 121 -279 155
rect -337 87 -325 121
rect -291 87 -279 121
rect -337 53 -279 87
rect -337 19 -325 53
rect -291 19 -279 53
rect -337 -15 -279 19
rect -337 -49 -325 -15
rect -291 -49 -279 -15
rect -337 -83 -279 -49
rect -337 -117 -325 -83
rect -291 -117 -279 -83
rect -337 -151 -279 -117
rect -337 -185 -325 -151
rect -291 -185 -279 -151
rect -337 -219 -279 -185
rect -337 -253 -325 -219
rect -291 -253 -279 -219
rect -337 -287 -279 -253
rect -337 -321 -325 -287
rect -291 -321 -279 -287
rect -337 -355 -279 -321
rect -337 -389 -325 -355
rect -291 -389 -279 -355
rect -337 -423 -279 -389
rect -337 -457 -325 -423
rect -291 -457 -279 -423
rect -337 -491 -279 -457
rect -337 -525 -325 -491
rect -291 -525 -279 -491
rect -337 -559 -279 -525
rect -337 -593 -325 -559
rect -291 -593 -279 -559
rect -337 -627 -279 -593
rect -337 -661 -325 -627
rect -291 -661 -279 -627
rect -337 -695 -279 -661
rect -337 -729 -325 -695
rect -291 -729 -279 -695
rect -337 -763 -279 -729
rect -337 -797 -325 -763
rect -291 -797 -279 -763
rect -337 -831 -279 -797
rect -337 -865 -325 -831
rect -291 -865 -279 -831
rect -337 -904 -279 -865
rect -29 937 29 976
rect -29 903 -17 937
rect 17 903 29 937
rect -29 869 29 903
rect -29 835 -17 869
rect 17 835 29 869
rect -29 801 29 835
rect -29 767 -17 801
rect 17 767 29 801
rect -29 733 29 767
rect -29 699 -17 733
rect 17 699 29 733
rect -29 665 29 699
rect -29 631 -17 665
rect 17 631 29 665
rect -29 597 29 631
rect -29 563 -17 597
rect 17 563 29 597
rect -29 529 29 563
rect -29 495 -17 529
rect 17 495 29 529
rect -29 461 29 495
rect -29 427 -17 461
rect 17 427 29 461
rect -29 393 29 427
rect -29 359 -17 393
rect 17 359 29 393
rect -29 325 29 359
rect -29 291 -17 325
rect 17 291 29 325
rect -29 257 29 291
rect -29 223 -17 257
rect 17 223 29 257
rect -29 189 29 223
rect -29 155 -17 189
rect 17 155 29 189
rect -29 121 29 155
rect -29 87 -17 121
rect 17 87 29 121
rect -29 53 29 87
rect -29 19 -17 53
rect 17 19 29 53
rect -29 -15 29 19
rect -29 -49 -17 -15
rect 17 -49 29 -15
rect -29 -83 29 -49
rect -29 -117 -17 -83
rect 17 -117 29 -83
rect -29 -151 29 -117
rect -29 -185 -17 -151
rect 17 -185 29 -151
rect -29 -219 29 -185
rect -29 -253 -17 -219
rect 17 -253 29 -219
rect -29 -287 29 -253
rect -29 -321 -17 -287
rect 17 -321 29 -287
rect -29 -355 29 -321
rect -29 -389 -17 -355
rect 17 -389 29 -355
rect -29 -423 29 -389
rect -29 -457 -17 -423
rect 17 -457 29 -423
rect -29 -491 29 -457
rect -29 -525 -17 -491
rect 17 -525 29 -491
rect -29 -559 29 -525
rect -29 -593 -17 -559
rect 17 -593 29 -559
rect -29 -627 29 -593
rect -29 -661 -17 -627
rect 17 -661 29 -627
rect -29 -695 29 -661
rect -29 -729 -17 -695
rect 17 -729 29 -695
rect -29 -763 29 -729
rect -29 -797 -17 -763
rect 17 -797 29 -763
rect -29 -831 29 -797
rect -29 -865 -17 -831
rect 17 -865 29 -831
rect -29 -904 29 -865
rect 279 937 337 976
rect 279 903 291 937
rect 325 903 337 937
rect 279 869 337 903
rect 279 835 291 869
rect 325 835 337 869
rect 279 801 337 835
rect 279 767 291 801
rect 325 767 337 801
rect 279 733 337 767
rect 279 699 291 733
rect 325 699 337 733
rect 279 665 337 699
rect 279 631 291 665
rect 325 631 337 665
rect 279 597 337 631
rect 279 563 291 597
rect 325 563 337 597
rect 279 529 337 563
rect 279 495 291 529
rect 325 495 337 529
rect 279 461 337 495
rect 279 427 291 461
rect 325 427 337 461
rect 279 393 337 427
rect 279 359 291 393
rect 325 359 337 393
rect 279 325 337 359
rect 279 291 291 325
rect 325 291 337 325
rect 279 257 337 291
rect 279 223 291 257
rect 325 223 337 257
rect 279 189 337 223
rect 279 155 291 189
rect 325 155 337 189
rect 279 121 337 155
rect 279 87 291 121
rect 325 87 337 121
rect 279 53 337 87
rect 279 19 291 53
rect 325 19 337 53
rect 279 -15 337 19
rect 279 -49 291 -15
rect 325 -49 337 -15
rect 279 -83 337 -49
rect 279 -117 291 -83
rect 325 -117 337 -83
rect 279 -151 337 -117
rect 279 -185 291 -151
rect 325 -185 337 -151
rect 279 -219 337 -185
rect 279 -253 291 -219
rect 325 -253 337 -219
rect 279 -287 337 -253
rect 279 -321 291 -287
rect 325 -321 337 -287
rect 279 -355 337 -321
rect 279 -389 291 -355
rect 325 -389 337 -355
rect 279 -423 337 -389
rect 279 -457 291 -423
rect 325 -457 337 -423
rect 279 -491 337 -457
rect 279 -525 291 -491
rect 325 -525 337 -491
rect 279 -559 337 -525
rect 279 -593 291 -559
rect 325 -593 337 -559
rect 279 -627 337 -593
rect 279 -661 291 -627
rect 325 -661 337 -627
rect 279 -695 337 -661
rect 279 -729 291 -695
rect 325 -729 337 -695
rect 279 -763 337 -729
rect 279 -797 291 -763
rect 325 -797 337 -763
rect 279 -831 337 -797
rect 279 -865 291 -831
rect 325 -865 337 -831
rect 279 -904 337 -865
rect 587 937 645 976
rect 587 903 599 937
rect 633 903 645 937
rect 587 869 645 903
rect 587 835 599 869
rect 633 835 645 869
rect 587 801 645 835
rect 587 767 599 801
rect 633 767 645 801
rect 587 733 645 767
rect 587 699 599 733
rect 633 699 645 733
rect 587 665 645 699
rect 587 631 599 665
rect 633 631 645 665
rect 587 597 645 631
rect 587 563 599 597
rect 633 563 645 597
rect 587 529 645 563
rect 587 495 599 529
rect 633 495 645 529
rect 587 461 645 495
rect 587 427 599 461
rect 633 427 645 461
rect 587 393 645 427
rect 587 359 599 393
rect 633 359 645 393
rect 587 325 645 359
rect 587 291 599 325
rect 633 291 645 325
rect 587 257 645 291
rect 587 223 599 257
rect 633 223 645 257
rect 587 189 645 223
rect 587 155 599 189
rect 633 155 645 189
rect 587 121 645 155
rect 587 87 599 121
rect 633 87 645 121
rect 587 53 645 87
rect 587 19 599 53
rect 633 19 645 53
rect 587 -15 645 19
rect 587 -49 599 -15
rect 633 -49 645 -15
rect 587 -83 645 -49
rect 587 -117 599 -83
rect 633 -117 645 -83
rect 587 -151 645 -117
rect 587 -185 599 -151
rect 633 -185 645 -151
rect 587 -219 645 -185
rect 587 -253 599 -219
rect 633 -253 645 -219
rect 587 -287 645 -253
rect 587 -321 599 -287
rect 633 -321 645 -287
rect 587 -355 645 -321
rect 587 -389 599 -355
rect 633 -389 645 -355
rect 587 -423 645 -389
rect 587 -457 599 -423
rect 633 -457 645 -423
rect 587 -491 645 -457
rect 587 -525 599 -491
rect 633 -525 645 -491
rect 587 -559 645 -525
rect 587 -593 599 -559
rect 633 -593 645 -559
rect 587 -627 645 -593
rect 587 -661 599 -627
rect 633 -661 645 -627
rect 587 -695 645 -661
rect 587 -729 599 -695
rect 633 -729 645 -695
rect 587 -763 645 -729
rect 587 -797 599 -763
rect 633 -797 645 -763
rect 587 -831 645 -797
rect 587 -865 599 -831
rect 633 -865 645 -831
rect 587 -904 645 -865
rect 895 937 953 976
rect 895 903 907 937
rect 941 903 953 937
rect 895 869 953 903
rect 895 835 907 869
rect 941 835 953 869
rect 895 801 953 835
rect 895 767 907 801
rect 941 767 953 801
rect 895 733 953 767
rect 895 699 907 733
rect 941 699 953 733
rect 895 665 953 699
rect 895 631 907 665
rect 941 631 953 665
rect 895 597 953 631
rect 895 563 907 597
rect 941 563 953 597
rect 895 529 953 563
rect 895 495 907 529
rect 941 495 953 529
rect 895 461 953 495
rect 895 427 907 461
rect 941 427 953 461
rect 895 393 953 427
rect 895 359 907 393
rect 941 359 953 393
rect 895 325 953 359
rect 895 291 907 325
rect 941 291 953 325
rect 895 257 953 291
rect 895 223 907 257
rect 941 223 953 257
rect 895 189 953 223
rect 895 155 907 189
rect 941 155 953 189
rect 895 121 953 155
rect 895 87 907 121
rect 941 87 953 121
rect 895 53 953 87
rect 895 19 907 53
rect 941 19 953 53
rect 895 -15 953 19
rect 895 -49 907 -15
rect 941 -49 953 -15
rect 895 -83 953 -49
rect 895 -117 907 -83
rect 941 -117 953 -83
rect 895 -151 953 -117
rect 895 -185 907 -151
rect 941 -185 953 -151
rect 895 -219 953 -185
rect 895 -253 907 -219
rect 941 -253 953 -219
rect 895 -287 953 -253
rect 895 -321 907 -287
rect 941 -321 953 -287
rect 895 -355 953 -321
rect 895 -389 907 -355
rect 941 -389 953 -355
rect 895 -423 953 -389
rect 895 -457 907 -423
rect 941 -457 953 -423
rect 895 -491 953 -457
rect 895 -525 907 -491
rect 941 -525 953 -491
rect 895 -559 953 -525
rect 895 -593 907 -559
rect 941 -593 953 -559
rect 895 -627 953 -593
rect 895 -661 907 -627
rect 941 -661 953 -627
rect 895 -695 953 -661
rect 895 -729 907 -695
rect 941 -729 953 -695
rect 895 -763 953 -729
rect 895 -797 907 -763
rect 941 -797 953 -763
rect 895 -831 953 -797
rect 895 -865 907 -831
rect 941 -865 953 -831
rect 895 -904 953 -865
rect 1203 937 1261 976
rect 1203 903 1215 937
rect 1249 903 1261 937
rect 1203 869 1261 903
rect 1203 835 1215 869
rect 1249 835 1261 869
rect 1203 801 1261 835
rect 1203 767 1215 801
rect 1249 767 1261 801
rect 1203 733 1261 767
rect 1203 699 1215 733
rect 1249 699 1261 733
rect 1203 665 1261 699
rect 1203 631 1215 665
rect 1249 631 1261 665
rect 1203 597 1261 631
rect 1203 563 1215 597
rect 1249 563 1261 597
rect 1203 529 1261 563
rect 1203 495 1215 529
rect 1249 495 1261 529
rect 1203 461 1261 495
rect 1203 427 1215 461
rect 1249 427 1261 461
rect 1203 393 1261 427
rect 1203 359 1215 393
rect 1249 359 1261 393
rect 1203 325 1261 359
rect 1203 291 1215 325
rect 1249 291 1261 325
rect 1203 257 1261 291
rect 1203 223 1215 257
rect 1249 223 1261 257
rect 1203 189 1261 223
rect 1203 155 1215 189
rect 1249 155 1261 189
rect 1203 121 1261 155
rect 1203 87 1215 121
rect 1249 87 1261 121
rect 1203 53 1261 87
rect 1203 19 1215 53
rect 1249 19 1261 53
rect 1203 -15 1261 19
rect 1203 -49 1215 -15
rect 1249 -49 1261 -15
rect 1203 -83 1261 -49
rect 1203 -117 1215 -83
rect 1249 -117 1261 -83
rect 1203 -151 1261 -117
rect 1203 -185 1215 -151
rect 1249 -185 1261 -151
rect 1203 -219 1261 -185
rect 1203 -253 1215 -219
rect 1249 -253 1261 -219
rect 1203 -287 1261 -253
rect 1203 -321 1215 -287
rect 1249 -321 1261 -287
rect 1203 -355 1261 -321
rect 1203 -389 1215 -355
rect 1249 -389 1261 -355
rect 1203 -423 1261 -389
rect 1203 -457 1215 -423
rect 1249 -457 1261 -423
rect 1203 -491 1261 -457
rect 1203 -525 1215 -491
rect 1249 -525 1261 -491
rect 1203 -559 1261 -525
rect 1203 -593 1215 -559
rect 1249 -593 1261 -559
rect 1203 -627 1261 -593
rect 1203 -661 1215 -627
rect 1249 -661 1261 -627
rect 1203 -695 1261 -661
rect 1203 -729 1215 -695
rect 1249 -729 1261 -695
rect 1203 -763 1261 -729
rect 1203 -797 1215 -763
rect 1249 -797 1261 -763
rect 1203 -831 1261 -797
rect 1203 -865 1215 -831
rect 1249 -865 1261 -831
rect 1203 -904 1261 -865
rect 1511 937 1569 976
rect 1511 903 1523 937
rect 1557 903 1569 937
rect 1511 869 1569 903
rect 1511 835 1523 869
rect 1557 835 1569 869
rect 1511 801 1569 835
rect 1511 767 1523 801
rect 1557 767 1569 801
rect 1511 733 1569 767
rect 1511 699 1523 733
rect 1557 699 1569 733
rect 1511 665 1569 699
rect 1511 631 1523 665
rect 1557 631 1569 665
rect 1511 597 1569 631
rect 1511 563 1523 597
rect 1557 563 1569 597
rect 1511 529 1569 563
rect 1511 495 1523 529
rect 1557 495 1569 529
rect 1511 461 1569 495
rect 1511 427 1523 461
rect 1557 427 1569 461
rect 1511 393 1569 427
rect 1511 359 1523 393
rect 1557 359 1569 393
rect 1511 325 1569 359
rect 1511 291 1523 325
rect 1557 291 1569 325
rect 1511 257 1569 291
rect 1511 223 1523 257
rect 1557 223 1569 257
rect 1511 189 1569 223
rect 1511 155 1523 189
rect 1557 155 1569 189
rect 1511 121 1569 155
rect 1511 87 1523 121
rect 1557 87 1569 121
rect 1511 53 1569 87
rect 1511 19 1523 53
rect 1557 19 1569 53
rect 1511 -15 1569 19
rect 1511 -49 1523 -15
rect 1557 -49 1569 -15
rect 1511 -83 1569 -49
rect 1511 -117 1523 -83
rect 1557 -117 1569 -83
rect 1511 -151 1569 -117
rect 1511 -185 1523 -151
rect 1557 -185 1569 -151
rect 1511 -219 1569 -185
rect 1511 -253 1523 -219
rect 1557 -253 1569 -219
rect 1511 -287 1569 -253
rect 1511 -321 1523 -287
rect 1557 -321 1569 -287
rect 1511 -355 1569 -321
rect 1511 -389 1523 -355
rect 1557 -389 1569 -355
rect 1511 -423 1569 -389
rect 1511 -457 1523 -423
rect 1557 -457 1569 -423
rect 1511 -491 1569 -457
rect 1511 -525 1523 -491
rect 1557 -525 1569 -491
rect 1511 -559 1569 -525
rect 1511 -593 1523 -559
rect 1557 -593 1569 -559
rect 1511 -627 1569 -593
rect 1511 -661 1523 -627
rect 1557 -661 1569 -627
rect 1511 -695 1569 -661
rect 1511 -729 1523 -695
rect 1557 -729 1569 -695
rect 1511 -763 1569 -729
rect 1511 -797 1523 -763
rect 1557 -797 1569 -763
rect 1511 -831 1569 -797
rect 1511 -865 1523 -831
rect 1557 -865 1569 -831
rect 1511 -904 1569 -865
rect 1819 937 1877 976
rect 1819 903 1831 937
rect 1865 903 1877 937
rect 1819 869 1877 903
rect 1819 835 1831 869
rect 1865 835 1877 869
rect 1819 801 1877 835
rect 1819 767 1831 801
rect 1865 767 1877 801
rect 1819 733 1877 767
rect 1819 699 1831 733
rect 1865 699 1877 733
rect 1819 665 1877 699
rect 1819 631 1831 665
rect 1865 631 1877 665
rect 1819 597 1877 631
rect 1819 563 1831 597
rect 1865 563 1877 597
rect 1819 529 1877 563
rect 1819 495 1831 529
rect 1865 495 1877 529
rect 1819 461 1877 495
rect 1819 427 1831 461
rect 1865 427 1877 461
rect 1819 393 1877 427
rect 1819 359 1831 393
rect 1865 359 1877 393
rect 1819 325 1877 359
rect 1819 291 1831 325
rect 1865 291 1877 325
rect 1819 257 1877 291
rect 1819 223 1831 257
rect 1865 223 1877 257
rect 1819 189 1877 223
rect 1819 155 1831 189
rect 1865 155 1877 189
rect 1819 121 1877 155
rect 1819 87 1831 121
rect 1865 87 1877 121
rect 1819 53 1877 87
rect 1819 19 1831 53
rect 1865 19 1877 53
rect 1819 -15 1877 19
rect 1819 -49 1831 -15
rect 1865 -49 1877 -15
rect 1819 -83 1877 -49
rect 1819 -117 1831 -83
rect 1865 -117 1877 -83
rect 1819 -151 1877 -117
rect 1819 -185 1831 -151
rect 1865 -185 1877 -151
rect 1819 -219 1877 -185
rect 1819 -253 1831 -219
rect 1865 -253 1877 -219
rect 1819 -287 1877 -253
rect 1819 -321 1831 -287
rect 1865 -321 1877 -287
rect 1819 -355 1877 -321
rect 1819 -389 1831 -355
rect 1865 -389 1877 -355
rect 1819 -423 1877 -389
rect 1819 -457 1831 -423
rect 1865 -457 1877 -423
rect 1819 -491 1877 -457
rect 1819 -525 1831 -491
rect 1865 -525 1877 -491
rect 1819 -559 1877 -525
rect 1819 -593 1831 -559
rect 1865 -593 1877 -559
rect 1819 -627 1877 -593
rect 1819 -661 1831 -627
rect 1865 -661 1877 -627
rect 1819 -695 1877 -661
rect 1819 -729 1831 -695
rect 1865 -729 1877 -695
rect 1819 -763 1877 -729
rect 1819 -797 1831 -763
rect 1865 -797 1877 -763
rect 1819 -831 1877 -797
rect 1819 -865 1831 -831
rect 1865 -865 1877 -831
rect 1819 -904 1877 -865
rect 2127 937 2185 976
rect 2127 903 2139 937
rect 2173 903 2185 937
rect 2127 869 2185 903
rect 2127 835 2139 869
rect 2173 835 2185 869
rect 2127 801 2185 835
rect 2127 767 2139 801
rect 2173 767 2185 801
rect 2127 733 2185 767
rect 2127 699 2139 733
rect 2173 699 2185 733
rect 2127 665 2185 699
rect 2127 631 2139 665
rect 2173 631 2185 665
rect 2127 597 2185 631
rect 2127 563 2139 597
rect 2173 563 2185 597
rect 2127 529 2185 563
rect 2127 495 2139 529
rect 2173 495 2185 529
rect 2127 461 2185 495
rect 2127 427 2139 461
rect 2173 427 2185 461
rect 2127 393 2185 427
rect 2127 359 2139 393
rect 2173 359 2185 393
rect 2127 325 2185 359
rect 2127 291 2139 325
rect 2173 291 2185 325
rect 2127 257 2185 291
rect 2127 223 2139 257
rect 2173 223 2185 257
rect 2127 189 2185 223
rect 2127 155 2139 189
rect 2173 155 2185 189
rect 2127 121 2185 155
rect 2127 87 2139 121
rect 2173 87 2185 121
rect 2127 53 2185 87
rect 2127 19 2139 53
rect 2173 19 2185 53
rect 2127 -15 2185 19
rect 2127 -49 2139 -15
rect 2173 -49 2185 -15
rect 2127 -83 2185 -49
rect 2127 -117 2139 -83
rect 2173 -117 2185 -83
rect 2127 -151 2185 -117
rect 2127 -185 2139 -151
rect 2173 -185 2185 -151
rect 2127 -219 2185 -185
rect 2127 -253 2139 -219
rect 2173 -253 2185 -219
rect 2127 -287 2185 -253
rect 2127 -321 2139 -287
rect 2173 -321 2185 -287
rect 2127 -355 2185 -321
rect 2127 -389 2139 -355
rect 2173 -389 2185 -355
rect 2127 -423 2185 -389
rect 2127 -457 2139 -423
rect 2173 -457 2185 -423
rect 2127 -491 2185 -457
rect 2127 -525 2139 -491
rect 2173 -525 2185 -491
rect 2127 -559 2185 -525
rect 2127 -593 2139 -559
rect 2173 -593 2185 -559
rect 2127 -627 2185 -593
rect 2127 -661 2139 -627
rect 2173 -661 2185 -627
rect 2127 -695 2185 -661
rect 2127 -729 2139 -695
rect 2173 -729 2185 -695
rect 2127 -763 2185 -729
rect 2127 -797 2139 -763
rect 2173 -797 2185 -763
rect 2127 -831 2185 -797
rect 2127 -865 2139 -831
rect 2173 -865 2185 -831
rect 2127 -904 2185 -865
rect 2435 937 2493 976
rect 2435 903 2447 937
rect 2481 903 2493 937
rect 2435 869 2493 903
rect 2435 835 2447 869
rect 2481 835 2493 869
rect 2435 801 2493 835
rect 2435 767 2447 801
rect 2481 767 2493 801
rect 2435 733 2493 767
rect 2435 699 2447 733
rect 2481 699 2493 733
rect 2435 665 2493 699
rect 2435 631 2447 665
rect 2481 631 2493 665
rect 2435 597 2493 631
rect 2435 563 2447 597
rect 2481 563 2493 597
rect 2435 529 2493 563
rect 2435 495 2447 529
rect 2481 495 2493 529
rect 2435 461 2493 495
rect 2435 427 2447 461
rect 2481 427 2493 461
rect 2435 393 2493 427
rect 2435 359 2447 393
rect 2481 359 2493 393
rect 2435 325 2493 359
rect 2435 291 2447 325
rect 2481 291 2493 325
rect 2435 257 2493 291
rect 2435 223 2447 257
rect 2481 223 2493 257
rect 2435 189 2493 223
rect 2435 155 2447 189
rect 2481 155 2493 189
rect 2435 121 2493 155
rect 2435 87 2447 121
rect 2481 87 2493 121
rect 2435 53 2493 87
rect 2435 19 2447 53
rect 2481 19 2493 53
rect 2435 -15 2493 19
rect 2435 -49 2447 -15
rect 2481 -49 2493 -15
rect 2435 -83 2493 -49
rect 2435 -117 2447 -83
rect 2481 -117 2493 -83
rect 2435 -151 2493 -117
rect 2435 -185 2447 -151
rect 2481 -185 2493 -151
rect 2435 -219 2493 -185
rect 2435 -253 2447 -219
rect 2481 -253 2493 -219
rect 2435 -287 2493 -253
rect 2435 -321 2447 -287
rect 2481 -321 2493 -287
rect 2435 -355 2493 -321
rect 2435 -389 2447 -355
rect 2481 -389 2493 -355
rect 2435 -423 2493 -389
rect 2435 -457 2447 -423
rect 2481 -457 2493 -423
rect 2435 -491 2493 -457
rect 2435 -525 2447 -491
rect 2481 -525 2493 -491
rect 2435 -559 2493 -525
rect 2435 -593 2447 -559
rect 2481 -593 2493 -559
rect 2435 -627 2493 -593
rect 2435 -661 2447 -627
rect 2481 -661 2493 -627
rect 2435 -695 2493 -661
rect 2435 -729 2447 -695
rect 2481 -729 2493 -695
rect 2435 -763 2493 -729
rect 2435 -797 2447 -763
rect 2481 -797 2493 -763
rect 2435 -831 2493 -797
rect 2435 -865 2447 -831
rect 2481 -865 2493 -831
rect 2435 -904 2493 -865
rect 2743 937 2801 976
rect 2743 903 2755 937
rect 2789 903 2801 937
rect 2743 869 2801 903
rect 2743 835 2755 869
rect 2789 835 2801 869
rect 2743 801 2801 835
rect 2743 767 2755 801
rect 2789 767 2801 801
rect 2743 733 2801 767
rect 2743 699 2755 733
rect 2789 699 2801 733
rect 2743 665 2801 699
rect 2743 631 2755 665
rect 2789 631 2801 665
rect 2743 597 2801 631
rect 2743 563 2755 597
rect 2789 563 2801 597
rect 2743 529 2801 563
rect 2743 495 2755 529
rect 2789 495 2801 529
rect 2743 461 2801 495
rect 2743 427 2755 461
rect 2789 427 2801 461
rect 2743 393 2801 427
rect 2743 359 2755 393
rect 2789 359 2801 393
rect 2743 325 2801 359
rect 2743 291 2755 325
rect 2789 291 2801 325
rect 2743 257 2801 291
rect 2743 223 2755 257
rect 2789 223 2801 257
rect 2743 189 2801 223
rect 2743 155 2755 189
rect 2789 155 2801 189
rect 2743 121 2801 155
rect 2743 87 2755 121
rect 2789 87 2801 121
rect 2743 53 2801 87
rect 2743 19 2755 53
rect 2789 19 2801 53
rect 2743 -15 2801 19
rect 2743 -49 2755 -15
rect 2789 -49 2801 -15
rect 2743 -83 2801 -49
rect 2743 -117 2755 -83
rect 2789 -117 2801 -83
rect 2743 -151 2801 -117
rect 2743 -185 2755 -151
rect 2789 -185 2801 -151
rect 2743 -219 2801 -185
rect 2743 -253 2755 -219
rect 2789 -253 2801 -219
rect 2743 -287 2801 -253
rect 2743 -321 2755 -287
rect 2789 -321 2801 -287
rect 2743 -355 2801 -321
rect 2743 -389 2755 -355
rect 2789 -389 2801 -355
rect 2743 -423 2801 -389
rect 2743 -457 2755 -423
rect 2789 -457 2801 -423
rect 2743 -491 2801 -457
rect 2743 -525 2755 -491
rect 2789 -525 2801 -491
rect 2743 -559 2801 -525
rect 2743 -593 2755 -559
rect 2789 -593 2801 -559
rect 2743 -627 2801 -593
rect 2743 -661 2755 -627
rect 2789 -661 2801 -627
rect 2743 -695 2801 -661
rect 2743 -729 2755 -695
rect 2789 -729 2801 -695
rect 2743 -763 2801 -729
rect 2743 -797 2755 -763
rect 2789 -797 2801 -763
rect 2743 -831 2801 -797
rect 2743 -865 2755 -831
rect 2789 -865 2801 -831
rect 2743 -904 2801 -865
<< mvpdiffc >>
rect -2789 903 -2755 937
rect -2789 835 -2755 869
rect -2789 767 -2755 801
rect -2789 699 -2755 733
rect -2789 631 -2755 665
rect -2789 563 -2755 597
rect -2789 495 -2755 529
rect -2789 427 -2755 461
rect -2789 359 -2755 393
rect -2789 291 -2755 325
rect -2789 223 -2755 257
rect -2789 155 -2755 189
rect -2789 87 -2755 121
rect -2789 19 -2755 53
rect -2789 -49 -2755 -15
rect -2789 -117 -2755 -83
rect -2789 -185 -2755 -151
rect -2789 -253 -2755 -219
rect -2789 -321 -2755 -287
rect -2789 -389 -2755 -355
rect -2789 -457 -2755 -423
rect -2789 -525 -2755 -491
rect -2789 -593 -2755 -559
rect -2789 -661 -2755 -627
rect -2789 -729 -2755 -695
rect -2789 -797 -2755 -763
rect -2789 -865 -2755 -831
rect -2481 903 -2447 937
rect -2481 835 -2447 869
rect -2481 767 -2447 801
rect -2481 699 -2447 733
rect -2481 631 -2447 665
rect -2481 563 -2447 597
rect -2481 495 -2447 529
rect -2481 427 -2447 461
rect -2481 359 -2447 393
rect -2481 291 -2447 325
rect -2481 223 -2447 257
rect -2481 155 -2447 189
rect -2481 87 -2447 121
rect -2481 19 -2447 53
rect -2481 -49 -2447 -15
rect -2481 -117 -2447 -83
rect -2481 -185 -2447 -151
rect -2481 -253 -2447 -219
rect -2481 -321 -2447 -287
rect -2481 -389 -2447 -355
rect -2481 -457 -2447 -423
rect -2481 -525 -2447 -491
rect -2481 -593 -2447 -559
rect -2481 -661 -2447 -627
rect -2481 -729 -2447 -695
rect -2481 -797 -2447 -763
rect -2481 -865 -2447 -831
rect -2173 903 -2139 937
rect -2173 835 -2139 869
rect -2173 767 -2139 801
rect -2173 699 -2139 733
rect -2173 631 -2139 665
rect -2173 563 -2139 597
rect -2173 495 -2139 529
rect -2173 427 -2139 461
rect -2173 359 -2139 393
rect -2173 291 -2139 325
rect -2173 223 -2139 257
rect -2173 155 -2139 189
rect -2173 87 -2139 121
rect -2173 19 -2139 53
rect -2173 -49 -2139 -15
rect -2173 -117 -2139 -83
rect -2173 -185 -2139 -151
rect -2173 -253 -2139 -219
rect -2173 -321 -2139 -287
rect -2173 -389 -2139 -355
rect -2173 -457 -2139 -423
rect -2173 -525 -2139 -491
rect -2173 -593 -2139 -559
rect -2173 -661 -2139 -627
rect -2173 -729 -2139 -695
rect -2173 -797 -2139 -763
rect -2173 -865 -2139 -831
rect -1865 903 -1831 937
rect -1865 835 -1831 869
rect -1865 767 -1831 801
rect -1865 699 -1831 733
rect -1865 631 -1831 665
rect -1865 563 -1831 597
rect -1865 495 -1831 529
rect -1865 427 -1831 461
rect -1865 359 -1831 393
rect -1865 291 -1831 325
rect -1865 223 -1831 257
rect -1865 155 -1831 189
rect -1865 87 -1831 121
rect -1865 19 -1831 53
rect -1865 -49 -1831 -15
rect -1865 -117 -1831 -83
rect -1865 -185 -1831 -151
rect -1865 -253 -1831 -219
rect -1865 -321 -1831 -287
rect -1865 -389 -1831 -355
rect -1865 -457 -1831 -423
rect -1865 -525 -1831 -491
rect -1865 -593 -1831 -559
rect -1865 -661 -1831 -627
rect -1865 -729 -1831 -695
rect -1865 -797 -1831 -763
rect -1865 -865 -1831 -831
rect -1557 903 -1523 937
rect -1557 835 -1523 869
rect -1557 767 -1523 801
rect -1557 699 -1523 733
rect -1557 631 -1523 665
rect -1557 563 -1523 597
rect -1557 495 -1523 529
rect -1557 427 -1523 461
rect -1557 359 -1523 393
rect -1557 291 -1523 325
rect -1557 223 -1523 257
rect -1557 155 -1523 189
rect -1557 87 -1523 121
rect -1557 19 -1523 53
rect -1557 -49 -1523 -15
rect -1557 -117 -1523 -83
rect -1557 -185 -1523 -151
rect -1557 -253 -1523 -219
rect -1557 -321 -1523 -287
rect -1557 -389 -1523 -355
rect -1557 -457 -1523 -423
rect -1557 -525 -1523 -491
rect -1557 -593 -1523 -559
rect -1557 -661 -1523 -627
rect -1557 -729 -1523 -695
rect -1557 -797 -1523 -763
rect -1557 -865 -1523 -831
rect -1249 903 -1215 937
rect -1249 835 -1215 869
rect -1249 767 -1215 801
rect -1249 699 -1215 733
rect -1249 631 -1215 665
rect -1249 563 -1215 597
rect -1249 495 -1215 529
rect -1249 427 -1215 461
rect -1249 359 -1215 393
rect -1249 291 -1215 325
rect -1249 223 -1215 257
rect -1249 155 -1215 189
rect -1249 87 -1215 121
rect -1249 19 -1215 53
rect -1249 -49 -1215 -15
rect -1249 -117 -1215 -83
rect -1249 -185 -1215 -151
rect -1249 -253 -1215 -219
rect -1249 -321 -1215 -287
rect -1249 -389 -1215 -355
rect -1249 -457 -1215 -423
rect -1249 -525 -1215 -491
rect -1249 -593 -1215 -559
rect -1249 -661 -1215 -627
rect -1249 -729 -1215 -695
rect -1249 -797 -1215 -763
rect -1249 -865 -1215 -831
rect -941 903 -907 937
rect -941 835 -907 869
rect -941 767 -907 801
rect -941 699 -907 733
rect -941 631 -907 665
rect -941 563 -907 597
rect -941 495 -907 529
rect -941 427 -907 461
rect -941 359 -907 393
rect -941 291 -907 325
rect -941 223 -907 257
rect -941 155 -907 189
rect -941 87 -907 121
rect -941 19 -907 53
rect -941 -49 -907 -15
rect -941 -117 -907 -83
rect -941 -185 -907 -151
rect -941 -253 -907 -219
rect -941 -321 -907 -287
rect -941 -389 -907 -355
rect -941 -457 -907 -423
rect -941 -525 -907 -491
rect -941 -593 -907 -559
rect -941 -661 -907 -627
rect -941 -729 -907 -695
rect -941 -797 -907 -763
rect -941 -865 -907 -831
rect -633 903 -599 937
rect -633 835 -599 869
rect -633 767 -599 801
rect -633 699 -599 733
rect -633 631 -599 665
rect -633 563 -599 597
rect -633 495 -599 529
rect -633 427 -599 461
rect -633 359 -599 393
rect -633 291 -599 325
rect -633 223 -599 257
rect -633 155 -599 189
rect -633 87 -599 121
rect -633 19 -599 53
rect -633 -49 -599 -15
rect -633 -117 -599 -83
rect -633 -185 -599 -151
rect -633 -253 -599 -219
rect -633 -321 -599 -287
rect -633 -389 -599 -355
rect -633 -457 -599 -423
rect -633 -525 -599 -491
rect -633 -593 -599 -559
rect -633 -661 -599 -627
rect -633 -729 -599 -695
rect -633 -797 -599 -763
rect -633 -865 -599 -831
rect -325 903 -291 937
rect -325 835 -291 869
rect -325 767 -291 801
rect -325 699 -291 733
rect -325 631 -291 665
rect -325 563 -291 597
rect -325 495 -291 529
rect -325 427 -291 461
rect -325 359 -291 393
rect -325 291 -291 325
rect -325 223 -291 257
rect -325 155 -291 189
rect -325 87 -291 121
rect -325 19 -291 53
rect -325 -49 -291 -15
rect -325 -117 -291 -83
rect -325 -185 -291 -151
rect -325 -253 -291 -219
rect -325 -321 -291 -287
rect -325 -389 -291 -355
rect -325 -457 -291 -423
rect -325 -525 -291 -491
rect -325 -593 -291 -559
rect -325 -661 -291 -627
rect -325 -729 -291 -695
rect -325 -797 -291 -763
rect -325 -865 -291 -831
rect -17 903 17 937
rect -17 835 17 869
rect -17 767 17 801
rect -17 699 17 733
rect -17 631 17 665
rect -17 563 17 597
rect -17 495 17 529
rect -17 427 17 461
rect -17 359 17 393
rect -17 291 17 325
rect -17 223 17 257
rect -17 155 17 189
rect -17 87 17 121
rect -17 19 17 53
rect -17 -49 17 -15
rect -17 -117 17 -83
rect -17 -185 17 -151
rect -17 -253 17 -219
rect -17 -321 17 -287
rect -17 -389 17 -355
rect -17 -457 17 -423
rect -17 -525 17 -491
rect -17 -593 17 -559
rect -17 -661 17 -627
rect -17 -729 17 -695
rect -17 -797 17 -763
rect -17 -865 17 -831
rect 291 903 325 937
rect 291 835 325 869
rect 291 767 325 801
rect 291 699 325 733
rect 291 631 325 665
rect 291 563 325 597
rect 291 495 325 529
rect 291 427 325 461
rect 291 359 325 393
rect 291 291 325 325
rect 291 223 325 257
rect 291 155 325 189
rect 291 87 325 121
rect 291 19 325 53
rect 291 -49 325 -15
rect 291 -117 325 -83
rect 291 -185 325 -151
rect 291 -253 325 -219
rect 291 -321 325 -287
rect 291 -389 325 -355
rect 291 -457 325 -423
rect 291 -525 325 -491
rect 291 -593 325 -559
rect 291 -661 325 -627
rect 291 -729 325 -695
rect 291 -797 325 -763
rect 291 -865 325 -831
rect 599 903 633 937
rect 599 835 633 869
rect 599 767 633 801
rect 599 699 633 733
rect 599 631 633 665
rect 599 563 633 597
rect 599 495 633 529
rect 599 427 633 461
rect 599 359 633 393
rect 599 291 633 325
rect 599 223 633 257
rect 599 155 633 189
rect 599 87 633 121
rect 599 19 633 53
rect 599 -49 633 -15
rect 599 -117 633 -83
rect 599 -185 633 -151
rect 599 -253 633 -219
rect 599 -321 633 -287
rect 599 -389 633 -355
rect 599 -457 633 -423
rect 599 -525 633 -491
rect 599 -593 633 -559
rect 599 -661 633 -627
rect 599 -729 633 -695
rect 599 -797 633 -763
rect 599 -865 633 -831
rect 907 903 941 937
rect 907 835 941 869
rect 907 767 941 801
rect 907 699 941 733
rect 907 631 941 665
rect 907 563 941 597
rect 907 495 941 529
rect 907 427 941 461
rect 907 359 941 393
rect 907 291 941 325
rect 907 223 941 257
rect 907 155 941 189
rect 907 87 941 121
rect 907 19 941 53
rect 907 -49 941 -15
rect 907 -117 941 -83
rect 907 -185 941 -151
rect 907 -253 941 -219
rect 907 -321 941 -287
rect 907 -389 941 -355
rect 907 -457 941 -423
rect 907 -525 941 -491
rect 907 -593 941 -559
rect 907 -661 941 -627
rect 907 -729 941 -695
rect 907 -797 941 -763
rect 907 -865 941 -831
rect 1215 903 1249 937
rect 1215 835 1249 869
rect 1215 767 1249 801
rect 1215 699 1249 733
rect 1215 631 1249 665
rect 1215 563 1249 597
rect 1215 495 1249 529
rect 1215 427 1249 461
rect 1215 359 1249 393
rect 1215 291 1249 325
rect 1215 223 1249 257
rect 1215 155 1249 189
rect 1215 87 1249 121
rect 1215 19 1249 53
rect 1215 -49 1249 -15
rect 1215 -117 1249 -83
rect 1215 -185 1249 -151
rect 1215 -253 1249 -219
rect 1215 -321 1249 -287
rect 1215 -389 1249 -355
rect 1215 -457 1249 -423
rect 1215 -525 1249 -491
rect 1215 -593 1249 -559
rect 1215 -661 1249 -627
rect 1215 -729 1249 -695
rect 1215 -797 1249 -763
rect 1215 -865 1249 -831
rect 1523 903 1557 937
rect 1523 835 1557 869
rect 1523 767 1557 801
rect 1523 699 1557 733
rect 1523 631 1557 665
rect 1523 563 1557 597
rect 1523 495 1557 529
rect 1523 427 1557 461
rect 1523 359 1557 393
rect 1523 291 1557 325
rect 1523 223 1557 257
rect 1523 155 1557 189
rect 1523 87 1557 121
rect 1523 19 1557 53
rect 1523 -49 1557 -15
rect 1523 -117 1557 -83
rect 1523 -185 1557 -151
rect 1523 -253 1557 -219
rect 1523 -321 1557 -287
rect 1523 -389 1557 -355
rect 1523 -457 1557 -423
rect 1523 -525 1557 -491
rect 1523 -593 1557 -559
rect 1523 -661 1557 -627
rect 1523 -729 1557 -695
rect 1523 -797 1557 -763
rect 1523 -865 1557 -831
rect 1831 903 1865 937
rect 1831 835 1865 869
rect 1831 767 1865 801
rect 1831 699 1865 733
rect 1831 631 1865 665
rect 1831 563 1865 597
rect 1831 495 1865 529
rect 1831 427 1865 461
rect 1831 359 1865 393
rect 1831 291 1865 325
rect 1831 223 1865 257
rect 1831 155 1865 189
rect 1831 87 1865 121
rect 1831 19 1865 53
rect 1831 -49 1865 -15
rect 1831 -117 1865 -83
rect 1831 -185 1865 -151
rect 1831 -253 1865 -219
rect 1831 -321 1865 -287
rect 1831 -389 1865 -355
rect 1831 -457 1865 -423
rect 1831 -525 1865 -491
rect 1831 -593 1865 -559
rect 1831 -661 1865 -627
rect 1831 -729 1865 -695
rect 1831 -797 1865 -763
rect 1831 -865 1865 -831
rect 2139 903 2173 937
rect 2139 835 2173 869
rect 2139 767 2173 801
rect 2139 699 2173 733
rect 2139 631 2173 665
rect 2139 563 2173 597
rect 2139 495 2173 529
rect 2139 427 2173 461
rect 2139 359 2173 393
rect 2139 291 2173 325
rect 2139 223 2173 257
rect 2139 155 2173 189
rect 2139 87 2173 121
rect 2139 19 2173 53
rect 2139 -49 2173 -15
rect 2139 -117 2173 -83
rect 2139 -185 2173 -151
rect 2139 -253 2173 -219
rect 2139 -321 2173 -287
rect 2139 -389 2173 -355
rect 2139 -457 2173 -423
rect 2139 -525 2173 -491
rect 2139 -593 2173 -559
rect 2139 -661 2173 -627
rect 2139 -729 2173 -695
rect 2139 -797 2173 -763
rect 2139 -865 2173 -831
rect 2447 903 2481 937
rect 2447 835 2481 869
rect 2447 767 2481 801
rect 2447 699 2481 733
rect 2447 631 2481 665
rect 2447 563 2481 597
rect 2447 495 2481 529
rect 2447 427 2481 461
rect 2447 359 2481 393
rect 2447 291 2481 325
rect 2447 223 2481 257
rect 2447 155 2481 189
rect 2447 87 2481 121
rect 2447 19 2481 53
rect 2447 -49 2481 -15
rect 2447 -117 2481 -83
rect 2447 -185 2481 -151
rect 2447 -253 2481 -219
rect 2447 -321 2481 -287
rect 2447 -389 2481 -355
rect 2447 -457 2481 -423
rect 2447 -525 2481 -491
rect 2447 -593 2481 -559
rect 2447 -661 2481 -627
rect 2447 -729 2481 -695
rect 2447 -797 2481 -763
rect 2447 -865 2481 -831
rect 2755 903 2789 937
rect 2755 835 2789 869
rect 2755 767 2789 801
rect 2755 699 2789 733
rect 2755 631 2789 665
rect 2755 563 2789 597
rect 2755 495 2789 529
rect 2755 427 2789 461
rect 2755 359 2789 393
rect 2755 291 2789 325
rect 2755 223 2789 257
rect 2755 155 2789 189
rect 2755 87 2789 121
rect 2755 19 2789 53
rect 2755 -49 2789 -15
rect 2755 -117 2789 -83
rect 2755 -185 2789 -151
rect 2755 -253 2789 -219
rect 2755 -321 2789 -287
rect 2755 -389 2789 -355
rect 2755 -457 2789 -423
rect 2755 -525 2789 -491
rect 2755 -593 2789 -559
rect 2755 -661 2789 -627
rect 2755 -729 2789 -695
rect 2755 -797 2789 -763
rect 2755 -865 2789 -831
<< poly >>
rect -2743 976 -2493 1002
rect -2435 976 -2185 1002
rect -2127 976 -1877 1002
rect -1819 976 -1569 1002
rect -1511 976 -1261 1002
rect -1203 976 -953 1002
rect -895 976 -645 1002
rect -587 976 -337 1002
rect -279 976 -29 1002
rect 29 976 279 1002
rect 337 976 587 1002
rect 645 976 895 1002
rect 953 976 1203 1002
rect 1261 976 1511 1002
rect 1569 976 1819 1002
rect 1877 976 2127 1002
rect 2185 976 2435 1002
rect 2493 976 2743 1002
rect -2743 -951 -2493 -904
rect -2743 -968 -2669 -951
rect -2705 -985 -2669 -968
rect -2635 -985 -2601 -951
rect -2567 -968 -2493 -951
rect -2435 -951 -2185 -904
rect -2435 -968 -2361 -951
rect -2567 -985 -2531 -968
rect -2705 -1001 -2531 -985
rect -2397 -985 -2361 -968
rect -2327 -985 -2293 -951
rect -2259 -968 -2185 -951
rect -2127 -951 -1877 -904
rect -2127 -968 -2053 -951
rect -2259 -985 -2223 -968
rect -2397 -1001 -2223 -985
rect -2089 -985 -2053 -968
rect -2019 -985 -1985 -951
rect -1951 -968 -1877 -951
rect -1819 -951 -1569 -904
rect -1819 -968 -1745 -951
rect -1951 -985 -1915 -968
rect -2089 -1001 -1915 -985
rect -1781 -985 -1745 -968
rect -1711 -985 -1677 -951
rect -1643 -968 -1569 -951
rect -1511 -951 -1261 -904
rect -1511 -968 -1437 -951
rect -1643 -985 -1607 -968
rect -1781 -1001 -1607 -985
rect -1473 -985 -1437 -968
rect -1403 -985 -1369 -951
rect -1335 -968 -1261 -951
rect -1203 -951 -953 -904
rect -1203 -968 -1129 -951
rect -1335 -985 -1299 -968
rect -1473 -1001 -1299 -985
rect -1165 -985 -1129 -968
rect -1095 -985 -1061 -951
rect -1027 -968 -953 -951
rect -895 -951 -645 -904
rect -895 -968 -821 -951
rect -1027 -985 -991 -968
rect -1165 -1001 -991 -985
rect -857 -985 -821 -968
rect -787 -985 -753 -951
rect -719 -968 -645 -951
rect -587 -951 -337 -904
rect -587 -968 -513 -951
rect -719 -985 -683 -968
rect -857 -1001 -683 -985
rect -549 -985 -513 -968
rect -479 -985 -445 -951
rect -411 -968 -337 -951
rect -279 -951 -29 -904
rect -279 -968 -205 -951
rect -411 -985 -375 -968
rect -549 -1001 -375 -985
rect -241 -985 -205 -968
rect -171 -985 -137 -951
rect -103 -968 -29 -951
rect 29 -951 279 -904
rect 29 -968 103 -951
rect -103 -985 -67 -968
rect -241 -1001 -67 -985
rect 67 -985 103 -968
rect 137 -985 171 -951
rect 205 -968 279 -951
rect 337 -951 587 -904
rect 337 -968 411 -951
rect 205 -985 241 -968
rect 67 -1001 241 -985
rect 375 -985 411 -968
rect 445 -985 479 -951
rect 513 -968 587 -951
rect 645 -951 895 -904
rect 645 -968 719 -951
rect 513 -985 549 -968
rect 375 -1001 549 -985
rect 683 -985 719 -968
rect 753 -985 787 -951
rect 821 -968 895 -951
rect 953 -951 1203 -904
rect 953 -968 1027 -951
rect 821 -985 857 -968
rect 683 -1001 857 -985
rect 991 -985 1027 -968
rect 1061 -985 1095 -951
rect 1129 -968 1203 -951
rect 1261 -951 1511 -904
rect 1261 -968 1335 -951
rect 1129 -985 1165 -968
rect 991 -1001 1165 -985
rect 1299 -985 1335 -968
rect 1369 -985 1403 -951
rect 1437 -968 1511 -951
rect 1569 -951 1819 -904
rect 1569 -968 1643 -951
rect 1437 -985 1473 -968
rect 1299 -1001 1473 -985
rect 1607 -985 1643 -968
rect 1677 -985 1711 -951
rect 1745 -968 1819 -951
rect 1877 -951 2127 -904
rect 1877 -968 1951 -951
rect 1745 -985 1781 -968
rect 1607 -1001 1781 -985
rect 1915 -985 1951 -968
rect 1985 -985 2019 -951
rect 2053 -968 2127 -951
rect 2185 -951 2435 -904
rect 2185 -968 2259 -951
rect 2053 -985 2089 -968
rect 1915 -1001 2089 -985
rect 2223 -985 2259 -968
rect 2293 -985 2327 -951
rect 2361 -968 2435 -951
rect 2493 -951 2743 -904
rect 2493 -968 2567 -951
rect 2361 -985 2397 -968
rect 2223 -1001 2397 -985
rect 2531 -985 2567 -968
rect 2601 -985 2635 -951
rect 2669 -968 2743 -951
rect 2669 -985 2705 -968
rect 2531 -1001 2705 -985
<< polycont >>
rect -2669 -985 -2635 -951
rect -2601 -985 -2567 -951
rect -2361 -985 -2327 -951
rect -2293 -985 -2259 -951
rect -2053 -985 -2019 -951
rect -1985 -985 -1951 -951
rect -1745 -985 -1711 -951
rect -1677 -985 -1643 -951
rect -1437 -985 -1403 -951
rect -1369 -985 -1335 -951
rect -1129 -985 -1095 -951
rect -1061 -985 -1027 -951
rect -821 -985 -787 -951
rect -753 -985 -719 -951
rect -513 -985 -479 -951
rect -445 -985 -411 -951
rect -205 -985 -171 -951
rect -137 -985 -103 -951
rect 103 -985 137 -951
rect 171 -985 205 -951
rect 411 -985 445 -951
rect 479 -985 513 -951
rect 719 -985 753 -951
rect 787 -985 821 -951
rect 1027 -985 1061 -951
rect 1095 -985 1129 -951
rect 1335 -985 1369 -951
rect 1403 -985 1437 -951
rect 1643 -985 1677 -951
rect 1711 -985 1745 -951
rect 1951 -985 1985 -951
rect 2019 -985 2053 -951
rect 2259 -985 2293 -951
rect 2327 -985 2361 -951
rect 2567 -985 2601 -951
rect 2635 -985 2669 -951
<< locali >>
rect -2789 953 -2755 980
rect -2789 881 -2755 903
rect -2789 809 -2755 835
rect -2789 737 -2755 767
rect -2789 665 -2755 699
rect -2789 597 -2755 631
rect -2789 529 -2755 559
rect -2789 461 -2755 487
rect -2789 393 -2755 415
rect -2789 325 -2755 343
rect -2789 257 -2755 271
rect -2789 189 -2755 199
rect -2789 121 -2755 127
rect -2789 53 -2755 55
rect -2789 17 -2755 19
rect -2789 -55 -2755 -49
rect -2789 -127 -2755 -117
rect -2789 -199 -2755 -185
rect -2789 -271 -2755 -253
rect -2789 -343 -2755 -321
rect -2789 -415 -2755 -389
rect -2789 -487 -2755 -457
rect -2789 -559 -2755 -525
rect -2789 -627 -2755 -593
rect -2789 -695 -2755 -665
rect -2789 -763 -2755 -737
rect -2789 -831 -2755 -809
rect -2789 -908 -2755 -881
rect -2481 953 -2447 980
rect -2481 881 -2447 903
rect -2481 809 -2447 835
rect -2481 737 -2447 767
rect -2481 665 -2447 699
rect -2481 597 -2447 631
rect -2481 529 -2447 559
rect -2481 461 -2447 487
rect -2481 393 -2447 415
rect -2481 325 -2447 343
rect -2481 257 -2447 271
rect -2481 189 -2447 199
rect -2481 121 -2447 127
rect -2481 53 -2447 55
rect -2481 17 -2447 19
rect -2481 -55 -2447 -49
rect -2481 -127 -2447 -117
rect -2481 -199 -2447 -185
rect -2481 -271 -2447 -253
rect -2481 -343 -2447 -321
rect -2481 -415 -2447 -389
rect -2481 -487 -2447 -457
rect -2481 -559 -2447 -525
rect -2481 -627 -2447 -593
rect -2481 -695 -2447 -665
rect -2481 -763 -2447 -737
rect -2481 -831 -2447 -809
rect -2481 -908 -2447 -881
rect -2173 953 -2139 980
rect -2173 881 -2139 903
rect -2173 809 -2139 835
rect -2173 737 -2139 767
rect -2173 665 -2139 699
rect -2173 597 -2139 631
rect -2173 529 -2139 559
rect -2173 461 -2139 487
rect -2173 393 -2139 415
rect -2173 325 -2139 343
rect -2173 257 -2139 271
rect -2173 189 -2139 199
rect -2173 121 -2139 127
rect -2173 53 -2139 55
rect -2173 17 -2139 19
rect -2173 -55 -2139 -49
rect -2173 -127 -2139 -117
rect -2173 -199 -2139 -185
rect -2173 -271 -2139 -253
rect -2173 -343 -2139 -321
rect -2173 -415 -2139 -389
rect -2173 -487 -2139 -457
rect -2173 -559 -2139 -525
rect -2173 -627 -2139 -593
rect -2173 -695 -2139 -665
rect -2173 -763 -2139 -737
rect -2173 -831 -2139 -809
rect -2173 -908 -2139 -881
rect -1865 953 -1831 980
rect -1865 881 -1831 903
rect -1865 809 -1831 835
rect -1865 737 -1831 767
rect -1865 665 -1831 699
rect -1865 597 -1831 631
rect -1865 529 -1831 559
rect -1865 461 -1831 487
rect -1865 393 -1831 415
rect -1865 325 -1831 343
rect -1865 257 -1831 271
rect -1865 189 -1831 199
rect -1865 121 -1831 127
rect -1865 53 -1831 55
rect -1865 17 -1831 19
rect -1865 -55 -1831 -49
rect -1865 -127 -1831 -117
rect -1865 -199 -1831 -185
rect -1865 -271 -1831 -253
rect -1865 -343 -1831 -321
rect -1865 -415 -1831 -389
rect -1865 -487 -1831 -457
rect -1865 -559 -1831 -525
rect -1865 -627 -1831 -593
rect -1865 -695 -1831 -665
rect -1865 -763 -1831 -737
rect -1865 -831 -1831 -809
rect -1865 -908 -1831 -881
rect -1557 953 -1523 980
rect -1557 881 -1523 903
rect -1557 809 -1523 835
rect -1557 737 -1523 767
rect -1557 665 -1523 699
rect -1557 597 -1523 631
rect -1557 529 -1523 559
rect -1557 461 -1523 487
rect -1557 393 -1523 415
rect -1557 325 -1523 343
rect -1557 257 -1523 271
rect -1557 189 -1523 199
rect -1557 121 -1523 127
rect -1557 53 -1523 55
rect -1557 17 -1523 19
rect -1557 -55 -1523 -49
rect -1557 -127 -1523 -117
rect -1557 -199 -1523 -185
rect -1557 -271 -1523 -253
rect -1557 -343 -1523 -321
rect -1557 -415 -1523 -389
rect -1557 -487 -1523 -457
rect -1557 -559 -1523 -525
rect -1557 -627 -1523 -593
rect -1557 -695 -1523 -665
rect -1557 -763 -1523 -737
rect -1557 -831 -1523 -809
rect -1557 -908 -1523 -881
rect -1249 953 -1215 980
rect -1249 881 -1215 903
rect -1249 809 -1215 835
rect -1249 737 -1215 767
rect -1249 665 -1215 699
rect -1249 597 -1215 631
rect -1249 529 -1215 559
rect -1249 461 -1215 487
rect -1249 393 -1215 415
rect -1249 325 -1215 343
rect -1249 257 -1215 271
rect -1249 189 -1215 199
rect -1249 121 -1215 127
rect -1249 53 -1215 55
rect -1249 17 -1215 19
rect -1249 -55 -1215 -49
rect -1249 -127 -1215 -117
rect -1249 -199 -1215 -185
rect -1249 -271 -1215 -253
rect -1249 -343 -1215 -321
rect -1249 -415 -1215 -389
rect -1249 -487 -1215 -457
rect -1249 -559 -1215 -525
rect -1249 -627 -1215 -593
rect -1249 -695 -1215 -665
rect -1249 -763 -1215 -737
rect -1249 -831 -1215 -809
rect -1249 -908 -1215 -881
rect -941 953 -907 980
rect -941 881 -907 903
rect -941 809 -907 835
rect -941 737 -907 767
rect -941 665 -907 699
rect -941 597 -907 631
rect -941 529 -907 559
rect -941 461 -907 487
rect -941 393 -907 415
rect -941 325 -907 343
rect -941 257 -907 271
rect -941 189 -907 199
rect -941 121 -907 127
rect -941 53 -907 55
rect -941 17 -907 19
rect -941 -55 -907 -49
rect -941 -127 -907 -117
rect -941 -199 -907 -185
rect -941 -271 -907 -253
rect -941 -343 -907 -321
rect -941 -415 -907 -389
rect -941 -487 -907 -457
rect -941 -559 -907 -525
rect -941 -627 -907 -593
rect -941 -695 -907 -665
rect -941 -763 -907 -737
rect -941 -831 -907 -809
rect -941 -908 -907 -881
rect -633 953 -599 980
rect -633 881 -599 903
rect -633 809 -599 835
rect -633 737 -599 767
rect -633 665 -599 699
rect -633 597 -599 631
rect -633 529 -599 559
rect -633 461 -599 487
rect -633 393 -599 415
rect -633 325 -599 343
rect -633 257 -599 271
rect -633 189 -599 199
rect -633 121 -599 127
rect -633 53 -599 55
rect -633 17 -599 19
rect -633 -55 -599 -49
rect -633 -127 -599 -117
rect -633 -199 -599 -185
rect -633 -271 -599 -253
rect -633 -343 -599 -321
rect -633 -415 -599 -389
rect -633 -487 -599 -457
rect -633 -559 -599 -525
rect -633 -627 -599 -593
rect -633 -695 -599 -665
rect -633 -763 -599 -737
rect -633 -831 -599 -809
rect -633 -908 -599 -881
rect -325 953 -291 980
rect -325 881 -291 903
rect -325 809 -291 835
rect -325 737 -291 767
rect -325 665 -291 699
rect -325 597 -291 631
rect -325 529 -291 559
rect -325 461 -291 487
rect -325 393 -291 415
rect -325 325 -291 343
rect -325 257 -291 271
rect -325 189 -291 199
rect -325 121 -291 127
rect -325 53 -291 55
rect -325 17 -291 19
rect -325 -55 -291 -49
rect -325 -127 -291 -117
rect -325 -199 -291 -185
rect -325 -271 -291 -253
rect -325 -343 -291 -321
rect -325 -415 -291 -389
rect -325 -487 -291 -457
rect -325 -559 -291 -525
rect -325 -627 -291 -593
rect -325 -695 -291 -665
rect -325 -763 -291 -737
rect -325 -831 -291 -809
rect -325 -908 -291 -881
rect -17 953 17 980
rect -17 881 17 903
rect -17 809 17 835
rect -17 737 17 767
rect -17 665 17 699
rect -17 597 17 631
rect -17 529 17 559
rect -17 461 17 487
rect -17 393 17 415
rect -17 325 17 343
rect -17 257 17 271
rect -17 189 17 199
rect -17 121 17 127
rect -17 53 17 55
rect -17 17 17 19
rect -17 -55 17 -49
rect -17 -127 17 -117
rect -17 -199 17 -185
rect -17 -271 17 -253
rect -17 -343 17 -321
rect -17 -415 17 -389
rect -17 -487 17 -457
rect -17 -559 17 -525
rect -17 -627 17 -593
rect -17 -695 17 -665
rect -17 -763 17 -737
rect -17 -831 17 -809
rect -17 -908 17 -881
rect 291 953 325 980
rect 291 881 325 903
rect 291 809 325 835
rect 291 737 325 767
rect 291 665 325 699
rect 291 597 325 631
rect 291 529 325 559
rect 291 461 325 487
rect 291 393 325 415
rect 291 325 325 343
rect 291 257 325 271
rect 291 189 325 199
rect 291 121 325 127
rect 291 53 325 55
rect 291 17 325 19
rect 291 -55 325 -49
rect 291 -127 325 -117
rect 291 -199 325 -185
rect 291 -271 325 -253
rect 291 -343 325 -321
rect 291 -415 325 -389
rect 291 -487 325 -457
rect 291 -559 325 -525
rect 291 -627 325 -593
rect 291 -695 325 -665
rect 291 -763 325 -737
rect 291 -831 325 -809
rect 291 -908 325 -881
rect 599 953 633 980
rect 599 881 633 903
rect 599 809 633 835
rect 599 737 633 767
rect 599 665 633 699
rect 599 597 633 631
rect 599 529 633 559
rect 599 461 633 487
rect 599 393 633 415
rect 599 325 633 343
rect 599 257 633 271
rect 599 189 633 199
rect 599 121 633 127
rect 599 53 633 55
rect 599 17 633 19
rect 599 -55 633 -49
rect 599 -127 633 -117
rect 599 -199 633 -185
rect 599 -271 633 -253
rect 599 -343 633 -321
rect 599 -415 633 -389
rect 599 -487 633 -457
rect 599 -559 633 -525
rect 599 -627 633 -593
rect 599 -695 633 -665
rect 599 -763 633 -737
rect 599 -831 633 -809
rect 599 -908 633 -881
rect 907 953 941 980
rect 907 881 941 903
rect 907 809 941 835
rect 907 737 941 767
rect 907 665 941 699
rect 907 597 941 631
rect 907 529 941 559
rect 907 461 941 487
rect 907 393 941 415
rect 907 325 941 343
rect 907 257 941 271
rect 907 189 941 199
rect 907 121 941 127
rect 907 53 941 55
rect 907 17 941 19
rect 907 -55 941 -49
rect 907 -127 941 -117
rect 907 -199 941 -185
rect 907 -271 941 -253
rect 907 -343 941 -321
rect 907 -415 941 -389
rect 907 -487 941 -457
rect 907 -559 941 -525
rect 907 -627 941 -593
rect 907 -695 941 -665
rect 907 -763 941 -737
rect 907 -831 941 -809
rect 907 -908 941 -881
rect 1215 953 1249 980
rect 1215 881 1249 903
rect 1215 809 1249 835
rect 1215 737 1249 767
rect 1215 665 1249 699
rect 1215 597 1249 631
rect 1215 529 1249 559
rect 1215 461 1249 487
rect 1215 393 1249 415
rect 1215 325 1249 343
rect 1215 257 1249 271
rect 1215 189 1249 199
rect 1215 121 1249 127
rect 1215 53 1249 55
rect 1215 17 1249 19
rect 1215 -55 1249 -49
rect 1215 -127 1249 -117
rect 1215 -199 1249 -185
rect 1215 -271 1249 -253
rect 1215 -343 1249 -321
rect 1215 -415 1249 -389
rect 1215 -487 1249 -457
rect 1215 -559 1249 -525
rect 1215 -627 1249 -593
rect 1215 -695 1249 -665
rect 1215 -763 1249 -737
rect 1215 -831 1249 -809
rect 1215 -908 1249 -881
rect 1523 953 1557 980
rect 1523 881 1557 903
rect 1523 809 1557 835
rect 1523 737 1557 767
rect 1523 665 1557 699
rect 1523 597 1557 631
rect 1523 529 1557 559
rect 1523 461 1557 487
rect 1523 393 1557 415
rect 1523 325 1557 343
rect 1523 257 1557 271
rect 1523 189 1557 199
rect 1523 121 1557 127
rect 1523 53 1557 55
rect 1523 17 1557 19
rect 1523 -55 1557 -49
rect 1523 -127 1557 -117
rect 1523 -199 1557 -185
rect 1523 -271 1557 -253
rect 1523 -343 1557 -321
rect 1523 -415 1557 -389
rect 1523 -487 1557 -457
rect 1523 -559 1557 -525
rect 1523 -627 1557 -593
rect 1523 -695 1557 -665
rect 1523 -763 1557 -737
rect 1523 -831 1557 -809
rect 1523 -908 1557 -881
rect 1831 953 1865 980
rect 1831 881 1865 903
rect 1831 809 1865 835
rect 1831 737 1865 767
rect 1831 665 1865 699
rect 1831 597 1865 631
rect 1831 529 1865 559
rect 1831 461 1865 487
rect 1831 393 1865 415
rect 1831 325 1865 343
rect 1831 257 1865 271
rect 1831 189 1865 199
rect 1831 121 1865 127
rect 1831 53 1865 55
rect 1831 17 1865 19
rect 1831 -55 1865 -49
rect 1831 -127 1865 -117
rect 1831 -199 1865 -185
rect 1831 -271 1865 -253
rect 1831 -343 1865 -321
rect 1831 -415 1865 -389
rect 1831 -487 1865 -457
rect 1831 -559 1865 -525
rect 1831 -627 1865 -593
rect 1831 -695 1865 -665
rect 1831 -763 1865 -737
rect 1831 -831 1865 -809
rect 1831 -908 1865 -881
rect 2139 953 2173 980
rect 2139 881 2173 903
rect 2139 809 2173 835
rect 2139 737 2173 767
rect 2139 665 2173 699
rect 2139 597 2173 631
rect 2139 529 2173 559
rect 2139 461 2173 487
rect 2139 393 2173 415
rect 2139 325 2173 343
rect 2139 257 2173 271
rect 2139 189 2173 199
rect 2139 121 2173 127
rect 2139 53 2173 55
rect 2139 17 2173 19
rect 2139 -55 2173 -49
rect 2139 -127 2173 -117
rect 2139 -199 2173 -185
rect 2139 -271 2173 -253
rect 2139 -343 2173 -321
rect 2139 -415 2173 -389
rect 2139 -487 2173 -457
rect 2139 -559 2173 -525
rect 2139 -627 2173 -593
rect 2139 -695 2173 -665
rect 2139 -763 2173 -737
rect 2139 -831 2173 -809
rect 2139 -908 2173 -881
rect 2447 953 2481 980
rect 2447 881 2481 903
rect 2447 809 2481 835
rect 2447 737 2481 767
rect 2447 665 2481 699
rect 2447 597 2481 631
rect 2447 529 2481 559
rect 2447 461 2481 487
rect 2447 393 2481 415
rect 2447 325 2481 343
rect 2447 257 2481 271
rect 2447 189 2481 199
rect 2447 121 2481 127
rect 2447 53 2481 55
rect 2447 17 2481 19
rect 2447 -55 2481 -49
rect 2447 -127 2481 -117
rect 2447 -199 2481 -185
rect 2447 -271 2481 -253
rect 2447 -343 2481 -321
rect 2447 -415 2481 -389
rect 2447 -487 2481 -457
rect 2447 -559 2481 -525
rect 2447 -627 2481 -593
rect 2447 -695 2481 -665
rect 2447 -763 2481 -737
rect 2447 -831 2481 -809
rect 2447 -908 2481 -881
rect 2755 953 2789 980
rect 2755 881 2789 903
rect 2755 809 2789 835
rect 2755 737 2789 767
rect 2755 665 2789 699
rect 2755 597 2789 631
rect 2755 529 2789 559
rect 2755 461 2789 487
rect 2755 393 2789 415
rect 2755 325 2789 343
rect 2755 257 2789 271
rect 2755 189 2789 199
rect 2755 121 2789 127
rect 2755 53 2789 55
rect 2755 17 2789 19
rect 2755 -55 2789 -49
rect 2755 -127 2789 -117
rect 2755 -199 2789 -185
rect 2755 -271 2789 -253
rect 2755 -343 2789 -321
rect 2755 -415 2789 -389
rect 2755 -487 2789 -457
rect 2755 -559 2789 -525
rect 2755 -627 2789 -593
rect 2755 -695 2789 -665
rect 2755 -763 2789 -737
rect 2755 -831 2789 -809
rect 2755 -908 2789 -881
rect -2705 -985 -2671 -951
rect -2635 -985 -2601 -951
rect -2565 -985 -2531 -951
rect -2397 -985 -2363 -951
rect -2327 -985 -2293 -951
rect -2257 -985 -2223 -951
rect -2089 -985 -2055 -951
rect -2019 -985 -1985 -951
rect -1949 -985 -1915 -951
rect -1781 -985 -1747 -951
rect -1711 -985 -1677 -951
rect -1641 -985 -1607 -951
rect -1473 -985 -1439 -951
rect -1403 -985 -1369 -951
rect -1333 -985 -1299 -951
rect -1165 -985 -1131 -951
rect -1095 -985 -1061 -951
rect -1025 -985 -991 -951
rect -857 -985 -823 -951
rect -787 -985 -753 -951
rect -717 -985 -683 -951
rect -549 -985 -515 -951
rect -479 -985 -445 -951
rect -409 -985 -375 -951
rect -241 -985 -207 -951
rect -171 -985 -137 -951
rect -101 -985 -67 -951
rect 67 -985 101 -951
rect 137 -985 171 -951
rect 207 -985 241 -951
rect 375 -985 409 -951
rect 445 -985 479 -951
rect 515 -985 549 -951
rect 683 -985 717 -951
rect 753 -985 787 -951
rect 823 -985 857 -951
rect 991 -985 1025 -951
rect 1061 -985 1095 -951
rect 1131 -985 1165 -951
rect 1299 -985 1333 -951
rect 1369 -985 1403 -951
rect 1439 -985 1473 -951
rect 1607 -985 1641 -951
rect 1677 -985 1711 -951
rect 1747 -985 1781 -951
rect 1915 -985 1949 -951
rect 1985 -985 2019 -951
rect 2055 -985 2089 -951
rect 2223 -985 2257 -951
rect 2293 -985 2327 -951
rect 2363 -985 2397 -951
rect 2531 -985 2565 -951
rect 2601 -985 2635 -951
rect 2671 -985 2705 -951
<< viali >>
rect -2789 937 -2755 953
rect -2789 919 -2755 937
rect -2789 869 -2755 881
rect -2789 847 -2755 869
rect -2789 801 -2755 809
rect -2789 775 -2755 801
rect -2789 733 -2755 737
rect -2789 703 -2755 733
rect -2789 631 -2755 665
rect -2789 563 -2755 593
rect -2789 559 -2755 563
rect -2789 495 -2755 521
rect -2789 487 -2755 495
rect -2789 427 -2755 449
rect -2789 415 -2755 427
rect -2789 359 -2755 377
rect -2789 343 -2755 359
rect -2789 291 -2755 305
rect -2789 271 -2755 291
rect -2789 223 -2755 233
rect -2789 199 -2755 223
rect -2789 155 -2755 161
rect -2789 127 -2755 155
rect -2789 87 -2755 89
rect -2789 55 -2755 87
rect -2789 -15 -2755 17
rect -2789 -17 -2755 -15
rect -2789 -83 -2755 -55
rect -2789 -89 -2755 -83
rect -2789 -151 -2755 -127
rect -2789 -161 -2755 -151
rect -2789 -219 -2755 -199
rect -2789 -233 -2755 -219
rect -2789 -287 -2755 -271
rect -2789 -305 -2755 -287
rect -2789 -355 -2755 -343
rect -2789 -377 -2755 -355
rect -2789 -423 -2755 -415
rect -2789 -449 -2755 -423
rect -2789 -491 -2755 -487
rect -2789 -521 -2755 -491
rect -2789 -593 -2755 -559
rect -2789 -661 -2755 -631
rect -2789 -665 -2755 -661
rect -2789 -729 -2755 -703
rect -2789 -737 -2755 -729
rect -2789 -797 -2755 -775
rect -2789 -809 -2755 -797
rect -2789 -865 -2755 -847
rect -2789 -881 -2755 -865
rect -2481 937 -2447 953
rect -2481 919 -2447 937
rect -2481 869 -2447 881
rect -2481 847 -2447 869
rect -2481 801 -2447 809
rect -2481 775 -2447 801
rect -2481 733 -2447 737
rect -2481 703 -2447 733
rect -2481 631 -2447 665
rect -2481 563 -2447 593
rect -2481 559 -2447 563
rect -2481 495 -2447 521
rect -2481 487 -2447 495
rect -2481 427 -2447 449
rect -2481 415 -2447 427
rect -2481 359 -2447 377
rect -2481 343 -2447 359
rect -2481 291 -2447 305
rect -2481 271 -2447 291
rect -2481 223 -2447 233
rect -2481 199 -2447 223
rect -2481 155 -2447 161
rect -2481 127 -2447 155
rect -2481 87 -2447 89
rect -2481 55 -2447 87
rect -2481 -15 -2447 17
rect -2481 -17 -2447 -15
rect -2481 -83 -2447 -55
rect -2481 -89 -2447 -83
rect -2481 -151 -2447 -127
rect -2481 -161 -2447 -151
rect -2481 -219 -2447 -199
rect -2481 -233 -2447 -219
rect -2481 -287 -2447 -271
rect -2481 -305 -2447 -287
rect -2481 -355 -2447 -343
rect -2481 -377 -2447 -355
rect -2481 -423 -2447 -415
rect -2481 -449 -2447 -423
rect -2481 -491 -2447 -487
rect -2481 -521 -2447 -491
rect -2481 -593 -2447 -559
rect -2481 -661 -2447 -631
rect -2481 -665 -2447 -661
rect -2481 -729 -2447 -703
rect -2481 -737 -2447 -729
rect -2481 -797 -2447 -775
rect -2481 -809 -2447 -797
rect -2481 -865 -2447 -847
rect -2481 -881 -2447 -865
rect -2173 937 -2139 953
rect -2173 919 -2139 937
rect -2173 869 -2139 881
rect -2173 847 -2139 869
rect -2173 801 -2139 809
rect -2173 775 -2139 801
rect -2173 733 -2139 737
rect -2173 703 -2139 733
rect -2173 631 -2139 665
rect -2173 563 -2139 593
rect -2173 559 -2139 563
rect -2173 495 -2139 521
rect -2173 487 -2139 495
rect -2173 427 -2139 449
rect -2173 415 -2139 427
rect -2173 359 -2139 377
rect -2173 343 -2139 359
rect -2173 291 -2139 305
rect -2173 271 -2139 291
rect -2173 223 -2139 233
rect -2173 199 -2139 223
rect -2173 155 -2139 161
rect -2173 127 -2139 155
rect -2173 87 -2139 89
rect -2173 55 -2139 87
rect -2173 -15 -2139 17
rect -2173 -17 -2139 -15
rect -2173 -83 -2139 -55
rect -2173 -89 -2139 -83
rect -2173 -151 -2139 -127
rect -2173 -161 -2139 -151
rect -2173 -219 -2139 -199
rect -2173 -233 -2139 -219
rect -2173 -287 -2139 -271
rect -2173 -305 -2139 -287
rect -2173 -355 -2139 -343
rect -2173 -377 -2139 -355
rect -2173 -423 -2139 -415
rect -2173 -449 -2139 -423
rect -2173 -491 -2139 -487
rect -2173 -521 -2139 -491
rect -2173 -593 -2139 -559
rect -2173 -661 -2139 -631
rect -2173 -665 -2139 -661
rect -2173 -729 -2139 -703
rect -2173 -737 -2139 -729
rect -2173 -797 -2139 -775
rect -2173 -809 -2139 -797
rect -2173 -865 -2139 -847
rect -2173 -881 -2139 -865
rect -1865 937 -1831 953
rect -1865 919 -1831 937
rect -1865 869 -1831 881
rect -1865 847 -1831 869
rect -1865 801 -1831 809
rect -1865 775 -1831 801
rect -1865 733 -1831 737
rect -1865 703 -1831 733
rect -1865 631 -1831 665
rect -1865 563 -1831 593
rect -1865 559 -1831 563
rect -1865 495 -1831 521
rect -1865 487 -1831 495
rect -1865 427 -1831 449
rect -1865 415 -1831 427
rect -1865 359 -1831 377
rect -1865 343 -1831 359
rect -1865 291 -1831 305
rect -1865 271 -1831 291
rect -1865 223 -1831 233
rect -1865 199 -1831 223
rect -1865 155 -1831 161
rect -1865 127 -1831 155
rect -1865 87 -1831 89
rect -1865 55 -1831 87
rect -1865 -15 -1831 17
rect -1865 -17 -1831 -15
rect -1865 -83 -1831 -55
rect -1865 -89 -1831 -83
rect -1865 -151 -1831 -127
rect -1865 -161 -1831 -151
rect -1865 -219 -1831 -199
rect -1865 -233 -1831 -219
rect -1865 -287 -1831 -271
rect -1865 -305 -1831 -287
rect -1865 -355 -1831 -343
rect -1865 -377 -1831 -355
rect -1865 -423 -1831 -415
rect -1865 -449 -1831 -423
rect -1865 -491 -1831 -487
rect -1865 -521 -1831 -491
rect -1865 -593 -1831 -559
rect -1865 -661 -1831 -631
rect -1865 -665 -1831 -661
rect -1865 -729 -1831 -703
rect -1865 -737 -1831 -729
rect -1865 -797 -1831 -775
rect -1865 -809 -1831 -797
rect -1865 -865 -1831 -847
rect -1865 -881 -1831 -865
rect -1557 937 -1523 953
rect -1557 919 -1523 937
rect -1557 869 -1523 881
rect -1557 847 -1523 869
rect -1557 801 -1523 809
rect -1557 775 -1523 801
rect -1557 733 -1523 737
rect -1557 703 -1523 733
rect -1557 631 -1523 665
rect -1557 563 -1523 593
rect -1557 559 -1523 563
rect -1557 495 -1523 521
rect -1557 487 -1523 495
rect -1557 427 -1523 449
rect -1557 415 -1523 427
rect -1557 359 -1523 377
rect -1557 343 -1523 359
rect -1557 291 -1523 305
rect -1557 271 -1523 291
rect -1557 223 -1523 233
rect -1557 199 -1523 223
rect -1557 155 -1523 161
rect -1557 127 -1523 155
rect -1557 87 -1523 89
rect -1557 55 -1523 87
rect -1557 -15 -1523 17
rect -1557 -17 -1523 -15
rect -1557 -83 -1523 -55
rect -1557 -89 -1523 -83
rect -1557 -151 -1523 -127
rect -1557 -161 -1523 -151
rect -1557 -219 -1523 -199
rect -1557 -233 -1523 -219
rect -1557 -287 -1523 -271
rect -1557 -305 -1523 -287
rect -1557 -355 -1523 -343
rect -1557 -377 -1523 -355
rect -1557 -423 -1523 -415
rect -1557 -449 -1523 -423
rect -1557 -491 -1523 -487
rect -1557 -521 -1523 -491
rect -1557 -593 -1523 -559
rect -1557 -661 -1523 -631
rect -1557 -665 -1523 -661
rect -1557 -729 -1523 -703
rect -1557 -737 -1523 -729
rect -1557 -797 -1523 -775
rect -1557 -809 -1523 -797
rect -1557 -865 -1523 -847
rect -1557 -881 -1523 -865
rect -1249 937 -1215 953
rect -1249 919 -1215 937
rect -1249 869 -1215 881
rect -1249 847 -1215 869
rect -1249 801 -1215 809
rect -1249 775 -1215 801
rect -1249 733 -1215 737
rect -1249 703 -1215 733
rect -1249 631 -1215 665
rect -1249 563 -1215 593
rect -1249 559 -1215 563
rect -1249 495 -1215 521
rect -1249 487 -1215 495
rect -1249 427 -1215 449
rect -1249 415 -1215 427
rect -1249 359 -1215 377
rect -1249 343 -1215 359
rect -1249 291 -1215 305
rect -1249 271 -1215 291
rect -1249 223 -1215 233
rect -1249 199 -1215 223
rect -1249 155 -1215 161
rect -1249 127 -1215 155
rect -1249 87 -1215 89
rect -1249 55 -1215 87
rect -1249 -15 -1215 17
rect -1249 -17 -1215 -15
rect -1249 -83 -1215 -55
rect -1249 -89 -1215 -83
rect -1249 -151 -1215 -127
rect -1249 -161 -1215 -151
rect -1249 -219 -1215 -199
rect -1249 -233 -1215 -219
rect -1249 -287 -1215 -271
rect -1249 -305 -1215 -287
rect -1249 -355 -1215 -343
rect -1249 -377 -1215 -355
rect -1249 -423 -1215 -415
rect -1249 -449 -1215 -423
rect -1249 -491 -1215 -487
rect -1249 -521 -1215 -491
rect -1249 -593 -1215 -559
rect -1249 -661 -1215 -631
rect -1249 -665 -1215 -661
rect -1249 -729 -1215 -703
rect -1249 -737 -1215 -729
rect -1249 -797 -1215 -775
rect -1249 -809 -1215 -797
rect -1249 -865 -1215 -847
rect -1249 -881 -1215 -865
rect -941 937 -907 953
rect -941 919 -907 937
rect -941 869 -907 881
rect -941 847 -907 869
rect -941 801 -907 809
rect -941 775 -907 801
rect -941 733 -907 737
rect -941 703 -907 733
rect -941 631 -907 665
rect -941 563 -907 593
rect -941 559 -907 563
rect -941 495 -907 521
rect -941 487 -907 495
rect -941 427 -907 449
rect -941 415 -907 427
rect -941 359 -907 377
rect -941 343 -907 359
rect -941 291 -907 305
rect -941 271 -907 291
rect -941 223 -907 233
rect -941 199 -907 223
rect -941 155 -907 161
rect -941 127 -907 155
rect -941 87 -907 89
rect -941 55 -907 87
rect -941 -15 -907 17
rect -941 -17 -907 -15
rect -941 -83 -907 -55
rect -941 -89 -907 -83
rect -941 -151 -907 -127
rect -941 -161 -907 -151
rect -941 -219 -907 -199
rect -941 -233 -907 -219
rect -941 -287 -907 -271
rect -941 -305 -907 -287
rect -941 -355 -907 -343
rect -941 -377 -907 -355
rect -941 -423 -907 -415
rect -941 -449 -907 -423
rect -941 -491 -907 -487
rect -941 -521 -907 -491
rect -941 -593 -907 -559
rect -941 -661 -907 -631
rect -941 -665 -907 -661
rect -941 -729 -907 -703
rect -941 -737 -907 -729
rect -941 -797 -907 -775
rect -941 -809 -907 -797
rect -941 -865 -907 -847
rect -941 -881 -907 -865
rect -633 937 -599 953
rect -633 919 -599 937
rect -633 869 -599 881
rect -633 847 -599 869
rect -633 801 -599 809
rect -633 775 -599 801
rect -633 733 -599 737
rect -633 703 -599 733
rect -633 631 -599 665
rect -633 563 -599 593
rect -633 559 -599 563
rect -633 495 -599 521
rect -633 487 -599 495
rect -633 427 -599 449
rect -633 415 -599 427
rect -633 359 -599 377
rect -633 343 -599 359
rect -633 291 -599 305
rect -633 271 -599 291
rect -633 223 -599 233
rect -633 199 -599 223
rect -633 155 -599 161
rect -633 127 -599 155
rect -633 87 -599 89
rect -633 55 -599 87
rect -633 -15 -599 17
rect -633 -17 -599 -15
rect -633 -83 -599 -55
rect -633 -89 -599 -83
rect -633 -151 -599 -127
rect -633 -161 -599 -151
rect -633 -219 -599 -199
rect -633 -233 -599 -219
rect -633 -287 -599 -271
rect -633 -305 -599 -287
rect -633 -355 -599 -343
rect -633 -377 -599 -355
rect -633 -423 -599 -415
rect -633 -449 -599 -423
rect -633 -491 -599 -487
rect -633 -521 -599 -491
rect -633 -593 -599 -559
rect -633 -661 -599 -631
rect -633 -665 -599 -661
rect -633 -729 -599 -703
rect -633 -737 -599 -729
rect -633 -797 -599 -775
rect -633 -809 -599 -797
rect -633 -865 -599 -847
rect -633 -881 -599 -865
rect -325 937 -291 953
rect -325 919 -291 937
rect -325 869 -291 881
rect -325 847 -291 869
rect -325 801 -291 809
rect -325 775 -291 801
rect -325 733 -291 737
rect -325 703 -291 733
rect -325 631 -291 665
rect -325 563 -291 593
rect -325 559 -291 563
rect -325 495 -291 521
rect -325 487 -291 495
rect -325 427 -291 449
rect -325 415 -291 427
rect -325 359 -291 377
rect -325 343 -291 359
rect -325 291 -291 305
rect -325 271 -291 291
rect -325 223 -291 233
rect -325 199 -291 223
rect -325 155 -291 161
rect -325 127 -291 155
rect -325 87 -291 89
rect -325 55 -291 87
rect -325 -15 -291 17
rect -325 -17 -291 -15
rect -325 -83 -291 -55
rect -325 -89 -291 -83
rect -325 -151 -291 -127
rect -325 -161 -291 -151
rect -325 -219 -291 -199
rect -325 -233 -291 -219
rect -325 -287 -291 -271
rect -325 -305 -291 -287
rect -325 -355 -291 -343
rect -325 -377 -291 -355
rect -325 -423 -291 -415
rect -325 -449 -291 -423
rect -325 -491 -291 -487
rect -325 -521 -291 -491
rect -325 -593 -291 -559
rect -325 -661 -291 -631
rect -325 -665 -291 -661
rect -325 -729 -291 -703
rect -325 -737 -291 -729
rect -325 -797 -291 -775
rect -325 -809 -291 -797
rect -325 -865 -291 -847
rect -325 -881 -291 -865
rect -17 937 17 953
rect -17 919 17 937
rect -17 869 17 881
rect -17 847 17 869
rect -17 801 17 809
rect -17 775 17 801
rect -17 733 17 737
rect -17 703 17 733
rect -17 631 17 665
rect -17 563 17 593
rect -17 559 17 563
rect -17 495 17 521
rect -17 487 17 495
rect -17 427 17 449
rect -17 415 17 427
rect -17 359 17 377
rect -17 343 17 359
rect -17 291 17 305
rect -17 271 17 291
rect -17 223 17 233
rect -17 199 17 223
rect -17 155 17 161
rect -17 127 17 155
rect -17 87 17 89
rect -17 55 17 87
rect -17 -15 17 17
rect -17 -17 17 -15
rect -17 -83 17 -55
rect -17 -89 17 -83
rect -17 -151 17 -127
rect -17 -161 17 -151
rect -17 -219 17 -199
rect -17 -233 17 -219
rect -17 -287 17 -271
rect -17 -305 17 -287
rect -17 -355 17 -343
rect -17 -377 17 -355
rect -17 -423 17 -415
rect -17 -449 17 -423
rect -17 -491 17 -487
rect -17 -521 17 -491
rect -17 -593 17 -559
rect -17 -661 17 -631
rect -17 -665 17 -661
rect -17 -729 17 -703
rect -17 -737 17 -729
rect -17 -797 17 -775
rect -17 -809 17 -797
rect -17 -865 17 -847
rect -17 -881 17 -865
rect 291 937 325 953
rect 291 919 325 937
rect 291 869 325 881
rect 291 847 325 869
rect 291 801 325 809
rect 291 775 325 801
rect 291 733 325 737
rect 291 703 325 733
rect 291 631 325 665
rect 291 563 325 593
rect 291 559 325 563
rect 291 495 325 521
rect 291 487 325 495
rect 291 427 325 449
rect 291 415 325 427
rect 291 359 325 377
rect 291 343 325 359
rect 291 291 325 305
rect 291 271 325 291
rect 291 223 325 233
rect 291 199 325 223
rect 291 155 325 161
rect 291 127 325 155
rect 291 87 325 89
rect 291 55 325 87
rect 291 -15 325 17
rect 291 -17 325 -15
rect 291 -83 325 -55
rect 291 -89 325 -83
rect 291 -151 325 -127
rect 291 -161 325 -151
rect 291 -219 325 -199
rect 291 -233 325 -219
rect 291 -287 325 -271
rect 291 -305 325 -287
rect 291 -355 325 -343
rect 291 -377 325 -355
rect 291 -423 325 -415
rect 291 -449 325 -423
rect 291 -491 325 -487
rect 291 -521 325 -491
rect 291 -593 325 -559
rect 291 -661 325 -631
rect 291 -665 325 -661
rect 291 -729 325 -703
rect 291 -737 325 -729
rect 291 -797 325 -775
rect 291 -809 325 -797
rect 291 -865 325 -847
rect 291 -881 325 -865
rect 599 937 633 953
rect 599 919 633 937
rect 599 869 633 881
rect 599 847 633 869
rect 599 801 633 809
rect 599 775 633 801
rect 599 733 633 737
rect 599 703 633 733
rect 599 631 633 665
rect 599 563 633 593
rect 599 559 633 563
rect 599 495 633 521
rect 599 487 633 495
rect 599 427 633 449
rect 599 415 633 427
rect 599 359 633 377
rect 599 343 633 359
rect 599 291 633 305
rect 599 271 633 291
rect 599 223 633 233
rect 599 199 633 223
rect 599 155 633 161
rect 599 127 633 155
rect 599 87 633 89
rect 599 55 633 87
rect 599 -15 633 17
rect 599 -17 633 -15
rect 599 -83 633 -55
rect 599 -89 633 -83
rect 599 -151 633 -127
rect 599 -161 633 -151
rect 599 -219 633 -199
rect 599 -233 633 -219
rect 599 -287 633 -271
rect 599 -305 633 -287
rect 599 -355 633 -343
rect 599 -377 633 -355
rect 599 -423 633 -415
rect 599 -449 633 -423
rect 599 -491 633 -487
rect 599 -521 633 -491
rect 599 -593 633 -559
rect 599 -661 633 -631
rect 599 -665 633 -661
rect 599 -729 633 -703
rect 599 -737 633 -729
rect 599 -797 633 -775
rect 599 -809 633 -797
rect 599 -865 633 -847
rect 599 -881 633 -865
rect 907 937 941 953
rect 907 919 941 937
rect 907 869 941 881
rect 907 847 941 869
rect 907 801 941 809
rect 907 775 941 801
rect 907 733 941 737
rect 907 703 941 733
rect 907 631 941 665
rect 907 563 941 593
rect 907 559 941 563
rect 907 495 941 521
rect 907 487 941 495
rect 907 427 941 449
rect 907 415 941 427
rect 907 359 941 377
rect 907 343 941 359
rect 907 291 941 305
rect 907 271 941 291
rect 907 223 941 233
rect 907 199 941 223
rect 907 155 941 161
rect 907 127 941 155
rect 907 87 941 89
rect 907 55 941 87
rect 907 -15 941 17
rect 907 -17 941 -15
rect 907 -83 941 -55
rect 907 -89 941 -83
rect 907 -151 941 -127
rect 907 -161 941 -151
rect 907 -219 941 -199
rect 907 -233 941 -219
rect 907 -287 941 -271
rect 907 -305 941 -287
rect 907 -355 941 -343
rect 907 -377 941 -355
rect 907 -423 941 -415
rect 907 -449 941 -423
rect 907 -491 941 -487
rect 907 -521 941 -491
rect 907 -593 941 -559
rect 907 -661 941 -631
rect 907 -665 941 -661
rect 907 -729 941 -703
rect 907 -737 941 -729
rect 907 -797 941 -775
rect 907 -809 941 -797
rect 907 -865 941 -847
rect 907 -881 941 -865
rect 1215 937 1249 953
rect 1215 919 1249 937
rect 1215 869 1249 881
rect 1215 847 1249 869
rect 1215 801 1249 809
rect 1215 775 1249 801
rect 1215 733 1249 737
rect 1215 703 1249 733
rect 1215 631 1249 665
rect 1215 563 1249 593
rect 1215 559 1249 563
rect 1215 495 1249 521
rect 1215 487 1249 495
rect 1215 427 1249 449
rect 1215 415 1249 427
rect 1215 359 1249 377
rect 1215 343 1249 359
rect 1215 291 1249 305
rect 1215 271 1249 291
rect 1215 223 1249 233
rect 1215 199 1249 223
rect 1215 155 1249 161
rect 1215 127 1249 155
rect 1215 87 1249 89
rect 1215 55 1249 87
rect 1215 -15 1249 17
rect 1215 -17 1249 -15
rect 1215 -83 1249 -55
rect 1215 -89 1249 -83
rect 1215 -151 1249 -127
rect 1215 -161 1249 -151
rect 1215 -219 1249 -199
rect 1215 -233 1249 -219
rect 1215 -287 1249 -271
rect 1215 -305 1249 -287
rect 1215 -355 1249 -343
rect 1215 -377 1249 -355
rect 1215 -423 1249 -415
rect 1215 -449 1249 -423
rect 1215 -491 1249 -487
rect 1215 -521 1249 -491
rect 1215 -593 1249 -559
rect 1215 -661 1249 -631
rect 1215 -665 1249 -661
rect 1215 -729 1249 -703
rect 1215 -737 1249 -729
rect 1215 -797 1249 -775
rect 1215 -809 1249 -797
rect 1215 -865 1249 -847
rect 1215 -881 1249 -865
rect 1523 937 1557 953
rect 1523 919 1557 937
rect 1523 869 1557 881
rect 1523 847 1557 869
rect 1523 801 1557 809
rect 1523 775 1557 801
rect 1523 733 1557 737
rect 1523 703 1557 733
rect 1523 631 1557 665
rect 1523 563 1557 593
rect 1523 559 1557 563
rect 1523 495 1557 521
rect 1523 487 1557 495
rect 1523 427 1557 449
rect 1523 415 1557 427
rect 1523 359 1557 377
rect 1523 343 1557 359
rect 1523 291 1557 305
rect 1523 271 1557 291
rect 1523 223 1557 233
rect 1523 199 1557 223
rect 1523 155 1557 161
rect 1523 127 1557 155
rect 1523 87 1557 89
rect 1523 55 1557 87
rect 1523 -15 1557 17
rect 1523 -17 1557 -15
rect 1523 -83 1557 -55
rect 1523 -89 1557 -83
rect 1523 -151 1557 -127
rect 1523 -161 1557 -151
rect 1523 -219 1557 -199
rect 1523 -233 1557 -219
rect 1523 -287 1557 -271
rect 1523 -305 1557 -287
rect 1523 -355 1557 -343
rect 1523 -377 1557 -355
rect 1523 -423 1557 -415
rect 1523 -449 1557 -423
rect 1523 -491 1557 -487
rect 1523 -521 1557 -491
rect 1523 -593 1557 -559
rect 1523 -661 1557 -631
rect 1523 -665 1557 -661
rect 1523 -729 1557 -703
rect 1523 -737 1557 -729
rect 1523 -797 1557 -775
rect 1523 -809 1557 -797
rect 1523 -865 1557 -847
rect 1523 -881 1557 -865
rect 1831 937 1865 953
rect 1831 919 1865 937
rect 1831 869 1865 881
rect 1831 847 1865 869
rect 1831 801 1865 809
rect 1831 775 1865 801
rect 1831 733 1865 737
rect 1831 703 1865 733
rect 1831 631 1865 665
rect 1831 563 1865 593
rect 1831 559 1865 563
rect 1831 495 1865 521
rect 1831 487 1865 495
rect 1831 427 1865 449
rect 1831 415 1865 427
rect 1831 359 1865 377
rect 1831 343 1865 359
rect 1831 291 1865 305
rect 1831 271 1865 291
rect 1831 223 1865 233
rect 1831 199 1865 223
rect 1831 155 1865 161
rect 1831 127 1865 155
rect 1831 87 1865 89
rect 1831 55 1865 87
rect 1831 -15 1865 17
rect 1831 -17 1865 -15
rect 1831 -83 1865 -55
rect 1831 -89 1865 -83
rect 1831 -151 1865 -127
rect 1831 -161 1865 -151
rect 1831 -219 1865 -199
rect 1831 -233 1865 -219
rect 1831 -287 1865 -271
rect 1831 -305 1865 -287
rect 1831 -355 1865 -343
rect 1831 -377 1865 -355
rect 1831 -423 1865 -415
rect 1831 -449 1865 -423
rect 1831 -491 1865 -487
rect 1831 -521 1865 -491
rect 1831 -593 1865 -559
rect 1831 -661 1865 -631
rect 1831 -665 1865 -661
rect 1831 -729 1865 -703
rect 1831 -737 1865 -729
rect 1831 -797 1865 -775
rect 1831 -809 1865 -797
rect 1831 -865 1865 -847
rect 1831 -881 1865 -865
rect 2139 937 2173 953
rect 2139 919 2173 937
rect 2139 869 2173 881
rect 2139 847 2173 869
rect 2139 801 2173 809
rect 2139 775 2173 801
rect 2139 733 2173 737
rect 2139 703 2173 733
rect 2139 631 2173 665
rect 2139 563 2173 593
rect 2139 559 2173 563
rect 2139 495 2173 521
rect 2139 487 2173 495
rect 2139 427 2173 449
rect 2139 415 2173 427
rect 2139 359 2173 377
rect 2139 343 2173 359
rect 2139 291 2173 305
rect 2139 271 2173 291
rect 2139 223 2173 233
rect 2139 199 2173 223
rect 2139 155 2173 161
rect 2139 127 2173 155
rect 2139 87 2173 89
rect 2139 55 2173 87
rect 2139 -15 2173 17
rect 2139 -17 2173 -15
rect 2139 -83 2173 -55
rect 2139 -89 2173 -83
rect 2139 -151 2173 -127
rect 2139 -161 2173 -151
rect 2139 -219 2173 -199
rect 2139 -233 2173 -219
rect 2139 -287 2173 -271
rect 2139 -305 2173 -287
rect 2139 -355 2173 -343
rect 2139 -377 2173 -355
rect 2139 -423 2173 -415
rect 2139 -449 2173 -423
rect 2139 -491 2173 -487
rect 2139 -521 2173 -491
rect 2139 -593 2173 -559
rect 2139 -661 2173 -631
rect 2139 -665 2173 -661
rect 2139 -729 2173 -703
rect 2139 -737 2173 -729
rect 2139 -797 2173 -775
rect 2139 -809 2173 -797
rect 2139 -865 2173 -847
rect 2139 -881 2173 -865
rect 2447 937 2481 953
rect 2447 919 2481 937
rect 2447 869 2481 881
rect 2447 847 2481 869
rect 2447 801 2481 809
rect 2447 775 2481 801
rect 2447 733 2481 737
rect 2447 703 2481 733
rect 2447 631 2481 665
rect 2447 563 2481 593
rect 2447 559 2481 563
rect 2447 495 2481 521
rect 2447 487 2481 495
rect 2447 427 2481 449
rect 2447 415 2481 427
rect 2447 359 2481 377
rect 2447 343 2481 359
rect 2447 291 2481 305
rect 2447 271 2481 291
rect 2447 223 2481 233
rect 2447 199 2481 223
rect 2447 155 2481 161
rect 2447 127 2481 155
rect 2447 87 2481 89
rect 2447 55 2481 87
rect 2447 -15 2481 17
rect 2447 -17 2481 -15
rect 2447 -83 2481 -55
rect 2447 -89 2481 -83
rect 2447 -151 2481 -127
rect 2447 -161 2481 -151
rect 2447 -219 2481 -199
rect 2447 -233 2481 -219
rect 2447 -287 2481 -271
rect 2447 -305 2481 -287
rect 2447 -355 2481 -343
rect 2447 -377 2481 -355
rect 2447 -423 2481 -415
rect 2447 -449 2481 -423
rect 2447 -491 2481 -487
rect 2447 -521 2481 -491
rect 2447 -593 2481 -559
rect 2447 -661 2481 -631
rect 2447 -665 2481 -661
rect 2447 -729 2481 -703
rect 2447 -737 2481 -729
rect 2447 -797 2481 -775
rect 2447 -809 2481 -797
rect 2447 -865 2481 -847
rect 2447 -881 2481 -865
rect 2755 937 2789 953
rect 2755 919 2789 937
rect 2755 869 2789 881
rect 2755 847 2789 869
rect 2755 801 2789 809
rect 2755 775 2789 801
rect 2755 733 2789 737
rect 2755 703 2789 733
rect 2755 631 2789 665
rect 2755 563 2789 593
rect 2755 559 2789 563
rect 2755 495 2789 521
rect 2755 487 2789 495
rect 2755 427 2789 449
rect 2755 415 2789 427
rect 2755 359 2789 377
rect 2755 343 2789 359
rect 2755 291 2789 305
rect 2755 271 2789 291
rect 2755 223 2789 233
rect 2755 199 2789 223
rect 2755 155 2789 161
rect 2755 127 2789 155
rect 2755 87 2789 89
rect 2755 55 2789 87
rect 2755 -15 2789 17
rect 2755 -17 2789 -15
rect 2755 -83 2789 -55
rect 2755 -89 2789 -83
rect 2755 -151 2789 -127
rect 2755 -161 2789 -151
rect 2755 -219 2789 -199
rect 2755 -233 2789 -219
rect 2755 -287 2789 -271
rect 2755 -305 2789 -287
rect 2755 -355 2789 -343
rect 2755 -377 2789 -355
rect 2755 -423 2789 -415
rect 2755 -449 2789 -423
rect 2755 -491 2789 -487
rect 2755 -521 2789 -491
rect 2755 -593 2789 -559
rect 2755 -661 2789 -631
rect 2755 -665 2789 -661
rect 2755 -729 2789 -703
rect 2755 -737 2789 -729
rect 2755 -797 2789 -775
rect 2755 -809 2789 -797
rect 2755 -865 2789 -847
rect 2755 -881 2789 -865
rect -2671 -985 -2669 -951
rect -2669 -985 -2637 -951
rect -2599 -985 -2567 -951
rect -2567 -985 -2565 -951
rect -2363 -985 -2361 -951
rect -2361 -985 -2329 -951
rect -2291 -985 -2259 -951
rect -2259 -985 -2257 -951
rect -2055 -985 -2053 -951
rect -2053 -985 -2021 -951
rect -1983 -985 -1951 -951
rect -1951 -985 -1949 -951
rect -1747 -985 -1745 -951
rect -1745 -985 -1713 -951
rect -1675 -985 -1643 -951
rect -1643 -985 -1641 -951
rect -1439 -985 -1437 -951
rect -1437 -985 -1405 -951
rect -1367 -985 -1335 -951
rect -1335 -985 -1333 -951
rect -1131 -985 -1129 -951
rect -1129 -985 -1097 -951
rect -1059 -985 -1027 -951
rect -1027 -985 -1025 -951
rect -823 -985 -821 -951
rect -821 -985 -789 -951
rect -751 -985 -719 -951
rect -719 -985 -717 -951
rect -515 -985 -513 -951
rect -513 -985 -481 -951
rect -443 -985 -411 -951
rect -411 -985 -409 -951
rect -207 -985 -205 -951
rect -205 -985 -173 -951
rect -135 -985 -103 -951
rect -103 -985 -101 -951
rect 101 -985 103 -951
rect 103 -985 135 -951
rect 173 -985 205 -951
rect 205 -985 207 -951
rect 409 -985 411 -951
rect 411 -985 443 -951
rect 481 -985 513 -951
rect 513 -985 515 -951
rect 717 -985 719 -951
rect 719 -985 751 -951
rect 789 -985 821 -951
rect 821 -985 823 -951
rect 1025 -985 1027 -951
rect 1027 -985 1059 -951
rect 1097 -985 1129 -951
rect 1129 -985 1131 -951
rect 1333 -985 1335 -951
rect 1335 -985 1367 -951
rect 1405 -985 1437 -951
rect 1437 -985 1439 -951
rect 1641 -985 1643 -951
rect 1643 -985 1675 -951
rect 1713 -985 1745 -951
rect 1745 -985 1747 -951
rect 1949 -985 1951 -951
rect 1951 -985 1983 -951
rect 2021 -985 2053 -951
rect 2053 -985 2055 -951
rect 2257 -985 2259 -951
rect 2259 -985 2291 -951
rect 2329 -985 2361 -951
rect 2361 -985 2363 -951
rect 2565 -985 2567 -951
rect 2567 -985 2599 -951
rect 2637 -985 2669 -951
rect 2669 -985 2671 -951
<< metal1 >>
rect -2795 953 -2749 976
rect -2795 919 -2789 953
rect -2755 919 -2749 953
rect -2795 881 -2749 919
rect -2795 847 -2789 881
rect -2755 847 -2749 881
rect -2795 809 -2749 847
rect -2795 775 -2789 809
rect -2755 775 -2749 809
rect -2795 737 -2749 775
rect -2795 703 -2789 737
rect -2755 703 -2749 737
rect -2795 665 -2749 703
rect -2795 631 -2789 665
rect -2755 631 -2749 665
rect -2795 593 -2749 631
rect -2795 559 -2789 593
rect -2755 559 -2749 593
rect -2795 521 -2749 559
rect -2795 487 -2789 521
rect -2755 487 -2749 521
rect -2795 449 -2749 487
rect -2795 415 -2789 449
rect -2755 415 -2749 449
rect -2795 377 -2749 415
rect -2795 343 -2789 377
rect -2755 343 -2749 377
rect -2795 305 -2749 343
rect -2795 271 -2789 305
rect -2755 271 -2749 305
rect -2795 233 -2749 271
rect -2795 199 -2789 233
rect -2755 199 -2749 233
rect -2795 161 -2749 199
rect -2795 127 -2789 161
rect -2755 127 -2749 161
rect -2795 89 -2749 127
rect -2795 55 -2789 89
rect -2755 55 -2749 89
rect -2795 17 -2749 55
rect -2795 -17 -2789 17
rect -2755 -17 -2749 17
rect -2795 -55 -2749 -17
rect -2795 -89 -2789 -55
rect -2755 -89 -2749 -55
rect -2795 -127 -2749 -89
rect -2795 -161 -2789 -127
rect -2755 -161 -2749 -127
rect -2795 -199 -2749 -161
rect -2795 -233 -2789 -199
rect -2755 -233 -2749 -199
rect -2795 -271 -2749 -233
rect -2795 -305 -2789 -271
rect -2755 -305 -2749 -271
rect -2795 -343 -2749 -305
rect -2795 -377 -2789 -343
rect -2755 -377 -2749 -343
rect -2795 -415 -2749 -377
rect -2795 -449 -2789 -415
rect -2755 -449 -2749 -415
rect -2795 -487 -2749 -449
rect -2795 -521 -2789 -487
rect -2755 -521 -2749 -487
rect -2795 -559 -2749 -521
rect -2795 -593 -2789 -559
rect -2755 -593 -2749 -559
rect -2795 -631 -2749 -593
rect -2795 -665 -2789 -631
rect -2755 -665 -2749 -631
rect -2795 -703 -2749 -665
rect -2795 -737 -2789 -703
rect -2755 -737 -2749 -703
rect -2795 -775 -2749 -737
rect -2795 -809 -2789 -775
rect -2755 -809 -2749 -775
rect -2795 -847 -2749 -809
rect -2795 -881 -2789 -847
rect -2755 -881 -2749 -847
rect -2795 -904 -2749 -881
rect -2487 953 -2441 976
rect -2487 919 -2481 953
rect -2447 919 -2441 953
rect -2487 881 -2441 919
rect -2487 847 -2481 881
rect -2447 847 -2441 881
rect -2487 809 -2441 847
rect -2487 775 -2481 809
rect -2447 775 -2441 809
rect -2487 737 -2441 775
rect -2487 703 -2481 737
rect -2447 703 -2441 737
rect -2487 665 -2441 703
rect -2487 631 -2481 665
rect -2447 631 -2441 665
rect -2487 593 -2441 631
rect -2487 559 -2481 593
rect -2447 559 -2441 593
rect -2487 521 -2441 559
rect -2487 487 -2481 521
rect -2447 487 -2441 521
rect -2487 449 -2441 487
rect -2487 415 -2481 449
rect -2447 415 -2441 449
rect -2487 377 -2441 415
rect -2487 343 -2481 377
rect -2447 343 -2441 377
rect -2487 305 -2441 343
rect -2487 271 -2481 305
rect -2447 271 -2441 305
rect -2487 233 -2441 271
rect -2487 199 -2481 233
rect -2447 199 -2441 233
rect -2487 161 -2441 199
rect -2487 127 -2481 161
rect -2447 127 -2441 161
rect -2487 89 -2441 127
rect -2487 55 -2481 89
rect -2447 55 -2441 89
rect -2487 17 -2441 55
rect -2487 -17 -2481 17
rect -2447 -17 -2441 17
rect -2487 -55 -2441 -17
rect -2487 -89 -2481 -55
rect -2447 -89 -2441 -55
rect -2487 -127 -2441 -89
rect -2487 -161 -2481 -127
rect -2447 -161 -2441 -127
rect -2487 -199 -2441 -161
rect -2487 -233 -2481 -199
rect -2447 -233 -2441 -199
rect -2487 -271 -2441 -233
rect -2487 -305 -2481 -271
rect -2447 -305 -2441 -271
rect -2487 -343 -2441 -305
rect -2487 -377 -2481 -343
rect -2447 -377 -2441 -343
rect -2487 -415 -2441 -377
rect -2487 -449 -2481 -415
rect -2447 -449 -2441 -415
rect -2487 -487 -2441 -449
rect -2487 -521 -2481 -487
rect -2447 -521 -2441 -487
rect -2487 -559 -2441 -521
rect -2487 -593 -2481 -559
rect -2447 -593 -2441 -559
rect -2487 -631 -2441 -593
rect -2487 -665 -2481 -631
rect -2447 -665 -2441 -631
rect -2487 -703 -2441 -665
rect -2487 -737 -2481 -703
rect -2447 -737 -2441 -703
rect -2487 -775 -2441 -737
rect -2487 -809 -2481 -775
rect -2447 -809 -2441 -775
rect -2487 -847 -2441 -809
rect -2487 -881 -2481 -847
rect -2447 -881 -2441 -847
rect -2487 -904 -2441 -881
rect -2179 953 -2133 976
rect -2179 919 -2173 953
rect -2139 919 -2133 953
rect -2179 881 -2133 919
rect -2179 847 -2173 881
rect -2139 847 -2133 881
rect -2179 809 -2133 847
rect -2179 775 -2173 809
rect -2139 775 -2133 809
rect -2179 737 -2133 775
rect -2179 703 -2173 737
rect -2139 703 -2133 737
rect -2179 665 -2133 703
rect -2179 631 -2173 665
rect -2139 631 -2133 665
rect -2179 593 -2133 631
rect -2179 559 -2173 593
rect -2139 559 -2133 593
rect -2179 521 -2133 559
rect -2179 487 -2173 521
rect -2139 487 -2133 521
rect -2179 449 -2133 487
rect -2179 415 -2173 449
rect -2139 415 -2133 449
rect -2179 377 -2133 415
rect -2179 343 -2173 377
rect -2139 343 -2133 377
rect -2179 305 -2133 343
rect -2179 271 -2173 305
rect -2139 271 -2133 305
rect -2179 233 -2133 271
rect -2179 199 -2173 233
rect -2139 199 -2133 233
rect -2179 161 -2133 199
rect -2179 127 -2173 161
rect -2139 127 -2133 161
rect -2179 89 -2133 127
rect -2179 55 -2173 89
rect -2139 55 -2133 89
rect -2179 17 -2133 55
rect -2179 -17 -2173 17
rect -2139 -17 -2133 17
rect -2179 -55 -2133 -17
rect -2179 -89 -2173 -55
rect -2139 -89 -2133 -55
rect -2179 -127 -2133 -89
rect -2179 -161 -2173 -127
rect -2139 -161 -2133 -127
rect -2179 -199 -2133 -161
rect -2179 -233 -2173 -199
rect -2139 -233 -2133 -199
rect -2179 -271 -2133 -233
rect -2179 -305 -2173 -271
rect -2139 -305 -2133 -271
rect -2179 -343 -2133 -305
rect -2179 -377 -2173 -343
rect -2139 -377 -2133 -343
rect -2179 -415 -2133 -377
rect -2179 -449 -2173 -415
rect -2139 -449 -2133 -415
rect -2179 -487 -2133 -449
rect -2179 -521 -2173 -487
rect -2139 -521 -2133 -487
rect -2179 -559 -2133 -521
rect -2179 -593 -2173 -559
rect -2139 -593 -2133 -559
rect -2179 -631 -2133 -593
rect -2179 -665 -2173 -631
rect -2139 -665 -2133 -631
rect -2179 -703 -2133 -665
rect -2179 -737 -2173 -703
rect -2139 -737 -2133 -703
rect -2179 -775 -2133 -737
rect -2179 -809 -2173 -775
rect -2139 -809 -2133 -775
rect -2179 -847 -2133 -809
rect -2179 -881 -2173 -847
rect -2139 -881 -2133 -847
rect -2179 -904 -2133 -881
rect -1871 953 -1825 976
rect -1871 919 -1865 953
rect -1831 919 -1825 953
rect -1871 881 -1825 919
rect -1871 847 -1865 881
rect -1831 847 -1825 881
rect -1871 809 -1825 847
rect -1871 775 -1865 809
rect -1831 775 -1825 809
rect -1871 737 -1825 775
rect -1871 703 -1865 737
rect -1831 703 -1825 737
rect -1871 665 -1825 703
rect -1871 631 -1865 665
rect -1831 631 -1825 665
rect -1871 593 -1825 631
rect -1871 559 -1865 593
rect -1831 559 -1825 593
rect -1871 521 -1825 559
rect -1871 487 -1865 521
rect -1831 487 -1825 521
rect -1871 449 -1825 487
rect -1871 415 -1865 449
rect -1831 415 -1825 449
rect -1871 377 -1825 415
rect -1871 343 -1865 377
rect -1831 343 -1825 377
rect -1871 305 -1825 343
rect -1871 271 -1865 305
rect -1831 271 -1825 305
rect -1871 233 -1825 271
rect -1871 199 -1865 233
rect -1831 199 -1825 233
rect -1871 161 -1825 199
rect -1871 127 -1865 161
rect -1831 127 -1825 161
rect -1871 89 -1825 127
rect -1871 55 -1865 89
rect -1831 55 -1825 89
rect -1871 17 -1825 55
rect -1871 -17 -1865 17
rect -1831 -17 -1825 17
rect -1871 -55 -1825 -17
rect -1871 -89 -1865 -55
rect -1831 -89 -1825 -55
rect -1871 -127 -1825 -89
rect -1871 -161 -1865 -127
rect -1831 -161 -1825 -127
rect -1871 -199 -1825 -161
rect -1871 -233 -1865 -199
rect -1831 -233 -1825 -199
rect -1871 -271 -1825 -233
rect -1871 -305 -1865 -271
rect -1831 -305 -1825 -271
rect -1871 -343 -1825 -305
rect -1871 -377 -1865 -343
rect -1831 -377 -1825 -343
rect -1871 -415 -1825 -377
rect -1871 -449 -1865 -415
rect -1831 -449 -1825 -415
rect -1871 -487 -1825 -449
rect -1871 -521 -1865 -487
rect -1831 -521 -1825 -487
rect -1871 -559 -1825 -521
rect -1871 -593 -1865 -559
rect -1831 -593 -1825 -559
rect -1871 -631 -1825 -593
rect -1871 -665 -1865 -631
rect -1831 -665 -1825 -631
rect -1871 -703 -1825 -665
rect -1871 -737 -1865 -703
rect -1831 -737 -1825 -703
rect -1871 -775 -1825 -737
rect -1871 -809 -1865 -775
rect -1831 -809 -1825 -775
rect -1871 -847 -1825 -809
rect -1871 -881 -1865 -847
rect -1831 -881 -1825 -847
rect -1871 -904 -1825 -881
rect -1563 953 -1517 976
rect -1563 919 -1557 953
rect -1523 919 -1517 953
rect -1563 881 -1517 919
rect -1563 847 -1557 881
rect -1523 847 -1517 881
rect -1563 809 -1517 847
rect -1563 775 -1557 809
rect -1523 775 -1517 809
rect -1563 737 -1517 775
rect -1563 703 -1557 737
rect -1523 703 -1517 737
rect -1563 665 -1517 703
rect -1563 631 -1557 665
rect -1523 631 -1517 665
rect -1563 593 -1517 631
rect -1563 559 -1557 593
rect -1523 559 -1517 593
rect -1563 521 -1517 559
rect -1563 487 -1557 521
rect -1523 487 -1517 521
rect -1563 449 -1517 487
rect -1563 415 -1557 449
rect -1523 415 -1517 449
rect -1563 377 -1517 415
rect -1563 343 -1557 377
rect -1523 343 -1517 377
rect -1563 305 -1517 343
rect -1563 271 -1557 305
rect -1523 271 -1517 305
rect -1563 233 -1517 271
rect -1563 199 -1557 233
rect -1523 199 -1517 233
rect -1563 161 -1517 199
rect -1563 127 -1557 161
rect -1523 127 -1517 161
rect -1563 89 -1517 127
rect -1563 55 -1557 89
rect -1523 55 -1517 89
rect -1563 17 -1517 55
rect -1563 -17 -1557 17
rect -1523 -17 -1517 17
rect -1563 -55 -1517 -17
rect -1563 -89 -1557 -55
rect -1523 -89 -1517 -55
rect -1563 -127 -1517 -89
rect -1563 -161 -1557 -127
rect -1523 -161 -1517 -127
rect -1563 -199 -1517 -161
rect -1563 -233 -1557 -199
rect -1523 -233 -1517 -199
rect -1563 -271 -1517 -233
rect -1563 -305 -1557 -271
rect -1523 -305 -1517 -271
rect -1563 -343 -1517 -305
rect -1563 -377 -1557 -343
rect -1523 -377 -1517 -343
rect -1563 -415 -1517 -377
rect -1563 -449 -1557 -415
rect -1523 -449 -1517 -415
rect -1563 -487 -1517 -449
rect -1563 -521 -1557 -487
rect -1523 -521 -1517 -487
rect -1563 -559 -1517 -521
rect -1563 -593 -1557 -559
rect -1523 -593 -1517 -559
rect -1563 -631 -1517 -593
rect -1563 -665 -1557 -631
rect -1523 -665 -1517 -631
rect -1563 -703 -1517 -665
rect -1563 -737 -1557 -703
rect -1523 -737 -1517 -703
rect -1563 -775 -1517 -737
rect -1563 -809 -1557 -775
rect -1523 -809 -1517 -775
rect -1563 -847 -1517 -809
rect -1563 -881 -1557 -847
rect -1523 -881 -1517 -847
rect -1563 -904 -1517 -881
rect -1255 953 -1209 976
rect -1255 919 -1249 953
rect -1215 919 -1209 953
rect -1255 881 -1209 919
rect -1255 847 -1249 881
rect -1215 847 -1209 881
rect -1255 809 -1209 847
rect -1255 775 -1249 809
rect -1215 775 -1209 809
rect -1255 737 -1209 775
rect -1255 703 -1249 737
rect -1215 703 -1209 737
rect -1255 665 -1209 703
rect -1255 631 -1249 665
rect -1215 631 -1209 665
rect -1255 593 -1209 631
rect -1255 559 -1249 593
rect -1215 559 -1209 593
rect -1255 521 -1209 559
rect -1255 487 -1249 521
rect -1215 487 -1209 521
rect -1255 449 -1209 487
rect -1255 415 -1249 449
rect -1215 415 -1209 449
rect -1255 377 -1209 415
rect -1255 343 -1249 377
rect -1215 343 -1209 377
rect -1255 305 -1209 343
rect -1255 271 -1249 305
rect -1215 271 -1209 305
rect -1255 233 -1209 271
rect -1255 199 -1249 233
rect -1215 199 -1209 233
rect -1255 161 -1209 199
rect -1255 127 -1249 161
rect -1215 127 -1209 161
rect -1255 89 -1209 127
rect -1255 55 -1249 89
rect -1215 55 -1209 89
rect -1255 17 -1209 55
rect -1255 -17 -1249 17
rect -1215 -17 -1209 17
rect -1255 -55 -1209 -17
rect -1255 -89 -1249 -55
rect -1215 -89 -1209 -55
rect -1255 -127 -1209 -89
rect -1255 -161 -1249 -127
rect -1215 -161 -1209 -127
rect -1255 -199 -1209 -161
rect -1255 -233 -1249 -199
rect -1215 -233 -1209 -199
rect -1255 -271 -1209 -233
rect -1255 -305 -1249 -271
rect -1215 -305 -1209 -271
rect -1255 -343 -1209 -305
rect -1255 -377 -1249 -343
rect -1215 -377 -1209 -343
rect -1255 -415 -1209 -377
rect -1255 -449 -1249 -415
rect -1215 -449 -1209 -415
rect -1255 -487 -1209 -449
rect -1255 -521 -1249 -487
rect -1215 -521 -1209 -487
rect -1255 -559 -1209 -521
rect -1255 -593 -1249 -559
rect -1215 -593 -1209 -559
rect -1255 -631 -1209 -593
rect -1255 -665 -1249 -631
rect -1215 -665 -1209 -631
rect -1255 -703 -1209 -665
rect -1255 -737 -1249 -703
rect -1215 -737 -1209 -703
rect -1255 -775 -1209 -737
rect -1255 -809 -1249 -775
rect -1215 -809 -1209 -775
rect -1255 -847 -1209 -809
rect -1255 -881 -1249 -847
rect -1215 -881 -1209 -847
rect -1255 -904 -1209 -881
rect -947 953 -901 976
rect -947 919 -941 953
rect -907 919 -901 953
rect -947 881 -901 919
rect -947 847 -941 881
rect -907 847 -901 881
rect -947 809 -901 847
rect -947 775 -941 809
rect -907 775 -901 809
rect -947 737 -901 775
rect -947 703 -941 737
rect -907 703 -901 737
rect -947 665 -901 703
rect -947 631 -941 665
rect -907 631 -901 665
rect -947 593 -901 631
rect -947 559 -941 593
rect -907 559 -901 593
rect -947 521 -901 559
rect -947 487 -941 521
rect -907 487 -901 521
rect -947 449 -901 487
rect -947 415 -941 449
rect -907 415 -901 449
rect -947 377 -901 415
rect -947 343 -941 377
rect -907 343 -901 377
rect -947 305 -901 343
rect -947 271 -941 305
rect -907 271 -901 305
rect -947 233 -901 271
rect -947 199 -941 233
rect -907 199 -901 233
rect -947 161 -901 199
rect -947 127 -941 161
rect -907 127 -901 161
rect -947 89 -901 127
rect -947 55 -941 89
rect -907 55 -901 89
rect -947 17 -901 55
rect -947 -17 -941 17
rect -907 -17 -901 17
rect -947 -55 -901 -17
rect -947 -89 -941 -55
rect -907 -89 -901 -55
rect -947 -127 -901 -89
rect -947 -161 -941 -127
rect -907 -161 -901 -127
rect -947 -199 -901 -161
rect -947 -233 -941 -199
rect -907 -233 -901 -199
rect -947 -271 -901 -233
rect -947 -305 -941 -271
rect -907 -305 -901 -271
rect -947 -343 -901 -305
rect -947 -377 -941 -343
rect -907 -377 -901 -343
rect -947 -415 -901 -377
rect -947 -449 -941 -415
rect -907 -449 -901 -415
rect -947 -487 -901 -449
rect -947 -521 -941 -487
rect -907 -521 -901 -487
rect -947 -559 -901 -521
rect -947 -593 -941 -559
rect -907 -593 -901 -559
rect -947 -631 -901 -593
rect -947 -665 -941 -631
rect -907 -665 -901 -631
rect -947 -703 -901 -665
rect -947 -737 -941 -703
rect -907 -737 -901 -703
rect -947 -775 -901 -737
rect -947 -809 -941 -775
rect -907 -809 -901 -775
rect -947 -847 -901 -809
rect -947 -881 -941 -847
rect -907 -881 -901 -847
rect -947 -904 -901 -881
rect -639 953 -593 976
rect -639 919 -633 953
rect -599 919 -593 953
rect -639 881 -593 919
rect -639 847 -633 881
rect -599 847 -593 881
rect -639 809 -593 847
rect -639 775 -633 809
rect -599 775 -593 809
rect -639 737 -593 775
rect -639 703 -633 737
rect -599 703 -593 737
rect -639 665 -593 703
rect -639 631 -633 665
rect -599 631 -593 665
rect -639 593 -593 631
rect -639 559 -633 593
rect -599 559 -593 593
rect -639 521 -593 559
rect -639 487 -633 521
rect -599 487 -593 521
rect -639 449 -593 487
rect -639 415 -633 449
rect -599 415 -593 449
rect -639 377 -593 415
rect -639 343 -633 377
rect -599 343 -593 377
rect -639 305 -593 343
rect -639 271 -633 305
rect -599 271 -593 305
rect -639 233 -593 271
rect -639 199 -633 233
rect -599 199 -593 233
rect -639 161 -593 199
rect -639 127 -633 161
rect -599 127 -593 161
rect -639 89 -593 127
rect -639 55 -633 89
rect -599 55 -593 89
rect -639 17 -593 55
rect -639 -17 -633 17
rect -599 -17 -593 17
rect -639 -55 -593 -17
rect -639 -89 -633 -55
rect -599 -89 -593 -55
rect -639 -127 -593 -89
rect -639 -161 -633 -127
rect -599 -161 -593 -127
rect -639 -199 -593 -161
rect -639 -233 -633 -199
rect -599 -233 -593 -199
rect -639 -271 -593 -233
rect -639 -305 -633 -271
rect -599 -305 -593 -271
rect -639 -343 -593 -305
rect -639 -377 -633 -343
rect -599 -377 -593 -343
rect -639 -415 -593 -377
rect -639 -449 -633 -415
rect -599 -449 -593 -415
rect -639 -487 -593 -449
rect -639 -521 -633 -487
rect -599 -521 -593 -487
rect -639 -559 -593 -521
rect -639 -593 -633 -559
rect -599 -593 -593 -559
rect -639 -631 -593 -593
rect -639 -665 -633 -631
rect -599 -665 -593 -631
rect -639 -703 -593 -665
rect -639 -737 -633 -703
rect -599 -737 -593 -703
rect -639 -775 -593 -737
rect -639 -809 -633 -775
rect -599 -809 -593 -775
rect -639 -847 -593 -809
rect -639 -881 -633 -847
rect -599 -881 -593 -847
rect -639 -904 -593 -881
rect -331 953 -285 976
rect -331 919 -325 953
rect -291 919 -285 953
rect -331 881 -285 919
rect -331 847 -325 881
rect -291 847 -285 881
rect -331 809 -285 847
rect -331 775 -325 809
rect -291 775 -285 809
rect -331 737 -285 775
rect -331 703 -325 737
rect -291 703 -285 737
rect -331 665 -285 703
rect -331 631 -325 665
rect -291 631 -285 665
rect -331 593 -285 631
rect -331 559 -325 593
rect -291 559 -285 593
rect -331 521 -285 559
rect -331 487 -325 521
rect -291 487 -285 521
rect -331 449 -285 487
rect -331 415 -325 449
rect -291 415 -285 449
rect -331 377 -285 415
rect -331 343 -325 377
rect -291 343 -285 377
rect -331 305 -285 343
rect -331 271 -325 305
rect -291 271 -285 305
rect -331 233 -285 271
rect -331 199 -325 233
rect -291 199 -285 233
rect -331 161 -285 199
rect -331 127 -325 161
rect -291 127 -285 161
rect -331 89 -285 127
rect -331 55 -325 89
rect -291 55 -285 89
rect -331 17 -285 55
rect -331 -17 -325 17
rect -291 -17 -285 17
rect -331 -55 -285 -17
rect -331 -89 -325 -55
rect -291 -89 -285 -55
rect -331 -127 -285 -89
rect -331 -161 -325 -127
rect -291 -161 -285 -127
rect -331 -199 -285 -161
rect -331 -233 -325 -199
rect -291 -233 -285 -199
rect -331 -271 -285 -233
rect -331 -305 -325 -271
rect -291 -305 -285 -271
rect -331 -343 -285 -305
rect -331 -377 -325 -343
rect -291 -377 -285 -343
rect -331 -415 -285 -377
rect -331 -449 -325 -415
rect -291 -449 -285 -415
rect -331 -487 -285 -449
rect -331 -521 -325 -487
rect -291 -521 -285 -487
rect -331 -559 -285 -521
rect -331 -593 -325 -559
rect -291 -593 -285 -559
rect -331 -631 -285 -593
rect -331 -665 -325 -631
rect -291 -665 -285 -631
rect -331 -703 -285 -665
rect -331 -737 -325 -703
rect -291 -737 -285 -703
rect -331 -775 -285 -737
rect -331 -809 -325 -775
rect -291 -809 -285 -775
rect -331 -847 -285 -809
rect -331 -881 -325 -847
rect -291 -881 -285 -847
rect -331 -904 -285 -881
rect -23 953 23 976
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -904 23 -881
rect 285 953 331 976
rect 285 919 291 953
rect 325 919 331 953
rect 285 881 331 919
rect 285 847 291 881
rect 325 847 331 881
rect 285 809 331 847
rect 285 775 291 809
rect 325 775 331 809
rect 285 737 331 775
rect 285 703 291 737
rect 325 703 331 737
rect 285 665 331 703
rect 285 631 291 665
rect 325 631 331 665
rect 285 593 331 631
rect 285 559 291 593
rect 325 559 331 593
rect 285 521 331 559
rect 285 487 291 521
rect 325 487 331 521
rect 285 449 331 487
rect 285 415 291 449
rect 325 415 331 449
rect 285 377 331 415
rect 285 343 291 377
rect 325 343 331 377
rect 285 305 331 343
rect 285 271 291 305
rect 325 271 331 305
rect 285 233 331 271
rect 285 199 291 233
rect 325 199 331 233
rect 285 161 331 199
rect 285 127 291 161
rect 325 127 331 161
rect 285 89 331 127
rect 285 55 291 89
rect 325 55 331 89
rect 285 17 331 55
rect 285 -17 291 17
rect 325 -17 331 17
rect 285 -55 331 -17
rect 285 -89 291 -55
rect 325 -89 331 -55
rect 285 -127 331 -89
rect 285 -161 291 -127
rect 325 -161 331 -127
rect 285 -199 331 -161
rect 285 -233 291 -199
rect 325 -233 331 -199
rect 285 -271 331 -233
rect 285 -305 291 -271
rect 325 -305 331 -271
rect 285 -343 331 -305
rect 285 -377 291 -343
rect 325 -377 331 -343
rect 285 -415 331 -377
rect 285 -449 291 -415
rect 325 -449 331 -415
rect 285 -487 331 -449
rect 285 -521 291 -487
rect 325 -521 331 -487
rect 285 -559 331 -521
rect 285 -593 291 -559
rect 325 -593 331 -559
rect 285 -631 331 -593
rect 285 -665 291 -631
rect 325 -665 331 -631
rect 285 -703 331 -665
rect 285 -737 291 -703
rect 325 -737 331 -703
rect 285 -775 331 -737
rect 285 -809 291 -775
rect 325 -809 331 -775
rect 285 -847 331 -809
rect 285 -881 291 -847
rect 325 -881 331 -847
rect 285 -904 331 -881
rect 593 953 639 976
rect 593 919 599 953
rect 633 919 639 953
rect 593 881 639 919
rect 593 847 599 881
rect 633 847 639 881
rect 593 809 639 847
rect 593 775 599 809
rect 633 775 639 809
rect 593 737 639 775
rect 593 703 599 737
rect 633 703 639 737
rect 593 665 639 703
rect 593 631 599 665
rect 633 631 639 665
rect 593 593 639 631
rect 593 559 599 593
rect 633 559 639 593
rect 593 521 639 559
rect 593 487 599 521
rect 633 487 639 521
rect 593 449 639 487
rect 593 415 599 449
rect 633 415 639 449
rect 593 377 639 415
rect 593 343 599 377
rect 633 343 639 377
rect 593 305 639 343
rect 593 271 599 305
rect 633 271 639 305
rect 593 233 639 271
rect 593 199 599 233
rect 633 199 639 233
rect 593 161 639 199
rect 593 127 599 161
rect 633 127 639 161
rect 593 89 639 127
rect 593 55 599 89
rect 633 55 639 89
rect 593 17 639 55
rect 593 -17 599 17
rect 633 -17 639 17
rect 593 -55 639 -17
rect 593 -89 599 -55
rect 633 -89 639 -55
rect 593 -127 639 -89
rect 593 -161 599 -127
rect 633 -161 639 -127
rect 593 -199 639 -161
rect 593 -233 599 -199
rect 633 -233 639 -199
rect 593 -271 639 -233
rect 593 -305 599 -271
rect 633 -305 639 -271
rect 593 -343 639 -305
rect 593 -377 599 -343
rect 633 -377 639 -343
rect 593 -415 639 -377
rect 593 -449 599 -415
rect 633 -449 639 -415
rect 593 -487 639 -449
rect 593 -521 599 -487
rect 633 -521 639 -487
rect 593 -559 639 -521
rect 593 -593 599 -559
rect 633 -593 639 -559
rect 593 -631 639 -593
rect 593 -665 599 -631
rect 633 -665 639 -631
rect 593 -703 639 -665
rect 593 -737 599 -703
rect 633 -737 639 -703
rect 593 -775 639 -737
rect 593 -809 599 -775
rect 633 -809 639 -775
rect 593 -847 639 -809
rect 593 -881 599 -847
rect 633 -881 639 -847
rect 593 -904 639 -881
rect 901 953 947 976
rect 901 919 907 953
rect 941 919 947 953
rect 901 881 947 919
rect 901 847 907 881
rect 941 847 947 881
rect 901 809 947 847
rect 901 775 907 809
rect 941 775 947 809
rect 901 737 947 775
rect 901 703 907 737
rect 941 703 947 737
rect 901 665 947 703
rect 901 631 907 665
rect 941 631 947 665
rect 901 593 947 631
rect 901 559 907 593
rect 941 559 947 593
rect 901 521 947 559
rect 901 487 907 521
rect 941 487 947 521
rect 901 449 947 487
rect 901 415 907 449
rect 941 415 947 449
rect 901 377 947 415
rect 901 343 907 377
rect 941 343 947 377
rect 901 305 947 343
rect 901 271 907 305
rect 941 271 947 305
rect 901 233 947 271
rect 901 199 907 233
rect 941 199 947 233
rect 901 161 947 199
rect 901 127 907 161
rect 941 127 947 161
rect 901 89 947 127
rect 901 55 907 89
rect 941 55 947 89
rect 901 17 947 55
rect 901 -17 907 17
rect 941 -17 947 17
rect 901 -55 947 -17
rect 901 -89 907 -55
rect 941 -89 947 -55
rect 901 -127 947 -89
rect 901 -161 907 -127
rect 941 -161 947 -127
rect 901 -199 947 -161
rect 901 -233 907 -199
rect 941 -233 947 -199
rect 901 -271 947 -233
rect 901 -305 907 -271
rect 941 -305 947 -271
rect 901 -343 947 -305
rect 901 -377 907 -343
rect 941 -377 947 -343
rect 901 -415 947 -377
rect 901 -449 907 -415
rect 941 -449 947 -415
rect 901 -487 947 -449
rect 901 -521 907 -487
rect 941 -521 947 -487
rect 901 -559 947 -521
rect 901 -593 907 -559
rect 941 -593 947 -559
rect 901 -631 947 -593
rect 901 -665 907 -631
rect 941 -665 947 -631
rect 901 -703 947 -665
rect 901 -737 907 -703
rect 941 -737 947 -703
rect 901 -775 947 -737
rect 901 -809 907 -775
rect 941 -809 947 -775
rect 901 -847 947 -809
rect 901 -881 907 -847
rect 941 -881 947 -847
rect 901 -904 947 -881
rect 1209 953 1255 976
rect 1209 919 1215 953
rect 1249 919 1255 953
rect 1209 881 1255 919
rect 1209 847 1215 881
rect 1249 847 1255 881
rect 1209 809 1255 847
rect 1209 775 1215 809
rect 1249 775 1255 809
rect 1209 737 1255 775
rect 1209 703 1215 737
rect 1249 703 1255 737
rect 1209 665 1255 703
rect 1209 631 1215 665
rect 1249 631 1255 665
rect 1209 593 1255 631
rect 1209 559 1215 593
rect 1249 559 1255 593
rect 1209 521 1255 559
rect 1209 487 1215 521
rect 1249 487 1255 521
rect 1209 449 1255 487
rect 1209 415 1215 449
rect 1249 415 1255 449
rect 1209 377 1255 415
rect 1209 343 1215 377
rect 1249 343 1255 377
rect 1209 305 1255 343
rect 1209 271 1215 305
rect 1249 271 1255 305
rect 1209 233 1255 271
rect 1209 199 1215 233
rect 1249 199 1255 233
rect 1209 161 1255 199
rect 1209 127 1215 161
rect 1249 127 1255 161
rect 1209 89 1255 127
rect 1209 55 1215 89
rect 1249 55 1255 89
rect 1209 17 1255 55
rect 1209 -17 1215 17
rect 1249 -17 1255 17
rect 1209 -55 1255 -17
rect 1209 -89 1215 -55
rect 1249 -89 1255 -55
rect 1209 -127 1255 -89
rect 1209 -161 1215 -127
rect 1249 -161 1255 -127
rect 1209 -199 1255 -161
rect 1209 -233 1215 -199
rect 1249 -233 1255 -199
rect 1209 -271 1255 -233
rect 1209 -305 1215 -271
rect 1249 -305 1255 -271
rect 1209 -343 1255 -305
rect 1209 -377 1215 -343
rect 1249 -377 1255 -343
rect 1209 -415 1255 -377
rect 1209 -449 1215 -415
rect 1249 -449 1255 -415
rect 1209 -487 1255 -449
rect 1209 -521 1215 -487
rect 1249 -521 1255 -487
rect 1209 -559 1255 -521
rect 1209 -593 1215 -559
rect 1249 -593 1255 -559
rect 1209 -631 1255 -593
rect 1209 -665 1215 -631
rect 1249 -665 1255 -631
rect 1209 -703 1255 -665
rect 1209 -737 1215 -703
rect 1249 -737 1255 -703
rect 1209 -775 1255 -737
rect 1209 -809 1215 -775
rect 1249 -809 1255 -775
rect 1209 -847 1255 -809
rect 1209 -881 1215 -847
rect 1249 -881 1255 -847
rect 1209 -904 1255 -881
rect 1517 953 1563 976
rect 1517 919 1523 953
rect 1557 919 1563 953
rect 1517 881 1563 919
rect 1517 847 1523 881
rect 1557 847 1563 881
rect 1517 809 1563 847
rect 1517 775 1523 809
rect 1557 775 1563 809
rect 1517 737 1563 775
rect 1517 703 1523 737
rect 1557 703 1563 737
rect 1517 665 1563 703
rect 1517 631 1523 665
rect 1557 631 1563 665
rect 1517 593 1563 631
rect 1517 559 1523 593
rect 1557 559 1563 593
rect 1517 521 1563 559
rect 1517 487 1523 521
rect 1557 487 1563 521
rect 1517 449 1563 487
rect 1517 415 1523 449
rect 1557 415 1563 449
rect 1517 377 1563 415
rect 1517 343 1523 377
rect 1557 343 1563 377
rect 1517 305 1563 343
rect 1517 271 1523 305
rect 1557 271 1563 305
rect 1517 233 1563 271
rect 1517 199 1523 233
rect 1557 199 1563 233
rect 1517 161 1563 199
rect 1517 127 1523 161
rect 1557 127 1563 161
rect 1517 89 1563 127
rect 1517 55 1523 89
rect 1557 55 1563 89
rect 1517 17 1563 55
rect 1517 -17 1523 17
rect 1557 -17 1563 17
rect 1517 -55 1563 -17
rect 1517 -89 1523 -55
rect 1557 -89 1563 -55
rect 1517 -127 1563 -89
rect 1517 -161 1523 -127
rect 1557 -161 1563 -127
rect 1517 -199 1563 -161
rect 1517 -233 1523 -199
rect 1557 -233 1563 -199
rect 1517 -271 1563 -233
rect 1517 -305 1523 -271
rect 1557 -305 1563 -271
rect 1517 -343 1563 -305
rect 1517 -377 1523 -343
rect 1557 -377 1563 -343
rect 1517 -415 1563 -377
rect 1517 -449 1523 -415
rect 1557 -449 1563 -415
rect 1517 -487 1563 -449
rect 1517 -521 1523 -487
rect 1557 -521 1563 -487
rect 1517 -559 1563 -521
rect 1517 -593 1523 -559
rect 1557 -593 1563 -559
rect 1517 -631 1563 -593
rect 1517 -665 1523 -631
rect 1557 -665 1563 -631
rect 1517 -703 1563 -665
rect 1517 -737 1523 -703
rect 1557 -737 1563 -703
rect 1517 -775 1563 -737
rect 1517 -809 1523 -775
rect 1557 -809 1563 -775
rect 1517 -847 1563 -809
rect 1517 -881 1523 -847
rect 1557 -881 1563 -847
rect 1517 -904 1563 -881
rect 1825 953 1871 976
rect 1825 919 1831 953
rect 1865 919 1871 953
rect 1825 881 1871 919
rect 1825 847 1831 881
rect 1865 847 1871 881
rect 1825 809 1871 847
rect 1825 775 1831 809
rect 1865 775 1871 809
rect 1825 737 1871 775
rect 1825 703 1831 737
rect 1865 703 1871 737
rect 1825 665 1871 703
rect 1825 631 1831 665
rect 1865 631 1871 665
rect 1825 593 1871 631
rect 1825 559 1831 593
rect 1865 559 1871 593
rect 1825 521 1871 559
rect 1825 487 1831 521
rect 1865 487 1871 521
rect 1825 449 1871 487
rect 1825 415 1831 449
rect 1865 415 1871 449
rect 1825 377 1871 415
rect 1825 343 1831 377
rect 1865 343 1871 377
rect 1825 305 1871 343
rect 1825 271 1831 305
rect 1865 271 1871 305
rect 1825 233 1871 271
rect 1825 199 1831 233
rect 1865 199 1871 233
rect 1825 161 1871 199
rect 1825 127 1831 161
rect 1865 127 1871 161
rect 1825 89 1871 127
rect 1825 55 1831 89
rect 1865 55 1871 89
rect 1825 17 1871 55
rect 1825 -17 1831 17
rect 1865 -17 1871 17
rect 1825 -55 1871 -17
rect 1825 -89 1831 -55
rect 1865 -89 1871 -55
rect 1825 -127 1871 -89
rect 1825 -161 1831 -127
rect 1865 -161 1871 -127
rect 1825 -199 1871 -161
rect 1825 -233 1831 -199
rect 1865 -233 1871 -199
rect 1825 -271 1871 -233
rect 1825 -305 1831 -271
rect 1865 -305 1871 -271
rect 1825 -343 1871 -305
rect 1825 -377 1831 -343
rect 1865 -377 1871 -343
rect 1825 -415 1871 -377
rect 1825 -449 1831 -415
rect 1865 -449 1871 -415
rect 1825 -487 1871 -449
rect 1825 -521 1831 -487
rect 1865 -521 1871 -487
rect 1825 -559 1871 -521
rect 1825 -593 1831 -559
rect 1865 -593 1871 -559
rect 1825 -631 1871 -593
rect 1825 -665 1831 -631
rect 1865 -665 1871 -631
rect 1825 -703 1871 -665
rect 1825 -737 1831 -703
rect 1865 -737 1871 -703
rect 1825 -775 1871 -737
rect 1825 -809 1831 -775
rect 1865 -809 1871 -775
rect 1825 -847 1871 -809
rect 1825 -881 1831 -847
rect 1865 -881 1871 -847
rect 1825 -904 1871 -881
rect 2133 953 2179 976
rect 2133 919 2139 953
rect 2173 919 2179 953
rect 2133 881 2179 919
rect 2133 847 2139 881
rect 2173 847 2179 881
rect 2133 809 2179 847
rect 2133 775 2139 809
rect 2173 775 2179 809
rect 2133 737 2179 775
rect 2133 703 2139 737
rect 2173 703 2179 737
rect 2133 665 2179 703
rect 2133 631 2139 665
rect 2173 631 2179 665
rect 2133 593 2179 631
rect 2133 559 2139 593
rect 2173 559 2179 593
rect 2133 521 2179 559
rect 2133 487 2139 521
rect 2173 487 2179 521
rect 2133 449 2179 487
rect 2133 415 2139 449
rect 2173 415 2179 449
rect 2133 377 2179 415
rect 2133 343 2139 377
rect 2173 343 2179 377
rect 2133 305 2179 343
rect 2133 271 2139 305
rect 2173 271 2179 305
rect 2133 233 2179 271
rect 2133 199 2139 233
rect 2173 199 2179 233
rect 2133 161 2179 199
rect 2133 127 2139 161
rect 2173 127 2179 161
rect 2133 89 2179 127
rect 2133 55 2139 89
rect 2173 55 2179 89
rect 2133 17 2179 55
rect 2133 -17 2139 17
rect 2173 -17 2179 17
rect 2133 -55 2179 -17
rect 2133 -89 2139 -55
rect 2173 -89 2179 -55
rect 2133 -127 2179 -89
rect 2133 -161 2139 -127
rect 2173 -161 2179 -127
rect 2133 -199 2179 -161
rect 2133 -233 2139 -199
rect 2173 -233 2179 -199
rect 2133 -271 2179 -233
rect 2133 -305 2139 -271
rect 2173 -305 2179 -271
rect 2133 -343 2179 -305
rect 2133 -377 2139 -343
rect 2173 -377 2179 -343
rect 2133 -415 2179 -377
rect 2133 -449 2139 -415
rect 2173 -449 2179 -415
rect 2133 -487 2179 -449
rect 2133 -521 2139 -487
rect 2173 -521 2179 -487
rect 2133 -559 2179 -521
rect 2133 -593 2139 -559
rect 2173 -593 2179 -559
rect 2133 -631 2179 -593
rect 2133 -665 2139 -631
rect 2173 -665 2179 -631
rect 2133 -703 2179 -665
rect 2133 -737 2139 -703
rect 2173 -737 2179 -703
rect 2133 -775 2179 -737
rect 2133 -809 2139 -775
rect 2173 -809 2179 -775
rect 2133 -847 2179 -809
rect 2133 -881 2139 -847
rect 2173 -881 2179 -847
rect 2133 -904 2179 -881
rect 2441 953 2487 976
rect 2441 919 2447 953
rect 2481 919 2487 953
rect 2441 881 2487 919
rect 2441 847 2447 881
rect 2481 847 2487 881
rect 2441 809 2487 847
rect 2441 775 2447 809
rect 2481 775 2487 809
rect 2441 737 2487 775
rect 2441 703 2447 737
rect 2481 703 2487 737
rect 2441 665 2487 703
rect 2441 631 2447 665
rect 2481 631 2487 665
rect 2441 593 2487 631
rect 2441 559 2447 593
rect 2481 559 2487 593
rect 2441 521 2487 559
rect 2441 487 2447 521
rect 2481 487 2487 521
rect 2441 449 2487 487
rect 2441 415 2447 449
rect 2481 415 2487 449
rect 2441 377 2487 415
rect 2441 343 2447 377
rect 2481 343 2487 377
rect 2441 305 2487 343
rect 2441 271 2447 305
rect 2481 271 2487 305
rect 2441 233 2487 271
rect 2441 199 2447 233
rect 2481 199 2487 233
rect 2441 161 2487 199
rect 2441 127 2447 161
rect 2481 127 2487 161
rect 2441 89 2487 127
rect 2441 55 2447 89
rect 2481 55 2487 89
rect 2441 17 2487 55
rect 2441 -17 2447 17
rect 2481 -17 2487 17
rect 2441 -55 2487 -17
rect 2441 -89 2447 -55
rect 2481 -89 2487 -55
rect 2441 -127 2487 -89
rect 2441 -161 2447 -127
rect 2481 -161 2487 -127
rect 2441 -199 2487 -161
rect 2441 -233 2447 -199
rect 2481 -233 2487 -199
rect 2441 -271 2487 -233
rect 2441 -305 2447 -271
rect 2481 -305 2487 -271
rect 2441 -343 2487 -305
rect 2441 -377 2447 -343
rect 2481 -377 2487 -343
rect 2441 -415 2487 -377
rect 2441 -449 2447 -415
rect 2481 -449 2487 -415
rect 2441 -487 2487 -449
rect 2441 -521 2447 -487
rect 2481 -521 2487 -487
rect 2441 -559 2487 -521
rect 2441 -593 2447 -559
rect 2481 -593 2487 -559
rect 2441 -631 2487 -593
rect 2441 -665 2447 -631
rect 2481 -665 2487 -631
rect 2441 -703 2487 -665
rect 2441 -737 2447 -703
rect 2481 -737 2487 -703
rect 2441 -775 2487 -737
rect 2441 -809 2447 -775
rect 2481 -809 2487 -775
rect 2441 -847 2487 -809
rect 2441 -881 2447 -847
rect 2481 -881 2487 -847
rect 2441 -904 2487 -881
rect 2749 953 2795 976
rect 2749 919 2755 953
rect 2789 919 2795 953
rect 2749 881 2795 919
rect 2749 847 2755 881
rect 2789 847 2795 881
rect 2749 809 2795 847
rect 2749 775 2755 809
rect 2789 775 2795 809
rect 2749 737 2795 775
rect 2749 703 2755 737
rect 2789 703 2795 737
rect 2749 665 2795 703
rect 2749 631 2755 665
rect 2789 631 2795 665
rect 2749 593 2795 631
rect 2749 559 2755 593
rect 2789 559 2795 593
rect 2749 521 2795 559
rect 2749 487 2755 521
rect 2789 487 2795 521
rect 2749 449 2795 487
rect 2749 415 2755 449
rect 2789 415 2795 449
rect 2749 377 2795 415
rect 2749 343 2755 377
rect 2789 343 2795 377
rect 2749 305 2795 343
rect 2749 271 2755 305
rect 2789 271 2795 305
rect 2749 233 2795 271
rect 2749 199 2755 233
rect 2789 199 2795 233
rect 2749 161 2795 199
rect 2749 127 2755 161
rect 2789 127 2795 161
rect 2749 89 2795 127
rect 2749 55 2755 89
rect 2789 55 2795 89
rect 2749 17 2795 55
rect 2749 -17 2755 17
rect 2789 -17 2795 17
rect 2749 -55 2795 -17
rect 2749 -89 2755 -55
rect 2789 -89 2795 -55
rect 2749 -127 2795 -89
rect 2749 -161 2755 -127
rect 2789 -161 2795 -127
rect 2749 -199 2795 -161
rect 2749 -233 2755 -199
rect 2789 -233 2795 -199
rect 2749 -271 2795 -233
rect 2749 -305 2755 -271
rect 2789 -305 2795 -271
rect 2749 -343 2795 -305
rect 2749 -377 2755 -343
rect 2789 -377 2795 -343
rect 2749 -415 2795 -377
rect 2749 -449 2755 -415
rect 2789 -449 2795 -415
rect 2749 -487 2795 -449
rect 2749 -521 2755 -487
rect 2789 -521 2795 -487
rect 2749 -559 2795 -521
rect 2749 -593 2755 -559
rect 2789 -593 2795 -559
rect 2749 -631 2795 -593
rect 2749 -665 2755 -631
rect 2789 -665 2795 -631
rect 2749 -703 2795 -665
rect 2749 -737 2755 -703
rect 2789 -737 2795 -703
rect 2749 -775 2795 -737
rect 2749 -809 2755 -775
rect 2789 -809 2795 -775
rect 2749 -847 2795 -809
rect 2749 -881 2755 -847
rect 2789 -881 2795 -847
rect 2749 -904 2795 -881
rect -2701 -951 -2535 -945
rect -2701 -985 -2671 -951
rect -2637 -985 -2599 -951
rect -2565 -985 -2535 -951
rect -2701 -991 -2535 -985
rect -2393 -951 -2227 -945
rect -2393 -985 -2363 -951
rect -2329 -985 -2291 -951
rect -2257 -985 -2227 -951
rect -2393 -991 -2227 -985
rect -2085 -951 -1919 -945
rect -2085 -985 -2055 -951
rect -2021 -985 -1983 -951
rect -1949 -985 -1919 -951
rect -2085 -991 -1919 -985
rect -1777 -951 -1611 -945
rect -1777 -985 -1747 -951
rect -1713 -985 -1675 -951
rect -1641 -985 -1611 -951
rect -1777 -991 -1611 -985
rect -1469 -951 -1303 -945
rect -1469 -985 -1439 -951
rect -1405 -985 -1367 -951
rect -1333 -985 -1303 -951
rect -1469 -991 -1303 -985
rect -1161 -951 -995 -945
rect -1161 -985 -1131 -951
rect -1097 -985 -1059 -951
rect -1025 -985 -995 -951
rect -1161 -991 -995 -985
rect -853 -951 -687 -945
rect -853 -985 -823 -951
rect -789 -985 -751 -951
rect -717 -985 -687 -951
rect -853 -991 -687 -985
rect -545 -951 -379 -945
rect -545 -985 -515 -951
rect -481 -985 -443 -951
rect -409 -985 -379 -951
rect -545 -991 -379 -985
rect -237 -951 -71 -945
rect -237 -985 -207 -951
rect -173 -985 -135 -951
rect -101 -985 -71 -951
rect -237 -991 -71 -985
rect 71 -951 237 -945
rect 71 -985 101 -951
rect 135 -985 173 -951
rect 207 -985 237 -951
rect 71 -991 237 -985
rect 379 -951 545 -945
rect 379 -985 409 -951
rect 443 -985 481 -951
rect 515 -985 545 -951
rect 379 -991 545 -985
rect 687 -951 853 -945
rect 687 -985 717 -951
rect 751 -985 789 -951
rect 823 -985 853 -951
rect 687 -991 853 -985
rect 995 -951 1161 -945
rect 995 -985 1025 -951
rect 1059 -985 1097 -951
rect 1131 -985 1161 -951
rect 995 -991 1161 -985
rect 1303 -951 1469 -945
rect 1303 -985 1333 -951
rect 1367 -985 1405 -951
rect 1439 -985 1469 -951
rect 1303 -991 1469 -985
rect 1611 -951 1777 -945
rect 1611 -985 1641 -951
rect 1675 -985 1713 -951
rect 1747 -985 1777 -951
rect 1611 -991 1777 -985
rect 1919 -951 2085 -945
rect 1919 -985 1949 -951
rect 1983 -985 2021 -951
rect 2055 -985 2085 -951
rect 1919 -991 2085 -985
rect 2227 -951 2393 -945
rect 2227 -985 2257 -951
rect 2291 -985 2329 -951
rect 2363 -985 2393 -951
rect 2227 -991 2393 -985
rect 2535 -951 2701 -945
rect 2535 -985 2565 -951
rect 2599 -985 2637 -951
rect 2671 -985 2701 -951
rect 2535 -991 2701 -985
<< end >>
