magic
tech sky130A
magscale 1 2
timestamp 1770083657
<< nwell >>
rect 1200 2100 9200 5200
rect 1200 -4200 1800 2100
rect 8600 -4200 9200 2100
rect 1200 -4600 9200 -4200
<< pwell >>
rect 2374 -2226 2526 -1774
rect 7874 -2226 8026 -1774
<< psubdiff >>
rect 2400 -2200 2500 -1800
rect 7900 -2200 8000 -1800
<< mvnsubdiff >>
rect 1300 5051 9100 5100
rect 1300 4949 1525 5051
rect 2035 4949 8365 5051
rect 8875 4949 9100 5051
rect 1300 4900 9100 4949
rect 1300 4873 1500 4900
rect 1300 -4273 1349 4873
rect 1451 -4273 1500 4873
rect 2080 4760 8280 4900
rect 8900 4873 9100 4900
rect 1300 -4300 1500 -4273
rect 8900 -4273 8949 4873
rect 9051 -4273 9100 4873
rect 8900 -4300 9100 -4273
rect 1300 -4349 9100 -4300
rect 1300 -4451 1545 -4349
rect 8855 -4451 9100 -4349
rect 1300 -4500 9100 -4451
<< mvnsubdiffcont >>
rect 1525 4949 2035 5051
rect 8365 4949 8875 5051
rect 1349 -4273 1451 4873
rect 8949 -4273 9051 4873
rect 1545 -4451 8855 -4349
<< locali >>
rect 1300 5051 9100 5100
rect 1300 4949 1525 5051
rect 2035 5047 8365 5051
rect 2035 5013 2113 5047
rect 2147 5013 2213 5047
rect 2247 5013 2313 5047
rect 2347 5013 2413 5047
rect 2447 5013 2513 5047
rect 2547 5013 2613 5047
rect 2647 5013 2713 5047
rect 2747 5013 2813 5047
rect 2847 5013 2913 5047
rect 2947 5013 3013 5047
rect 3047 5013 3113 5047
rect 3147 5013 3213 5047
rect 3247 5013 3313 5047
rect 3347 5013 3413 5047
rect 3447 5013 3513 5047
rect 3547 5013 3613 5047
rect 3647 5013 3713 5047
rect 3747 5013 3813 5047
rect 3847 5013 3913 5047
rect 3947 5013 4013 5047
rect 4047 5013 4113 5047
rect 4147 5013 4213 5047
rect 4247 5013 4313 5047
rect 4347 5013 4413 5047
rect 4447 5013 4513 5047
rect 4547 5013 4613 5047
rect 4647 5013 4713 5047
rect 4747 5013 4813 5047
rect 4847 5013 4913 5047
rect 4947 5013 5013 5047
rect 5047 5013 5113 5047
rect 5147 5013 5213 5047
rect 5247 5013 5313 5047
rect 5347 5013 5413 5047
rect 5447 5013 5513 5047
rect 5547 5013 5613 5047
rect 5647 5013 5713 5047
rect 5747 5013 5813 5047
rect 5847 5013 5913 5047
rect 5947 5013 6013 5047
rect 6047 5013 6113 5047
rect 6147 5013 6213 5047
rect 6247 5013 6313 5047
rect 6347 5013 6413 5047
rect 6447 5013 6513 5047
rect 6547 5013 6613 5047
rect 6647 5013 6713 5047
rect 6747 5013 6813 5047
rect 6847 5013 6913 5047
rect 6947 5013 7013 5047
rect 7047 5013 7113 5047
rect 7147 5013 7213 5047
rect 7247 5013 7313 5047
rect 7347 5013 7413 5047
rect 7447 5013 7513 5047
rect 7547 5013 7613 5047
rect 7647 5013 7713 5047
rect 7747 5013 7813 5047
rect 7847 5013 7913 5047
rect 7947 5013 8013 5047
rect 8047 5013 8113 5047
rect 8147 5013 8213 5047
rect 8247 5013 8365 5047
rect 2035 4949 8365 5013
rect 8875 4949 9100 5051
rect 1300 4947 9100 4949
rect 1300 4913 2113 4947
rect 2147 4913 2213 4947
rect 2247 4913 2313 4947
rect 2347 4913 2413 4947
rect 2447 4913 2513 4947
rect 2547 4913 2613 4947
rect 2647 4913 2713 4947
rect 2747 4913 2813 4947
rect 2847 4913 2913 4947
rect 2947 4913 3013 4947
rect 3047 4913 3113 4947
rect 3147 4913 3213 4947
rect 3247 4913 3313 4947
rect 3347 4913 3413 4947
rect 3447 4913 3513 4947
rect 3547 4913 3613 4947
rect 3647 4913 3713 4947
rect 3747 4913 3813 4947
rect 3847 4913 3913 4947
rect 3947 4913 4013 4947
rect 4047 4913 4113 4947
rect 4147 4913 4213 4947
rect 4247 4913 4313 4947
rect 4347 4913 4413 4947
rect 4447 4913 4513 4947
rect 4547 4913 4613 4947
rect 4647 4913 4713 4947
rect 4747 4913 4813 4947
rect 4847 4913 4913 4947
rect 4947 4913 5013 4947
rect 5047 4913 5113 4947
rect 5147 4913 5213 4947
rect 5247 4913 5313 4947
rect 5347 4913 5413 4947
rect 5447 4913 5513 4947
rect 5547 4913 5613 4947
rect 5647 4913 5713 4947
rect 5747 4913 5813 4947
rect 5847 4913 5913 4947
rect 5947 4913 6013 4947
rect 6047 4913 6113 4947
rect 6147 4913 6213 4947
rect 6247 4913 6313 4947
rect 6347 4913 6413 4947
rect 6447 4913 6513 4947
rect 6547 4913 6613 4947
rect 6647 4913 6713 4947
rect 6747 4913 6813 4947
rect 6847 4913 6913 4947
rect 6947 4913 7013 4947
rect 7047 4913 7113 4947
rect 7147 4913 7213 4947
rect 7247 4913 7313 4947
rect 7347 4913 7413 4947
rect 7447 4913 7513 4947
rect 7547 4913 7613 4947
rect 7647 4913 7713 4947
rect 7747 4913 7813 4947
rect 7847 4913 7913 4947
rect 7947 4913 8013 4947
rect 8047 4913 8113 4947
rect 8147 4913 8213 4947
rect 8247 4913 9100 4947
rect 1300 4873 9100 4913
rect 1300 -4273 1349 4873
rect 1451 4847 8949 4873
rect 1451 4813 2113 4847
rect 2147 4813 2213 4847
rect 2247 4813 2313 4847
rect 2347 4813 2413 4847
rect 2447 4813 2513 4847
rect 2547 4813 2613 4847
rect 2647 4813 2713 4847
rect 2747 4813 2813 4847
rect 2847 4813 2913 4847
rect 2947 4813 3013 4847
rect 3047 4813 3113 4847
rect 3147 4813 3213 4847
rect 3247 4813 3313 4847
rect 3347 4813 3413 4847
rect 3447 4813 3513 4847
rect 3547 4813 3613 4847
rect 3647 4813 3713 4847
rect 3747 4813 3813 4847
rect 3847 4813 3913 4847
rect 3947 4813 4013 4847
rect 4047 4813 4113 4847
rect 4147 4813 4213 4847
rect 4247 4813 4313 4847
rect 4347 4813 4413 4847
rect 4447 4813 4513 4847
rect 4547 4813 4613 4847
rect 4647 4813 4713 4847
rect 4747 4813 4813 4847
rect 4847 4813 4913 4847
rect 4947 4813 5013 4847
rect 5047 4813 5113 4847
rect 5147 4813 5213 4847
rect 5247 4813 5313 4847
rect 5347 4813 5413 4847
rect 5447 4813 5513 4847
rect 5547 4813 5613 4847
rect 5647 4813 5713 4847
rect 5747 4813 5813 4847
rect 5847 4813 5913 4847
rect 5947 4813 6013 4847
rect 6047 4813 6113 4847
rect 6147 4813 6213 4847
rect 6247 4813 6313 4847
rect 6347 4813 6413 4847
rect 6447 4813 6513 4847
rect 6547 4813 6613 4847
rect 6647 4813 6713 4847
rect 6747 4813 6813 4847
rect 6847 4813 6913 4847
rect 6947 4813 7013 4847
rect 7047 4813 7113 4847
rect 7147 4813 7213 4847
rect 7247 4813 7313 4847
rect 7347 4813 7413 4847
rect 7447 4813 7513 4847
rect 7547 4813 7613 4847
rect 7647 4813 7713 4847
rect 7747 4813 7813 4847
rect 7847 4813 7913 4847
rect 7947 4813 8013 4847
rect 8047 4813 8113 4847
rect 8147 4813 8213 4847
rect 8247 4813 8949 4847
rect 1451 4760 8949 4813
rect 1451 2496 2176 4760
rect 8216 2500 8949 4760
rect 4760 2496 8949 2500
rect 1451 2100 8949 2496
rect 1451 2098 4800 2100
rect 1451 -4273 1500 2098
rect 1560 -1800 2400 2000
rect 8000 -1800 8840 2000
rect 1560 -1883 4920 -1800
rect 1560 -1917 2563 -1883
rect 2597 -1917 2683 -1883
rect 2717 -1917 2803 -1883
rect 2837 -1917 2923 -1883
rect 2957 -1917 3043 -1883
rect 3077 -1917 3163 -1883
rect 3197 -1917 3283 -1883
rect 3317 -1917 3403 -1883
rect 3437 -1917 3523 -1883
rect 3557 -1917 3643 -1883
rect 3677 -1917 3763 -1883
rect 3797 -1917 3883 -1883
rect 3917 -1917 4003 -1883
rect 4037 -1917 4123 -1883
rect 4157 -1917 4243 -1883
rect 4277 -1917 4363 -1883
rect 4397 -1917 4483 -1883
rect 4517 -1917 4603 -1883
rect 4637 -1917 4723 -1883
rect 4757 -1917 4843 -1883
rect 4877 -1917 4920 -1883
rect 1560 -2003 4920 -1917
rect 1560 -2037 2443 -2003
rect 2477 -2037 2563 -2003
rect 2597 -2037 2683 -2003
rect 2717 -2037 2803 -2003
rect 2837 -2037 2923 -2003
rect 2957 -2037 3043 -2003
rect 3077 -2037 3163 -2003
rect 3197 -2037 3283 -2003
rect 3317 -2037 3403 -2003
rect 3437 -2037 3523 -2003
rect 3557 -2037 3643 -2003
rect 3677 -2037 3763 -2003
rect 3797 -2037 3883 -2003
rect 3917 -2037 4003 -2003
rect 4037 -2037 4123 -2003
rect 4157 -2037 4243 -2003
rect 4277 -2037 4363 -2003
rect 4397 -2037 4483 -2003
rect 4517 -2037 4603 -2003
rect 4637 -2037 4723 -2003
rect 4757 -2037 4843 -2003
rect 4877 -2037 4920 -2003
rect 1560 -2123 4920 -2037
rect 1560 -2140 2443 -2123
rect 1560 -4100 2225 -2140
rect 2400 -2157 2443 -2140
rect 2477 -2157 2563 -2123
rect 2597 -2157 2683 -2123
rect 2717 -2157 2803 -2123
rect 2837 -2157 2923 -2123
rect 2957 -2157 3043 -2123
rect 3077 -2157 3163 -2123
rect 3197 -2157 3283 -2123
rect 3317 -2157 3403 -2123
rect 3437 -2157 3523 -2123
rect 3557 -2157 3643 -2123
rect 3677 -2157 3763 -2123
rect 3797 -2157 3883 -2123
rect 3917 -2157 4003 -2123
rect 4037 -2157 4123 -2123
rect 4157 -2157 4243 -2123
rect 4277 -2157 4363 -2123
rect 4397 -2157 4483 -2123
rect 4517 -2157 4603 -2123
rect 4637 -2157 4723 -2123
rect 4757 -2157 4843 -2123
rect 4877 -2157 4920 -2123
rect 2400 -2200 4920 -2157
rect 5480 -1883 8840 -1800
rect 5480 -1917 5523 -1883
rect 5557 -1917 5643 -1883
rect 5677 -1917 5763 -1883
rect 5797 -1917 5883 -1883
rect 5917 -1917 6003 -1883
rect 6037 -1917 6123 -1883
rect 6157 -1917 6243 -1883
rect 6277 -1917 6363 -1883
rect 6397 -1917 6483 -1883
rect 6517 -1917 6603 -1883
rect 6637 -1917 6723 -1883
rect 6757 -1917 6843 -1883
rect 6877 -1917 6963 -1883
rect 6997 -1917 7083 -1883
rect 7117 -1917 7203 -1883
rect 7237 -1917 7323 -1883
rect 7357 -1917 7443 -1883
rect 7477 -1917 7563 -1883
rect 7597 -1917 7683 -1883
rect 7717 -1917 7803 -1883
rect 7837 -1917 7923 -1883
rect 7957 -1917 8840 -1883
rect 5480 -2003 8840 -1917
rect 5480 -2037 5523 -2003
rect 5557 -2037 5643 -2003
rect 5677 -2037 5763 -2003
rect 5797 -2037 5883 -2003
rect 5917 -2037 6003 -2003
rect 6037 -2037 6123 -2003
rect 6157 -2037 6243 -2003
rect 6277 -2037 6363 -2003
rect 6397 -2037 6483 -2003
rect 6517 -2037 6603 -2003
rect 6637 -2037 6723 -2003
rect 6757 -2037 6843 -2003
rect 6877 -2037 6963 -2003
rect 6997 -2037 7083 -2003
rect 7117 -2037 7203 -2003
rect 7237 -2037 7323 -2003
rect 7357 -2037 7443 -2003
rect 7477 -2037 7563 -2003
rect 7597 -2037 7683 -2003
rect 7717 -2037 7803 -2003
rect 7837 -2037 7923 -2003
rect 7957 -2037 8840 -2003
rect 5480 -2123 8840 -2037
rect 5480 -2157 5523 -2123
rect 5557 -2157 5643 -2123
rect 5677 -2157 5763 -2123
rect 5797 -2157 5883 -2123
rect 5917 -2157 6003 -2123
rect 6037 -2157 6123 -2123
rect 6157 -2157 6243 -2123
rect 6277 -2157 6363 -2123
rect 6397 -2157 6483 -2123
rect 6517 -2157 6603 -2123
rect 6637 -2157 6723 -2123
rect 6757 -2157 6843 -2123
rect 6877 -2157 6963 -2123
rect 6997 -2157 7083 -2123
rect 7117 -2157 7203 -2123
rect 7237 -2157 7323 -2123
rect 7357 -2157 7443 -2123
rect 7477 -2157 7563 -2123
rect 7597 -2157 7683 -2123
rect 7717 -2157 7803 -2123
rect 7837 -2157 7923 -2123
rect 7957 -2157 8840 -2123
rect 5480 -2160 8840 -2157
rect 5480 -2200 8000 -2160
rect 8200 -4100 8840 -2160
rect 1560 -4260 8840 -4100
rect 1300 -4300 1500 -4273
rect 8900 -4273 8949 2100
rect 9051 -4273 9100 4873
rect 8900 -4300 9100 -4273
rect 1300 -4349 9100 -4300
rect 1300 -4451 1545 -4349
rect 8855 -4451 9100 -4349
rect 1300 -4500 9100 -4451
<< viali >>
rect 2113 5013 2147 5047
rect 2213 5013 2247 5047
rect 2313 5013 2347 5047
rect 2413 5013 2447 5047
rect 2513 5013 2547 5047
rect 2613 5013 2647 5047
rect 2713 5013 2747 5047
rect 2813 5013 2847 5047
rect 2913 5013 2947 5047
rect 3013 5013 3047 5047
rect 3113 5013 3147 5047
rect 3213 5013 3247 5047
rect 3313 5013 3347 5047
rect 3413 5013 3447 5047
rect 3513 5013 3547 5047
rect 3613 5013 3647 5047
rect 3713 5013 3747 5047
rect 3813 5013 3847 5047
rect 3913 5013 3947 5047
rect 4013 5013 4047 5047
rect 4113 5013 4147 5047
rect 4213 5013 4247 5047
rect 4313 5013 4347 5047
rect 4413 5013 4447 5047
rect 4513 5013 4547 5047
rect 4613 5013 4647 5047
rect 4713 5013 4747 5047
rect 4813 5013 4847 5047
rect 4913 5013 4947 5047
rect 5013 5013 5047 5047
rect 5113 5013 5147 5047
rect 5213 5013 5247 5047
rect 5313 5013 5347 5047
rect 5413 5013 5447 5047
rect 5513 5013 5547 5047
rect 5613 5013 5647 5047
rect 5713 5013 5747 5047
rect 5813 5013 5847 5047
rect 5913 5013 5947 5047
rect 6013 5013 6047 5047
rect 6113 5013 6147 5047
rect 6213 5013 6247 5047
rect 6313 5013 6347 5047
rect 6413 5013 6447 5047
rect 6513 5013 6547 5047
rect 6613 5013 6647 5047
rect 6713 5013 6747 5047
rect 6813 5013 6847 5047
rect 6913 5013 6947 5047
rect 7013 5013 7047 5047
rect 7113 5013 7147 5047
rect 7213 5013 7247 5047
rect 7313 5013 7347 5047
rect 7413 5013 7447 5047
rect 7513 5013 7547 5047
rect 7613 5013 7647 5047
rect 7713 5013 7747 5047
rect 7813 5013 7847 5047
rect 7913 5013 7947 5047
rect 8013 5013 8047 5047
rect 8113 5013 8147 5047
rect 8213 5013 8247 5047
rect 2113 4913 2147 4947
rect 2213 4913 2247 4947
rect 2313 4913 2347 4947
rect 2413 4913 2447 4947
rect 2513 4913 2547 4947
rect 2613 4913 2647 4947
rect 2713 4913 2747 4947
rect 2813 4913 2847 4947
rect 2913 4913 2947 4947
rect 3013 4913 3047 4947
rect 3113 4913 3147 4947
rect 3213 4913 3247 4947
rect 3313 4913 3347 4947
rect 3413 4913 3447 4947
rect 3513 4913 3547 4947
rect 3613 4913 3647 4947
rect 3713 4913 3747 4947
rect 3813 4913 3847 4947
rect 3913 4913 3947 4947
rect 4013 4913 4047 4947
rect 4113 4913 4147 4947
rect 4213 4913 4247 4947
rect 4313 4913 4347 4947
rect 4413 4913 4447 4947
rect 4513 4913 4547 4947
rect 4613 4913 4647 4947
rect 4713 4913 4747 4947
rect 4813 4913 4847 4947
rect 4913 4913 4947 4947
rect 5013 4913 5047 4947
rect 5113 4913 5147 4947
rect 5213 4913 5247 4947
rect 5313 4913 5347 4947
rect 5413 4913 5447 4947
rect 5513 4913 5547 4947
rect 5613 4913 5647 4947
rect 5713 4913 5747 4947
rect 5813 4913 5847 4947
rect 5913 4913 5947 4947
rect 6013 4913 6047 4947
rect 6113 4913 6147 4947
rect 6213 4913 6247 4947
rect 6313 4913 6347 4947
rect 6413 4913 6447 4947
rect 6513 4913 6547 4947
rect 6613 4913 6647 4947
rect 6713 4913 6747 4947
rect 6813 4913 6847 4947
rect 6913 4913 6947 4947
rect 7013 4913 7047 4947
rect 7113 4913 7147 4947
rect 7213 4913 7247 4947
rect 7313 4913 7347 4947
rect 7413 4913 7447 4947
rect 7513 4913 7547 4947
rect 7613 4913 7647 4947
rect 7713 4913 7747 4947
rect 7813 4913 7847 4947
rect 7913 4913 7947 4947
rect 8013 4913 8047 4947
rect 8113 4913 8147 4947
rect 8213 4913 8247 4947
rect 2113 4813 2147 4847
rect 2213 4813 2247 4847
rect 2313 4813 2347 4847
rect 2413 4813 2447 4847
rect 2513 4813 2547 4847
rect 2613 4813 2647 4847
rect 2713 4813 2747 4847
rect 2813 4813 2847 4847
rect 2913 4813 2947 4847
rect 3013 4813 3047 4847
rect 3113 4813 3147 4847
rect 3213 4813 3247 4847
rect 3313 4813 3347 4847
rect 3413 4813 3447 4847
rect 3513 4813 3547 4847
rect 3613 4813 3647 4847
rect 3713 4813 3747 4847
rect 3813 4813 3847 4847
rect 3913 4813 3947 4847
rect 4013 4813 4047 4847
rect 4113 4813 4147 4847
rect 4213 4813 4247 4847
rect 4313 4813 4347 4847
rect 4413 4813 4447 4847
rect 4513 4813 4547 4847
rect 4613 4813 4647 4847
rect 4713 4813 4747 4847
rect 4813 4813 4847 4847
rect 4913 4813 4947 4847
rect 5013 4813 5047 4847
rect 5113 4813 5147 4847
rect 5213 4813 5247 4847
rect 5313 4813 5347 4847
rect 5413 4813 5447 4847
rect 5513 4813 5547 4847
rect 5613 4813 5647 4847
rect 5713 4813 5747 4847
rect 5813 4813 5847 4847
rect 5913 4813 5947 4847
rect 6013 4813 6047 4847
rect 6113 4813 6147 4847
rect 6213 4813 6247 4847
rect 6313 4813 6347 4847
rect 6413 4813 6447 4847
rect 6513 4813 6547 4847
rect 6613 4813 6647 4847
rect 6713 4813 6747 4847
rect 6813 4813 6847 4847
rect 6913 4813 6947 4847
rect 7013 4813 7047 4847
rect 7113 4813 7147 4847
rect 7213 4813 7247 4847
rect 7313 4813 7347 4847
rect 7413 4813 7447 4847
rect 7513 4813 7547 4847
rect 7613 4813 7647 4847
rect 7713 4813 7747 4847
rect 7813 4813 7847 4847
rect 7913 4813 7947 4847
rect 8013 4813 8047 4847
rect 8113 4813 8147 4847
rect 8213 4813 8247 4847
rect 2563 -1917 2597 -1883
rect 2683 -1917 2717 -1883
rect 2803 -1917 2837 -1883
rect 2923 -1917 2957 -1883
rect 3043 -1917 3077 -1883
rect 3163 -1917 3197 -1883
rect 3283 -1917 3317 -1883
rect 3403 -1917 3437 -1883
rect 3523 -1917 3557 -1883
rect 3643 -1917 3677 -1883
rect 3763 -1917 3797 -1883
rect 3883 -1917 3917 -1883
rect 4003 -1917 4037 -1883
rect 4123 -1917 4157 -1883
rect 4243 -1917 4277 -1883
rect 4363 -1917 4397 -1883
rect 4483 -1917 4517 -1883
rect 4603 -1917 4637 -1883
rect 4723 -1917 4757 -1883
rect 4843 -1917 4877 -1883
rect 2443 -2037 2477 -2003
rect 2563 -2037 2597 -2003
rect 2683 -2037 2717 -2003
rect 2803 -2037 2837 -2003
rect 2923 -2037 2957 -2003
rect 3043 -2037 3077 -2003
rect 3163 -2037 3197 -2003
rect 3283 -2037 3317 -2003
rect 3403 -2037 3437 -2003
rect 3523 -2037 3557 -2003
rect 3643 -2037 3677 -2003
rect 3763 -2037 3797 -2003
rect 3883 -2037 3917 -2003
rect 4003 -2037 4037 -2003
rect 4123 -2037 4157 -2003
rect 4243 -2037 4277 -2003
rect 4363 -2037 4397 -2003
rect 4483 -2037 4517 -2003
rect 4603 -2037 4637 -2003
rect 4723 -2037 4757 -2003
rect 4843 -2037 4877 -2003
rect 2443 -2157 2477 -2123
rect 2563 -2157 2597 -2123
rect 2683 -2157 2717 -2123
rect 2803 -2157 2837 -2123
rect 2923 -2157 2957 -2123
rect 3043 -2157 3077 -2123
rect 3163 -2157 3197 -2123
rect 3283 -2157 3317 -2123
rect 3403 -2157 3437 -2123
rect 3523 -2157 3557 -2123
rect 3643 -2157 3677 -2123
rect 3763 -2157 3797 -2123
rect 3883 -2157 3917 -2123
rect 4003 -2157 4037 -2123
rect 4123 -2157 4157 -2123
rect 4243 -2157 4277 -2123
rect 4363 -2157 4397 -2123
rect 4483 -2157 4517 -2123
rect 4603 -2157 4637 -2123
rect 4723 -2157 4757 -2123
rect 4843 -2157 4877 -2123
rect 5523 -1917 5557 -1883
rect 5643 -1917 5677 -1883
rect 5763 -1917 5797 -1883
rect 5883 -1917 5917 -1883
rect 6003 -1917 6037 -1883
rect 6123 -1917 6157 -1883
rect 6243 -1917 6277 -1883
rect 6363 -1917 6397 -1883
rect 6483 -1917 6517 -1883
rect 6603 -1917 6637 -1883
rect 6723 -1917 6757 -1883
rect 6843 -1917 6877 -1883
rect 6963 -1917 6997 -1883
rect 7083 -1917 7117 -1883
rect 7203 -1917 7237 -1883
rect 7323 -1917 7357 -1883
rect 7443 -1917 7477 -1883
rect 7563 -1917 7597 -1883
rect 7683 -1917 7717 -1883
rect 7803 -1917 7837 -1883
rect 7923 -1917 7957 -1883
rect 5523 -2037 5557 -2003
rect 5643 -2037 5677 -2003
rect 5763 -2037 5797 -2003
rect 5883 -2037 5917 -2003
rect 6003 -2037 6037 -2003
rect 6123 -2037 6157 -2003
rect 6243 -2037 6277 -2003
rect 6363 -2037 6397 -2003
rect 6483 -2037 6517 -2003
rect 6603 -2037 6637 -2003
rect 6723 -2037 6757 -2003
rect 6843 -2037 6877 -2003
rect 6963 -2037 6997 -2003
rect 7083 -2037 7117 -2003
rect 7203 -2037 7237 -2003
rect 7323 -2037 7357 -2003
rect 7443 -2037 7477 -2003
rect 7563 -2037 7597 -2003
rect 7683 -2037 7717 -2003
rect 7803 -2037 7837 -2003
rect 7923 -2037 7957 -2003
rect 5523 -2157 5557 -2123
rect 5643 -2157 5677 -2123
rect 5763 -2157 5797 -2123
rect 5883 -2157 5917 -2123
rect 6003 -2157 6037 -2123
rect 6123 -2157 6157 -2123
rect 6243 -2157 6277 -2123
rect 6363 -2157 6397 -2123
rect 6483 -2157 6517 -2123
rect 6603 -2157 6637 -2123
rect 6723 -2157 6757 -2123
rect 6843 -2157 6877 -2123
rect 6963 -2157 6997 -2123
rect 7083 -2157 7117 -2123
rect 7203 -2157 7237 -2123
rect 7323 -2157 7357 -2123
rect 7443 -2157 7477 -2123
rect 7563 -2157 7597 -2123
rect 7683 -2157 7717 -2123
rect 7803 -2157 7837 -2123
rect 7923 -2157 7957 -2123
<< metal1 >>
rect 2080 5047 8280 5100
rect 2080 5013 2113 5047
rect 2147 5013 2213 5047
rect 2247 5013 2313 5047
rect 2347 5013 2413 5047
rect 2447 5013 2513 5047
rect 2547 5013 2613 5047
rect 2647 5013 2713 5047
rect 2747 5013 2813 5047
rect 2847 5013 2913 5047
rect 2947 5013 3013 5047
rect 3047 5013 3113 5047
rect 3147 5013 3213 5047
rect 3247 5013 3313 5047
rect 3347 5013 3413 5047
rect 3447 5013 3513 5047
rect 3547 5013 3613 5047
rect 3647 5013 3713 5047
rect 3747 5013 3813 5047
rect 3847 5013 3913 5047
rect 3947 5013 4013 5047
rect 4047 5013 4113 5047
rect 4147 5013 4213 5047
rect 4247 5013 4313 5047
rect 4347 5013 4413 5047
rect 4447 5013 4513 5047
rect 4547 5013 4613 5047
rect 4647 5013 4713 5047
rect 4747 5013 4813 5047
rect 4847 5013 4913 5047
rect 4947 5013 5013 5047
rect 5047 5013 5113 5047
rect 5147 5013 5213 5047
rect 5247 5013 5313 5047
rect 5347 5013 5413 5047
rect 5447 5013 5513 5047
rect 5547 5013 5613 5047
rect 5647 5013 5713 5047
rect 5747 5013 5813 5047
rect 5847 5013 5913 5047
rect 5947 5013 6013 5047
rect 6047 5013 6113 5047
rect 6147 5013 6213 5047
rect 6247 5013 6313 5047
rect 6347 5013 6413 5047
rect 6447 5013 6513 5047
rect 6547 5013 6613 5047
rect 6647 5013 6713 5047
rect 6747 5013 6813 5047
rect 6847 5013 6913 5047
rect 6947 5013 7013 5047
rect 7047 5013 7113 5047
rect 7147 5013 7213 5047
rect 7247 5013 7313 5047
rect 7347 5013 7413 5047
rect 7447 5013 7513 5047
rect 7547 5013 7613 5047
rect 7647 5013 7713 5047
rect 7747 5013 7813 5047
rect 7847 5013 7913 5047
rect 7947 5013 8013 5047
rect 8047 5013 8113 5047
rect 8147 5013 8213 5047
rect 8247 5013 8280 5047
rect 2080 4947 8280 5013
rect 2080 4913 2113 4947
rect 2147 4913 2213 4947
rect 2247 4913 2313 4947
rect 2347 4913 2413 4947
rect 2447 4913 2513 4947
rect 2547 4913 2613 4947
rect 2647 4913 2713 4947
rect 2747 4913 2813 4947
rect 2847 4913 2913 4947
rect 2947 4913 3013 4947
rect 3047 4913 3113 4947
rect 3147 4913 3213 4947
rect 3247 4913 3313 4947
rect 3347 4913 3413 4947
rect 3447 4913 3513 4947
rect 3547 4913 3613 4947
rect 3647 4913 3713 4947
rect 3747 4913 3813 4947
rect 3847 4913 3913 4947
rect 3947 4913 4013 4947
rect 4047 4913 4113 4947
rect 4147 4913 4213 4947
rect 4247 4913 4313 4947
rect 4347 4913 4413 4947
rect 4447 4913 4513 4947
rect 4547 4913 4613 4947
rect 4647 4913 4713 4947
rect 4747 4913 4813 4947
rect 4847 4913 4913 4947
rect 4947 4913 5013 4947
rect 5047 4913 5113 4947
rect 5147 4913 5213 4947
rect 5247 4913 5313 4947
rect 5347 4913 5413 4947
rect 5447 4913 5513 4947
rect 5547 4913 5613 4947
rect 5647 4913 5713 4947
rect 5747 4913 5813 4947
rect 5847 4913 5913 4947
rect 5947 4913 6013 4947
rect 6047 4913 6113 4947
rect 6147 4913 6213 4947
rect 6247 4913 6313 4947
rect 6347 4913 6413 4947
rect 6447 4913 6513 4947
rect 6547 4913 6613 4947
rect 6647 4913 6713 4947
rect 6747 4913 6813 4947
rect 6847 4913 6913 4947
rect 6947 4913 7013 4947
rect 7047 4913 7113 4947
rect 7147 4913 7213 4947
rect 7247 4913 7313 4947
rect 7347 4913 7413 4947
rect 7447 4913 7513 4947
rect 7547 4913 7613 4947
rect 7647 4913 7713 4947
rect 7747 4913 7813 4947
rect 7847 4913 7913 4947
rect 7947 4913 8013 4947
rect 8047 4913 8113 4947
rect 8147 4913 8213 4947
rect 8247 4913 8280 4947
rect 2080 4847 8280 4913
rect 2080 4813 2113 4847
rect 2147 4813 2213 4847
rect 2247 4813 2313 4847
rect 2347 4813 2413 4847
rect 2447 4813 2513 4847
rect 2547 4813 2613 4847
rect 2647 4813 2713 4847
rect 2747 4813 2813 4847
rect 2847 4813 2913 4847
rect 2947 4813 3013 4847
rect 3047 4813 3113 4847
rect 3147 4813 3213 4847
rect 3247 4813 3313 4847
rect 3347 4813 3413 4847
rect 3447 4813 3513 4847
rect 3547 4813 3613 4847
rect 3647 4813 3713 4847
rect 3747 4813 3813 4847
rect 3847 4813 3913 4847
rect 3947 4813 4013 4847
rect 4047 4813 4113 4847
rect 4147 4813 4213 4847
rect 4247 4813 4313 4847
rect 4347 4813 4413 4847
rect 4447 4813 4513 4847
rect 4547 4813 4613 4847
rect 4647 4813 4713 4847
rect 4747 4813 4813 4847
rect 4847 4813 4913 4847
rect 4947 4813 5013 4847
rect 5047 4813 5113 4847
rect 5147 4813 5213 4847
rect 5247 4813 5313 4847
rect 5347 4813 5413 4847
rect 5447 4813 5513 4847
rect 5547 4813 5613 4847
rect 5647 4813 5713 4847
rect 5747 4813 5813 4847
rect 5847 4813 5913 4847
rect 5947 4813 6013 4847
rect 6047 4813 6113 4847
rect 6147 4813 6213 4847
rect 6247 4813 6313 4847
rect 6347 4813 6413 4847
rect 6447 4813 6513 4847
rect 6547 4813 6613 4847
rect 6647 4813 6713 4847
rect 6747 4813 6813 4847
rect 6847 4813 6913 4847
rect 6947 4813 7013 4847
rect 7047 4813 7113 4847
rect 7147 4813 7213 4847
rect 7247 4813 7313 4847
rect 7347 4813 7413 4847
rect 7447 4813 7513 4847
rect 7547 4813 7613 4847
rect 7647 4813 7713 4847
rect 7747 4813 7813 4847
rect 7847 4813 7913 4847
rect 7947 4813 8013 4847
rect 8047 4813 8113 4847
rect 8147 4813 8213 4847
rect 8247 4813 8280 4847
rect 2080 4760 8280 4813
rect 5000 2276 5400 2300
rect 5000 2224 5024 2276
rect 5076 2224 5104 2276
rect 5156 2224 5244 2276
rect 5296 2224 5324 2276
rect 5376 2224 5400 2276
rect 5000 2176 5400 2224
rect 5000 2124 5024 2176
rect 5076 2124 5104 2176
rect 5156 2124 5244 2176
rect 5296 2124 5324 2176
rect 5376 2124 5400 2176
rect 5000 2100 5400 2124
rect 2400 -1883 4920 -1800
rect 2400 -1917 2563 -1883
rect 2597 -1917 2683 -1883
rect 2717 -1917 2803 -1883
rect 2837 -1917 2923 -1883
rect 2957 -1917 3043 -1883
rect 3077 -1917 3163 -1883
rect 3197 -1917 3283 -1883
rect 3317 -1917 3403 -1883
rect 3437 -1917 3523 -1883
rect 3557 -1917 3643 -1883
rect 3677 -1917 3763 -1883
rect 3797 -1917 3883 -1883
rect 3917 -1917 4003 -1883
rect 4037 -1917 4123 -1883
rect 4157 -1917 4243 -1883
rect 4277 -1917 4363 -1883
rect 4397 -1917 4483 -1883
rect 4517 -1917 4603 -1883
rect 4637 -1917 4723 -1883
rect 4757 -1917 4843 -1883
rect 4877 -1917 4920 -1883
rect 2400 -2003 4920 -1917
rect 2400 -2037 2443 -2003
rect 2477 -2037 2563 -2003
rect 2597 -2037 2683 -2003
rect 2717 -2037 2803 -2003
rect 2837 -2037 2923 -2003
rect 2957 -2037 3043 -2003
rect 3077 -2037 3163 -2003
rect 3197 -2037 3283 -2003
rect 3317 -2037 3403 -2003
rect 3437 -2037 3523 -2003
rect 3557 -2037 3643 -2003
rect 3677 -2037 3763 -2003
rect 3797 -2037 3883 -2003
rect 3917 -2037 4003 -2003
rect 4037 -2037 4123 -2003
rect 4157 -2037 4243 -2003
rect 4277 -2037 4363 -2003
rect 4397 -2037 4483 -2003
rect 4517 -2037 4603 -2003
rect 4637 -2037 4723 -2003
rect 4757 -2037 4843 -2003
rect 4877 -2037 4920 -2003
rect 2400 -2123 4920 -2037
rect 2400 -2157 2443 -2123
rect 2477 -2157 2563 -2123
rect 2597 -2157 2683 -2123
rect 2717 -2157 2803 -2123
rect 2837 -2157 2923 -2123
rect 2957 -2157 3043 -2123
rect 3077 -2157 3163 -2123
rect 3197 -2157 3283 -2123
rect 3317 -2157 3403 -2123
rect 3437 -2157 3523 -2123
rect 3557 -2157 3643 -2123
rect 3677 -2157 3763 -2123
rect 3797 -2157 3883 -2123
rect 3917 -2157 4003 -2123
rect 4037 -2157 4123 -2123
rect 4157 -2157 4243 -2123
rect 4277 -2157 4363 -2123
rect 4397 -2157 4483 -2123
rect 4517 -2157 4603 -2123
rect 4637 -2157 4723 -2123
rect 4757 -2157 4843 -2123
rect 4877 -2157 4920 -2123
rect 2400 -2200 4920 -2157
rect 5480 -1883 8000 -1800
rect 5480 -1917 5523 -1883
rect 5557 -1917 5643 -1883
rect 5677 -1917 5763 -1883
rect 5797 -1917 5883 -1883
rect 5917 -1917 6003 -1883
rect 6037 -1917 6123 -1883
rect 6157 -1917 6243 -1883
rect 6277 -1917 6363 -1883
rect 6397 -1917 6483 -1883
rect 6517 -1917 6603 -1883
rect 6637 -1917 6723 -1883
rect 6757 -1917 6843 -1883
rect 6877 -1917 6963 -1883
rect 6997 -1917 7083 -1883
rect 7117 -1917 7203 -1883
rect 7237 -1917 7323 -1883
rect 7357 -1917 7443 -1883
rect 7477 -1917 7563 -1883
rect 7597 -1917 7683 -1883
rect 7717 -1917 7803 -1883
rect 7837 -1917 7923 -1883
rect 7957 -1917 8000 -1883
rect 5480 -2003 8000 -1917
rect 5480 -2037 5523 -2003
rect 5557 -2037 5643 -2003
rect 5677 -2037 5763 -2003
rect 5797 -2037 5883 -2003
rect 5917 -2037 6003 -2003
rect 6037 -2037 6123 -2003
rect 6157 -2037 6243 -2003
rect 6277 -2037 6363 -2003
rect 6397 -2037 6483 -2003
rect 6517 -2037 6603 -2003
rect 6637 -2037 6723 -2003
rect 6757 -2037 6843 -2003
rect 6877 -2037 6963 -2003
rect 6997 -2037 7083 -2003
rect 7117 -2037 7203 -2003
rect 7237 -2037 7323 -2003
rect 7357 -2037 7443 -2003
rect 7477 -2037 7563 -2003
rect 7597 -2037 7683 -2003
rect 7717 -2037 7803 -2003
rect 7837 -2037 7923 -2003
rect 7957 -2037 8000 -2003
rect 5480 -2123 8000 -2037
rect 5480 -2157 5523 -2123
rect 5557 -2157 5643 -2123
rect 5677 -2157 5763 -2123
rect 5797 -2157 5883 -2123
rect 5917 -2157 6003 -2123
rect 6037 -2157 6123 -2123
rect 6157 -2157 6243 -2123
rect 6277 -2157 6363 -2123
rect 6397 -2157 6483 -2123
rect 6517 -2157 6603 -2123
rect 6637 -2157 6723 -2123
rect 6757 -2157 6843 -2123
rect 6877 -2157 6963 -2123
rect 6997 -2157 7083 -2123
rect 7117 -2157 7203 -2123
rect 7237 -2157 7323 -2123
rect 7357 -2157 7443 -2123
rect 7477 -2157 7563 -2123
rect 7597 -2157 7683 -2123
rect 7717 -2157 7803 -2123
rect 7837 -2157 7923 -2123
rect 7957 -2157 8000 -2123
rect 5480 -2200 8000 -2157
<< via1 >>
rect 5024 2224 5076 2276
rect 5104 2224 5156 2276
rect 5244 2224 5296 2276
rect 5324 2224 5376 2276
rect 5024 2124 5076 2176
rect 5104 2124 5156 2176
rect 5244 2124 5296 2176
rect 5324 2124 5376 2176
<< metal2 >>
rect 1400 3500 2000 3900
rect 8400 3500 9000 3900
rect 1400 1800 1600 3500
rect 1700 2276 8700 2300
rect 1700 2224 5024 2276
rect 5076 2224 5104 2276
rect 5156 2224 5244 2276
rect 5296 2224 5324 2276
rect 5376 2224 8700 2276
rect 1700 2176 8700 2224
rect 1700 2124 5024 2176
rect 5076 2124 5104 2176
rect 5156 2124 5244 2176
rect 5296 2124 5324 2176
rect 5376 2124 8700 2176
rect 1700 2100 8700 2124
rect 1700 1800 1900 2100
rect 8500 1800 8700 2100
rect 8800 1800 9000 3500
rect 5100 -3320 5300 -1900
use differential-pair  differential-pair_0
timestamp 1770083657
transform 1 0 1100 0 1 -1600
box 300 -500 7900 3626
use mirror-load  mirror-load_0
timestamp 1770083657
transform 1 0 840 0 1 2540
box 900 -500 7800 2366
use y  y_0
timestamp 1770083657
transform 1 0 104 0 1 -3222
box 1800 -1800 8400 1126
<< end >>
