magic
tech sky130A
magscale 1 2
timestamp 1769411983
<< mvnmos >>
rect -1235 -502 -1135 440
rect -1077 -502 -977 440
rect -919 -502 -819 440
rect -761 -502 -661 440
rect -603 -502 -503 440
rect -445 -502 -345 440
rect -287 -502 -187 440
rect -129 -502 -29 440
rect 29 -502 129 440
rect 187 -502 287 440
rect 345 -502 445 440
rect 503 -502 603 440
rect 661 -502 761 440
rect 819 -502 919 440
rect 977 -502 1077 440
rect 1135 -502 1235 440
<< mvndiff >>
rect -1293 428 -1235 440
rect -1293 -490 -1281 428
rect -1247 -490 -1235 428
rect -1293 -502 -1235 -490
rect -1135 428 -1077 440
rect -1135 -490 -1123 428
rect -1089 -490 -1077 428
rect -1135 -502 -1077 -490
rect -977 428 -919 440
rect -977 -490 -965 428
rect -931 -490 -919 428
rect -977 -502 -919 -490
rect -819 428 -761 440
rect -819 -490 -807 428
rect -773 -490 -761 428
rect -819 -502 -761 -490
rect -661 428 -603 440
rect -661 -490 -649 428
rect -615 -490 -603 428
rect -661 -502 -603 -490
rect -503 428 -445 440
rect -503 -490 -491 428
rect -457 -490 -445 428
rect -503 -502 -445 -490
rect -345 428 -287 440
rect -345 -490 -333 428
rect -299 -490 -287 428
rect -345 -502 -287 -490
rect -187 428 -129 440
rect -187 -490 -175 428
rect -141 -490 -129 428
rect -187 -502 -129 -490
rect -29 428 29 440
rect -29 -490 -17 428
rect 17 -490 29 428
rect -29 -502 29 -490
rect 129 428 187 440
rect 129 -490 141 428
rect 175 -490 187 428
rect 129 -502 187 -490
rect 287 428 345 440
rect 287 -490 299 428
rect 333 -490 345 428
rect 287 -502 345 -490
rect 445 428 503 440
rect 445 -490 457 428
rect 491 -490 503 428
rect 445 -502 503 -490
rect 603 428 661 440
rect 603 -490 615 428
rect 649 -490 661 428
rect 603 -502 661 -490
rect 761 428 819 440
rect 761 -490 773 428
rect 807 -490 819 428
rect 761 -502 819 -490
rect 919 428 977 440
rect 919 -490 931 428
rect 965 -490 977 428
rect 919 -502 977 -490
rect 1077 428 1135 440
rect 1077 -490 1089 428
rect 1123 -490 1135 428
rect 1077 -502 1135 -490
rect 1235 428 1293 440
rect 1235 -490 1247 428
rect 1281 -490 1293 428
rect 1235 -502 1293 -490
<< mvndiffc >>
rect -1281 -490 -1247 428
rect -1123 -490 -1089 428
rect -965 -490 -931 428
rect -807 -490 -773 428
rect -649 -490 -615 428
rect -491 -490 -457 428
rect -333 -490 -299 428
rect -175 -490 -141 428
rect -17 -490 17 428
rect 141 -490 175 428
rect 299 -490 333 428
rect 457 -490 491 428
rect 615 -490 649 428
rect 773 -490 807 428
rect 931 -490 965 428
rect 1089 -490 1123 428
rect 1247 -490 1281 428
<< poly >>
rect -1235 512 -1135 528
rect -1235 478 -1219 512
rect -1151 478 -1135 512
rect -1235 440 -1135 478
rect -1077 512 -977 528
rect -1077 478 -1061 512
rect -993 478 -977 512
rect -1077 440 -977 478
rect -919 512 -819 528
rect -919 478 -903 512
rect -835 478 -819 512
rect -919 440 -819 478
rect -761 512 -661 528
rect -761 478 -745 512
rect -677 478 -661 512
rect -761 440 -661 478
rect -603 512 -503 528
rect -603 478 -587 512
rect -519 478 -503 512
rect -603 440 -503 478
rect -445 512 -345 528
rect -445 478 -429 512
rect -361 478 -345 512
rect -445 440 -345 478
rect -287 512 -187 528
rect -287 478 -271 512
rect -203 478 -187 512
rect -287 440 -187 478
rect -129 512 -29 528
rect -129 478 -113 512
rect -45 478 -29 512
rect -129 440 -29 478
rect 29 512 129 528
rect 29 478 45 512
rect 113 478 129 512
rect 29 440 129 478
rect 187 512 287 528
rect 187 478 203 512
rect 271 478 287 512
rect 187 440 287 478
rect 345 512 445 528
rect 345 478 361 512
rect 429 478 445 512
rect 345 440 445 478
rect 503 512 603 528
rect 503 478 519 512
rect 587 478 603 512
rect 503 440 603 478
rect 661 512 761 528
rect 661 478 677 512
rect 745 478 761 512
rect 661 440 761 478
rect 819 512 919 528
rect 819 478 835 512
rect 903 478 919 512
rect 819 440 919 478
rect 977 512 1077 528
rect 977 478 993 512
rect 1061 478 1077 512
rect 977 440 1077 478
rect 1135 512 1235 528
rect 1135 478 1151 512
rect 1219 478 1235 512
rect 1135 440 1235 478
rect -1235 -528 -1135 -502
rect -1077 -528 -977 -502
rect -919 -528 -819 -502
rect -761 -528 -661 -502
rect -603 -528 -503 -502
rect -445 -528 -345 -502
rect -287 -528 -187 -502
rect -129 -528 -29 -502
rect 29 -528 129 -502
rect 187 -528 287 -502
rect 345 -528 445 -502
rect 503 -528 603 -502
rect 661 -528 761 -502
rect 819 -528 919 -502
rect 977 -528 1077 -502
rect 1135 -528 1235 -502
<< polycont >>
rect -1219 478 -1151 512
rect -1061 478 -993 512
rect -903 478 -835 512
rect -745 478 -677 512
rect -587 478 -519 512
rect -429 478 -361 512
rect -271 478 -203 512
rect -113 478 -45 512
rect 45 478 113 512
rect 203 478 271 512
rect 361 478 429 512
rect 519 478 587 512
rect 677 478 745 512
rect 835 478 903 512
rect 993 478 1061 512
rect 1151 478 1219 512
<< locali >>
rect -1235 478 -1219 512
rect -1151 478 -1135 512
rect -1077 478 -1061 512
rect -993 478 -977 512
rect -919 478 -903 512
rect -835 478 -819 512
rect -761 478 -745 512
rect -677 478 -661 512
rect -603 478 -587 512
rect -519 478 -503 512
rect -445 478 -429 512
rect -361 478 -345 512
rect -287 478 -271 512
rect -203 478 -187 512
rect -129 478 -113 512
rect -45 478 -29 512
rect 29 478 45 512
rect 113 478 129 512
rect 187 478 203 512
rect 271 478 287 512
rect 345 478 361 512
rect 429 478 445 512
rect 503 478 519 512
rect 587 478 603 512
rect 661 478 677 512
rect 745 478 761 512
rect 819 478 835 512
rect 903 478 919 512
rect 977 478 993 512
rect 1061 478 1077 512
rect 1135 478 1151 512
rect 1219 478 1235 512
rect -1281 428 -1247 444
rect -1281 -506 -1247 -490
rect -1123 428 -1089 444
rect -1123 -506 -1089 -490
rect -965 428 -931 444
rect -965 -506 -931 -490
rect -807 428 -773 444
rect -807 -506 -773 -490
rect -649 428 -615 444
rect -649 -506 -615 -490
rect -491 428 -457 444
rect -491 -506 -457 -490
rect -333 428 -299 444
rect -333 -506 -299 -490
rect -175 428 -141 444
rect -175 -506 -141 -490
rect -17 428 17 444
rect -17 -506 17 -490
rect 141 428 175 444
rect 141 -506 175 -490
rect 299 428 333 444
rect 299 -506 333 -490
rect 457 428 491 444
rect 457 -506 491 -490
rect 615 428 649 444
rect 615 -506 649 -490
rect 773 428 807 444
rect 773 -506 807 -490
rect 931 428 965 444
rect 931 -506 965 -490
rect 1089 428 1123 444
rect 1089 -506 1123 -490
rect 1247 428 1281 444
rect 1247 -506 1281 -490
<< viali >>
rect -1219 478 -1151 512
rect -1061 478 -993 512
rect -903 478 -835 512
rect -745 478 -677 512
rect -587 478 -519 512
rect -429 478 -361 512
rect -271 478 -203 512
rect -113 478 -45 512
rect 45 478 113 512
rect 203 478 271 512
rect 361 478 429 512
rect 519 478 587 512
rect 677 478 745 512
rect 835 478 903 512
rect 993 478 1061 512
rect 1151 478 1219 512
rect -1281 -490 -1247 428
rect -1123 -490 -1089 428
rect -965 -490 -931 428
rect -807 -490 -773 428
rect -649 -490 -615 428
rect -491 -490 -457 428
rect -333 -490 -299 428
rect -175 -490 -141 428
rect -17 -490 17 428
rect 141 -490 175 428
rect 299 -490 333 428
rect 457 -490 491 428
rect 615 -490 649 428
rect 773 -490 807 428
rect 931 -490 965 428
rect 1089 -490 1123 428
rect 1247 -490 1281 428
<< metal1 >>
rect -1231 512 -1139 518
rect -1231 478 -1219 512
rect -1151 478 -1139 512
rect -1231 472 -1139 478
rect -1073 512 -981 518
rect -1073 478 -1061 512
rect -993 478 -981 512
rect -1073 472 -981 478
rect -915 512 -823 518
rect -915 478 -903 512
rect -835 478 -823 512
rect -915 472 -823 478
rect -757 512 -665 518
rect -757 478 -745 512
rect -677 478 -665 512
rect -757 472 -665 478
rect -599 512 -507 518
rect -599 478 -587 512
rect -519 478 -507 512
rect -599 472 -507 478
rect -441 512 -349 518
rect -441 478 -429 512
rect -361 478 -349 512
rect -441 472 -349 478
rect -283 512 -191 518
rect -283 478 -271 512
rect -203 478 -191 512
rect -283 472 -191 478
rect -125 512 -33 518
rect -125 478 -113 512
rect -45 478 -33 512
rect -125 472 -33 478
rect 33 512 125 518
rect 33 478 45 512
rect 113 478 125 512
rect 33 472 125 478
rect 191 512 283 518
rect 191 478 203 512
rect 271 478 283 512
rect 191 472 283 478
rect 349 512 441 518
rect 349 478 361 512
rect 429 478 441 512
rect 349 472 441 478
rect 507 512 599 518
rect 507 478 519 512
rect 587 478 599 512
rect 507 472 599 478
rect 665 512 757 518
rect 665 478 677 512
rect 745 478 757 512
rect 665 472 757 478
rect 823 512 915 518
rect 823 478 835 512
rect 903 478 915 512
rect 823 472 915 478
rect 981 512 1073 518
rect 981 478 993 512
rect 1061 478 1073 512
rect 981 472 1073 478
rect 1139 512 1231 518
rect 1139 478 1151 512
rect 1219 478 1231 512
rect 1139 472 1231 478
rect -1287 428 -1241 440
rect -1287 -490 -1281 428
rect -1247 -490 -1241 428
rect -1287 -502 -1241 -490
rect -1129 428 -1083 440
rect -1129 -490 -1123 428
rect -1089 -490 -1083 428
rect -1129 -502 -1083 -490
rect -971 428 -925 440
rect -971 -490 -965 428
rect -931 -490 -925 428
rect -971 -502 -925 -490
rect -813 428 -767 440
rect -813 -490 -807 428
rect -773 -490 -767 428
rect -813 -502 -767 -490
rect -655 428 -609 440
rect -655 -490 -649 428
rect -615 -490 -609 428
rect -655 -502 -609 -490
rect -497 428 -451 440
rect -497 -490 -491 428
rect -457 -490 -451 428
rect -497 -502 -451 -490
rect -339 428 -293 440
rect -339 -490 -333 428
rect -299 -490 -293 428
rect -339 -502 -293 -490
rect -181 428 -135 440
rect -181 -490 -175 428
rect -141 -490 -135 428
rect -181 -502 -135 -490
rect -23 428 23 440
rect -23 -490 -17 428
rect 17 -490 23 428
rect -23 -502 23 -490
rect 135 428 181 440
rect 135 -490 141 428
rect 175 -490 181 428
rect 135 -502 181 -490
rect 293 428 339 440
rect 293 -490 299 428
rect 333 -490 339 428
rect 293 -502 339 -490
rect 451 428 497 440
rect 451 -490 457 428
rect 491 -490 497 428
rect 451 -502 497 -490
rect 609 428 655 440
rect 609 -490 615 428
rect 649 -490 655 428
rect 609 -502 655 -490
rect 767 428 813 440
rect 767 -490 773 428
rect 807 -490 813 428
rect 767 -502 813 -490
rect 925 428 971 440
rect 925 -490 931 428
rect 965 -490 971 428
rect 925 -502 971 -490
rect 1083 428 1129 440
rect 1083 -490 1089 428
rect 1123 -490 1129 428
rect 1083 -502 1129 -490
rect 1241 428 1287 440
rect 1241 -490 1247 428
rect 1281 -490 1287 428
rect 1241 -502 1287 -490
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.7125 l 0.5 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
