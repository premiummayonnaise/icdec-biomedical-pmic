magic
tech sky130A
magscale 1 2
timestamp 1770112220
<< mvnmos >>
rect -587 -719 -337 781
rect -279 -719 -29 781
rect 29 -719 279 781
rect 337 -719 587 781
<< mvndiff >>
rect -645 769 -587 781
rect -645 -707 -633 769
rect -599 -707 -587 769
rect -645 -719 -587 -707
rect -337 769 -279 781
rect -337 -707 -325 769
rect -291 -707 -279 769
rect -337 -719 -279 -707
rect -29 769 29 781
rect -29 -707 -17 769
rect 17 -707 29 769
rect -29 -719 29 -707
rect 279 769 337 781
rect 279 -707 291 769
rect 325 -707 337 769
rect 279 -719 337 -707
rect 587 769 645 781
rect 587 -707 599 769
rect 633 -707 645 769
rect 587 -719 645 -707
<< mvndiffc >>
rect -633 -707 -599 769
rect -325 -707 -291 769
rect -17 -707 17 769
rect 291 -707 325 769
rect 599 -707 633 769
<< poly >>
rect -587 781 -337 807
rect -279 781 -29 807
rect 29 781 279 807
rect 337 781 587 807
rect -587 -757 -337 -719
rect -587 -791 -571 -757
rect -353 -791 -337 -757
rect -587 -807 -337 -791
rect -279 -757 -29 -719
rect -279 -791 -263 -757
rect -45 -791 -29 -757
rect -279 -807 -29 -791
rect 29 -757 279 -719
rect 29 -791 45 -757
rect 263 -791 279 -757
rect 29 -807 279 -791
rect 337 -757 587 -719
rect 337 -791 353 -757
rect 571 -791 587 -757
rect 337 -807 587 -791
<< polycont >>
rect -571 -791 -353 -757
rect -263 -791 -45 -757
rect 45 -791 263 -757
rect 353 -791 571 -757
<< locali >>
rect -633 769 -599 785
rect -633 -723 -599 -707
rect -325 769 -291 785
rect -325 -723 -291 -707
rect -17 769 17 785
rect -17 -723 17 -707
rect 291 769 325 785
rect 291 -723 325 -707
rect 599 769 633 785
rect 599 -723 633 -707
rect -587 -791 -571 -757
rect -353 -791 -337 -757
rect -279 -791 -263 -757
rect -45 -791 -29 -757
rect 29 -791 45 -757
rect 263 -791 279 -757
rect 337 -791 353 -757
rect 571 -791 587 -757
<< viali >>
rect -633 -707 -599 769
rect -325 -707 -291 769
rect -17 -707 17 769
rect 291 -707 325 769
rect 599 -707 633 769
rect -571 -791 -353 -757
rect -263 -791 -45 -757
rect 45 -791 263 -757
rect 353 -791 571 -757
<< metal1 >>
rect -639 769 -593 781
rect -639 -707 -633 769
rect -599 -707 -593 769
rect -639 -719 -593 -707
rect -331 769 -285 781
rect -331 -707 -325 769
rect -291 -707 -285 769
rect -331 -719 -285 -707
rect -23 769 23 781
rect -23 -707 -17 769
rect 17 -707 23 769
rect -23 -719 23 -707
rect 285 769 331 781
rect 285 -707 291 769
rect 325 -707 331 769
rect 285 -719 331 -707
rect 593 769 639 781
rect 593 -707 599 769
rect 633 -707 639 769
rect 593 -719 639 -707
rect -583 -757 -341 -751
rect -583 -791 -571 -757
rect -353 -791 -341 -757
rect -583 -797 -341 -791
rect -275 -757 -33 -751
rect -275 -791 -263 -757
rect -45 -791 -33 -757
rect -275 -797 -33 -791
rect 33 -757 275 -751
rect 33 -791 45 -757
rect 263 -791 275 -757
rect 33 -797 275 -791
rect 341 -757 583 -751
rect 341 -791 353 -757
rect 571 -791 583 -757
rect 341 -797 583 -791
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
