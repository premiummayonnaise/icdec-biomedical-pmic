magic
tech sky130A
magscale 1 2
timestamp 1768760819
<< mvnmos >>
rect -339 -189 -89 127
rect 89 -189 339 127
<< mvndiff >>
rect -397 115 -339 127
rect -397 -177 -385 115
rect -351 -177 -339 115
rect -397 -189 -339 -177
rect -89 115 -31 127
rect -89 -177 -77 115
rect -43 -177 -31 115
rect -89 -189 -31 -177
rect 31 115 89 127
rect 31 -177 43 115
rect 77 -177 89 115
rect 31 -189 89 -177
rect 339 115 397 127
rect 339 -177 351 115
rect 385 -177 397 115
rect 339 -189 397 -177
<< mvndiffc >>
rect -385 -177 -351 115
rect -77 -177 -43 115
rect 43 -177 77 115
rect 351 -177 385 115
<< poly >>
rect -339 199 -89 215
rect -339 165 -323 199
rect -105 165 -89 199
rect -339 127 -89 165
rect 89 199 339 215
rect 89 165 105 199
rect 323 165 339 199
rect 89 127 339 165
rect -339 -215 -89 -189
rect 89 -215 339 -189
<< polycont >>
rect -323 165 -105 199
rect 105 165 323 199
<< locali >>
rect -339 165 -323 199
rect -105 165 -89 199
rect 89 165 105 199
rect 323 165 339 199
rect -385 115 -351 131
rect -385 -193 -351 -177
rect -77 115 -43 131
rect -77 -193 -43 -177
rect 43 115 77 131
rect 43 -193 77 -177
rect 351 115 385 131
rect 351 -193 385 -177
<< viali >>
rect -323 165 -105 199
rect 105 165 323 199
rect -385 -177 -351 115
rect -77 -177 -43 115
rect 43 -177 77 115
rect 351 -177 385 115
<< metal1 >>
rect -335 199 -93 205
rect -335 165 -323 199
rect -105 165 -93 199
rect -335 159 -93 165
rect 93 199 335 205
rect 93 165 105 199
rect 323 165 335 199
rect 93 159 335 165
rect -391 115 -345 127
rect -391 -177 -385 115
rect -351 -177 -345 115
rect -391 -189 -345 -177
rect -83 115 -37 127
rect -83 -177 -77 115
rect -43 -177 -37 115
rect -83 -189 -37 -177
rect 37 115 83 127
rect 37 -177 43 115
rect 77 -177 83 115
rect 37 -189 83 -177
rect 345 115 391 127
rect 345 -177 351 115
rect 385 -177 391 115
rect 345 -189 391 -177
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.58 l 1.25 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
