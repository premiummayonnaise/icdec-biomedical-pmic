magic
tech sky130A
magscale 1 2
timestamp 1770117167
<< pwell >>
rect -280 -674 280 674
<< mvnmos >>
rect -50 -416 50 416
<< mvndiff >>
rect -108 404 -50 416
rect -108 -404 -96 404
rect -62 -404 -50 404
rect -108 -416 -50 -404
rect 50 404 108 416
rect 50 -404 62 404
rect 96 -404 108 404
rect 50 -416 108 -404
<< mvndiffc >>
rect -96 -404 -62 404
rect 62 -404 96 404
<< mvpsubdiff >>
rect -244 580 244 638
rect -244 530 -186 580
rect -244 -530 -232 530
rect -198 -530 -186 530
rect -244 -580 -186 -530
rect 186 -580 244 580
rect -244 -638 244 -580
<< mvpsubdiffcont >>
rect -232 -530 -198 530
<< poly >>
rect -50 488 50 504
rect -50 454 -34 488
rect 34 454 50 488
rect -50 416 50 454
rect -50 -454 50 -416
rect -50 -488 -34 -454
rect 34 -488 50 -454
rect -50 -504 50 -488
<< polycont >>
rect -34 454 34 488
rect -34 -488 34 -454
<< locali >>
rect -232 592 232 626
rect -232 530 -198 592
rect -50 454 -34 488
rect 34 454 50 488
rect -96 404 -62 420
rect -96 -420 -62 -404
rect 62 404 96 420
rect 62 -420 96 -404
rect -50 -488 -34 -454
rect 34 -488 50 -454
rect -232 -592 -198 -530
rect 198 -592 232 592
rect -232 -626 232 -592
<< viali >>
rect -34 454 34 488
rect -96 -404 -62 404
rect 62 -404 96 404
rect -34 -488 34 -454
<< metal1 >>
rect -46 488 46 494
rect -46 454 -34 488
rect 34 454 46 488
rect -46 448 46 454
rect -102 404 -56 416
rect -102 -404 -96 404
rect -62 -404 -56 404
rect -102 -416 -56 -404
rect 56 404 102 416
rect 56 -404 62 404
rect 96 -404 102 404
rect 56 -416 102 -404
rect -46 -454 46 -448
rect -46 -488 -34 -454
rect 34 -488 46 -454
rect -46 -494 46 -488
<< labels >>
rlabel mvpsubdiff 0 -609 0 -609 0 B
port 1 nsew
rlabel mvndiffc -79 0 -79 0 0 D
port 2 nsew
rlabel mvndiffc 79 0 79 0 0 S
port 3 nsew
rlabel polycont 0 471 0 471 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -215 -609 215 609
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.16 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
