magic
tech sky130A
magscale 1 2
timestamp 1770134472
<< pwell >>
rect -617 -527 617 527
<< mvnmos >>
rect -387 -269 -237 331
rect -179 -269 -29 331
rect 29 -269 179 331
rect 237 -269 387 331
<< mvndiff >>
rect -445 319 -387 331
rect -445 -257 -433 319
rect -399 -257 -387 319
rect -445 -269 -387 -257
rect -237 319 -179 331
rect -237 -257 -225 319
rect -191 -257 -179 319
rect -237 -269 -179 -257
rect -29 319 29 331
rect -29 -257 -17 319
rect 17 -257 29 319
rect -29 -269 29 -257
rect 179 319 237 331
rect 179 -257 191 319
rect 225 -257 237 319
rect 179 -269 237 -257
rect 387 319 445 331
rect 387 -257 399 319
rect 433 -257 445 319
rect 387 -269 445 -257
<< mvndiffc >>
rect -433 -257 -399 319
rect -225 -257 -191 319
rect -17 -257 17 319
rect 191 -257 225 319
rect 399 -257 433 319
<< mvpsubdiff >>
rect -581 479 581 491
rect -581 445 -473 479
rect 473 445 581 479
rect -581 433 581 445
rect -581 -433 -523 433
rect 523 -433 581 433
rect -581 -445 581 -433
rect -581 -479 -473 -445
rect 473 -479 581 -445
rect -581 -491 581 -479
<< mvpsubdiffcont >>
rect -473 445 473 479
rect -473 -479 473 -445
<< poly >>
rect -387 331 -237 357
rect -179 331 -29 357
rect 29 331 179 357
rect 237 331 387 357
rect -387 -307 -237 -269
rect -387 -341 -371 -307
rect -253 -341 -237 -307
rect -387 -357 -237 -341
rect -179 -307 -29 -269
rect -179 -341 -163 -307
rect -45 -341 -29 -307
rect -179 -357 -29 -341
rect 29 -307 179 -269
rect 29 -341 45 -307
rect 163 -341 179 -307
rect 29 -357 179 -341
rect 237 -307 387 -269
rect 237 -341 253 -307
rect 371 -341 387 -307
rect 237 -357 387 -341
<< polycont >>
rect -371 -341 -253 -307
rect -163 -341 -45 -307
rect 45 -341 163 -307
rect 253 -341 371 -307
<< locali >>
rect -569 445 -473 479
rect 473 445 569 479
rect -569 -445 -535 445
rect -433 319 -399 335
rect -433 -273 -399 -257
rect -225 319 -191 335
rect -225 -273 -191 -257
rect -17 319 17 335
rect -17 -273 17 -257
rect 191 319 225 335
rect 191 -273 225 -257
rect 399 319 433 335
rect 399 -273 433 -257
rect -387 -341 -371 -307
rect -253 -341 -237 -307
rect -179 -341 -163 -307
rect -45 -341 -29 -307
rect 29 -341 45 -307
rect 163 -341 179 -307
rect 237 -341 253 -307
rect 371 -341 387 -307
rect 535 -445 569 445
rect -569 -479 -473 -445
rect 473 -479 569 -445
<< viali >>
rect -433 -257 -399 319
rect -225 -257 -191 319
rect -17 -257 17 319
rect 191 -257 225 319
rect 399 -257 433 319
rect -371 -341 -253 -307
rect -163 -341 -45 -307
rect 45 -341 163 -307
rect 253 -341 371 -307
<< metal1 >>
rect -439 319 -393 331
rect -439 -257 -433 319
rect -399 -257 -393 319
rect -439 -269 -393 -257
rect -231 319 -185 331
rect -231 -257 -225 319
rect -191 -257 -185 319
rect -231 -269 -185 -257
rect -23 319 23 331
rect -23 -257 -17 319
rect 17 -257 23 319
rect -23 -269 23 -257
rect 185 319 231 331
rect 185 -257 191 319
rect 225 -257 231 319
rect 185 -269 231 -257
rect 393 319 439 331
rect 393 -257 399 319
rect 433 -257 439 319
rect 393 -269 439 -257
rect -383 -307 -241 -301
rect -383 -341 -371 -307
rect -253 -341 -241 -307
rect -383 -347 -241 -341
rect -175 -307 -33 -301
rect -175 -341 -163 -307
rect -45 -341 -33 -307
rect -175 -347 -33 -341
rect 33 -307 175 -301
rect 33 -341 45 -307
rect 163 -341 175 -307
rect 33 -347 175 -341
rect 241 -307 383 -301
rect 241 -341 253 -307
rect 371 -341 383 -307
rect 241 -347 383 -341
<< labels >>
rlabel mvpsubdiffcont 0 -462 0 -462 0 B
port 1 nsew
rlabel mvndiffc -416 31 -416 31 0 D0
port 2 nsew
rlabel polycont -312 -324 -312 -324 0 G0
port 3 nsew
rlabel mvndiffc -208 31 -208 31 0 S1
port 4 nsew
rlabel polycont -104 -324 -104 -324 0 G1
port 5 nsew
rlabel mvndiffc 0 31 0 31 0 D2
port 6 nsew
rlabel polycont 104 -324 104 -324 0 G2
port 7 nsew
rlabel mvndiffc 208 31 208 31 0 S3
port 8 nsew
rlabel polycont 312 -324 312 -324 0 G3
port 9 nsew
<< properties >>
string FIXED_BBOX -552 -462 552 462
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 0.75 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
