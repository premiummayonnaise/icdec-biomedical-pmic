magic
tech sky130A
magscale 1 2
timestamp 1770112220
<< pwell >>
rect -2663 -1008 2663 1008
<< mvnmos >>
rect -2435 -750 -2185 750
rect -2127 -750 -1877 750
rect -1819 -750 -1569 750
rect -1511 -750 -1261 750
rect -1203 -750 -953 750
rect -895 -750 -645 750
rect -587 -750 -337 750
rect -279 -750 -29 750
rect 29 -750 279 750
rect 337 -750 587 750
rect 645 -750 895 750
rect 953 -750 1203 750
rect 1261 -750 1511 750
rect 1569 -750 1819 750
rect 1877 -750 2127 750
rect 2185 -750 2435 750
<< mvndiff >>
rect -2493 738 -2435 750
rect -2493 -738 -2481 738
rect -2447 -738 -2435 738
rect -2493 -750 -2435 -738
rect -2185 738 -2127 750
rect -2185 -738 -2173 738
rect -2139 -738 -2127 738
rect -2185 -750 -2127 -738
rect -1877 738 -1819 750
rect -1877 -738 -1865 738
rect -1831 -738 -1819 738
rect -1877 -750 -1819 -738
rect -1569 738 -1511 750
rect -1569 -738 -1557 738
rect -1523 -738 -1511 738
rect -1569 -750 -1511 -738
rect -1261 738 -1203 750
rect -1261 -738 -1249 738
rect -1215 -738 -1203 738
rect -1261 -750 -1203 -738
rect -953 738 -895 750
rect -953 -738 -941 738
rect -907 -738 -895 738
rect -953 -750 -895 -738
rect -645 738 -587 750
rect -645 -738 -633 738
rect -599 -738 -587 738
rect -645 -750 -587 -738
rect -337 738 -279 750
rect -337 -738 -325 738
rect -291 -738 -279 738
rect -337 -750 -279 -738
rect -29 738 29 750
rect -29 -738 -17 738
rect 17 -738 29 738
rect -29 -750 29 -738
rect 279 738 337 750
rect 279 -738 291 738
rect 325 -738 337 738
rect 279 -750 337 -738
rect 587 738 645 750
rect 587 -738 599 738
rect 633 -738 645 738
rect 587 -750 645 -738
rect 895 738 953 750
rect 895 -738 907 738
rect 941 -738 953 738
rect 895 -750 953 -738
rect 1203 738 1261 750
rect 1203 -738 1215 738
rect 1249 -738 1261 738
rect 1203 -750 1261 -738
rect 1511 738 1569 750
rect 1511 -738 1523 738
rect 1557 -738 1569 738
rect 1511 -750 1569 -738
rect 1819 738 1877 750
rect 1819 -738 1831 738
rect 1865 -738 1877 738
rect 1819 -750 1877 -738
rect 2127 738 2185 750
rect 2127 -738 2139 738
rect 2173 -738 2185 738
rect 2127 -750 2185 -738
rect 2435 738 2493 750
rect 2435 -738 2447 738
rect 2481 -738 2493 738
rect 2435 -750 2493 -738
<< mvndiffc >>
rect -2481 -738 -2447 738
rect -2173 -738 -2139 738
rect -1865 -738 -1831 738
rect -1557 -738 -1523 738
rect -1249 -738 -1215 738
rect -941 -738 -907 738
rect -633 -738 -599 738
rect -325 -738 -291 738
rect -17 -738 17 738
rect 291 -738 325 738
rect 599 -738 633 738
rect 907 -738 941 738
rect 1215 -738 1249 738
rect 1523 -738 1557 738
rect 1831 -738 1865 738
rect 2139 -738 2173 738
rect 2447 -738 2481 738
<< mvpsubdiff >>
rect -2627 960 2627 972
rect -2627 926 -2519 960
rect 2519 926 2627 960
rect -2627 914 2627 926
rect -2627 864 -2569 914
rect -2627 -864 -2615 864
rect -2581 -864 -2569 864
rect 2569 864 2627 914
rect -2627 -914 -2569 -864
rect 2569 -864 2581 864
rect 2615 -864 2627 864
rect 2569 -914 2627 -864
rect -2627 -926 2627 -914
rect -2627 -960 -2519 -926
rect 2519 -960 2627 -926
rect -2627 -972 2627 -960
<< mvpsubdiffcont >>
rect -2519 926 2519 960
rect -2615 -864 -2581 864
rect 2581 -864 2615 864
rect -2519 -960 2519 -926
<< poly >>
rect -2435 822 -2185 838
rect -2435 788 -2419 822
rect -2201 788 -2185 822
rect -2435 750 -2185 788
rect -2127 822 -1877 838
rect -2127 788 -2111 822
rect -1893 788 -1877 822
rect -2127 750 -1877 788
rect -1819 822 -1569 838
rect -1819 788 -1803 822
rect -1585 788 -1569 822
rect -1819 750 -1569 788
rect -1511 822 -1261 838
rect -1511 788 -1495 822
rect -1277 788 -1261 822
rect -1511 750 -1261 788
rect -1203 822 -953 838
rect -1203 788 -1187 822
rect -969 788 -953 822
rect -1203 750 -953 788
rect -895 822 -645 838
rect -895 788 -879 822
rect -661 788 -645 822
rect -895 750 -645 788
rect -587 822 -337 838
rect -587 788 -571 822
rect -353 788 -337 822
rect -587 750 -337 788
rect -279 822 -29 838
rect -279 788 -263 822
rect -45 788 -29 822
rect -279 750 -29 788
rect 29 822 279 838
rect 29 788 45 822
rect 263 788 279 822
rect 29 750 279 788
rect 337 822 587 838
rect 337 788 353 822
rect 571 788 587 822
rect 337 750 587 788
rect 645 822 895 838
rect 645 788 661 822
rect 879 788 895 822
rect 645 750 895 788
rect 953 822 1203 838
rect 953 788 969 822
rect 1187 788 1203 822
rect 953 750 1203 788
rect 1261 822 1511 838
rect 1261 788 1277 822
rect 1495 788 1511 822
rect 1261 750 1511 788
rect 1569 822 1819 838
rect 1569 788 1585 822
rect 1803 788 1819 822
rect 1569 750 1819 788
rect 1877 822 2127 838
rect 1877 788 1893 822
rect 2111 788 2127 822
rect 1877 750 2127 788
rect 2185 822 2435 838
rect 2185 788 2201 822
rect 2419 788 2435 822
rect 2185 750 2435 788
rect -2435 -788 -2185 -750
rect -2435 -822 -2419 -788
rect -2201 -822 -2185 -788
rect -2435 -838 -2185 -822
rect -2127 -788 -1877 -750
rect -2127 -822 -2111 -788
rect -1893 -822 -1877 -788
rect -2127 -838 -1877 -822
rect -1819 -788 -1569 -750
rect -1819 -822 -1803 -788
rect -1585 -822 -1569 -788
rect -1819 -838 -1569 -822
rect -1511 -788 -1261 -750
rect -1511 -822 -1495 -788
rect -1277 -822 -1261 -788
rect -1511 -838 -1261 -822
rect -1203 -788 -953 -750
rect -1203 -822 -1187 -788
rect -969 -822 -953 -788
rect -1203 -838 -953 -822
rect -895 -788 -645 -750
rect -895 -822 -879 -788
rect -661 -822 -645 -788
rect -895 -838 -645 -822
rect -587 -788 -337 -750
rect -587 -822 -571 -788
rect -353 -822 -337 -788
rect -587 -838 -337 -822
rect -279 -788 -29 -750
rect -279 -822 -263 -788
rect -45 -822 -29 -788
rect -279 -838 -29 -822
rect 29 -788 279 -750
rect 29 -822 45 -788
rect 263 -822 279 -788
rect 29 -838 279 -822
rect 337 -788 587 -750
rect 337 -822 353 -788
rect 571 -822 587 -788
rect 337 -838 587 -822
rect 645 -788 895 -750
rect 645 -822 661 -788
rect 879 -822 895 -788
rect 645 -838 895 -822
rect 953 -788 1203 -750
rect 953 -822 969 -788
rect 1187 -822 1203 -788
rect 953 -838 1203 -822
rect 1261 -788 1511 -750
rect 1261 -822 1277 -788
rect 1495 -822 1511 -788
rect 1261 -838 1511 -822
rect 1569 -788 1819 -750
rect 1569 -822 1585 -788
rect 1803 -822 1819 -788
rect 1569 -838 1819 -822
rect 1877 -788 2127 -750
rect 1877 -822 1893 -788
rect 2111 -822 2127 -788
rect 1877 -838 2127 -822
rect 2185 -788 2435 -750
rect 2185 -822 2201 -788
rect 2419 -822 2435 -788
rect 2185 -838 2435 -822
<< polycont >>
rect -2419 788 -2201 822
rect -2111 788 -1893 822
rect -1803 788 -1585 822
rect -1495 788 -1277 822
rect -1187 788 -969 822
rect -879 788 -661 822
rect -571 788 -353 822
rect -263 788 -45 822
rect 45 788 263 822
rect 353 788 571 822
rect 661 788 879 822
rect 969 788 1187 822
rect 1277 788 1495 822
rect 1585 788 1803 822
rect 1893 788 2111 822
rect 2201 788 2419 822
rect -2419 -822 -2201 -788
rect -2111 -822 -1893 -788
rect -1803 -822 -1585 -788
rect -1495 -822 -1277 -788
rect -1187 -822 -969 -788
rect -879 -822 -661 -788
rect -571 -822 -353 -788
rect -263 -822 -45 -788
rect 45 -822 263 -788
rect 353 -822 571 -788
rect 661 -822 879 -788
rect 969 -822 1187 -788
rect 1277 -822 1495 -788
rect 1585 -822 1803 -788
rect 1893 -822 2111 -788
rect 2201 -822 2419 -788
<< locali >>
rect -2615 926 -2519 960
rect 2519 926 2615 960
rect -2615 864 -2581 926
rect 2581 864 2615 926
rect -2435 788 -2419 822
rect -2201 788 -2185 822
rect -2127 788 -2111 822
rect -1893 788 -1877 822
rect -1819 788 -1803 822
rect -1585 788 -1569 822
rect -1511 788 -1495 822
rect -1277 788 -1261 822
rect -1203 788 -1187 822
rect -969 788 -953 822
rect -895 788 -879 822
rect -661 788 -645 822
rect -587 788 -571 822
rect -353 788 -337 822
rect -279 788 -263 822
rect -45 788 -29 822
rect 29 788 45 822
rect 263 788 279 822
rect 337 788 353 822
rect 571 788 587 822
rect 645 788 661 822
rect 879 788 895 822
rect 953 788 969 822
rect 1187 788 1203 822
rect 1261 788 1277 822
rect 1495 788 1511 822
rect 1569 788 1585 822
rect 1803 788 1819 822
rect 1877 788 1893 822
rect 2111 788 2127 822
rect 2185 788 2201 822
rect 2419 788 2435 822
rect -2481 738 -2447 754
rect -2481 -754 -2447 -738
rect -2173 738 -2139 754
rect -2173 -754 -2139 -738
rect -1865 738 -1831 754
rect -1865 -754 -1831 -738
rect -1557 738 -1523 754
rect -1557 -754 -1523 -738
rect -1249 738 -1215 754
rect -1249 -754 -1215 -738
rect -941 738 -907 754
rect -941 -754 -907 -738
rect -633 738 -599 754
rect -633 -754 -599 -738
rect -325 738 -291 754
rect -325 -754 -291 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 291 738 325 754
rect 291 -754 325 -738
rect 599 738 633 754
rect 599 -754 633 -738
rect 907 738 941 754
rect 907 -754 941 -738
rect 1215 738 1249 754
rect 1215 -754 1249 -738
rect 1523 738 1557 754
rect 1523 -754 1557 -738
rect 1831 738 1865 754
rect 1831 -754 1865 -738
rect 2139 738 2173 754
rect 2139 -754 2173 -738
rect 2447 738 2481 754
rect 2447 -754 2481 -738
rect -2435 -822 -2419 -788
rect -2201 -822 -2185 -788
rect -2127 -822 -2111 -788
rect -1893 -822 -1877 -788
rect -1819 -822 -1803 -788
rect -1585 -822 -1569 -788
rect -1511 -822 -1495 -788
rect -1277 -822 -1261 -788
rect -1203 -822 -1187 -788
rect -969 -822 -953 -788
rect -895 -822 -879 -788
rect -661 -822 -645 -788
rect -587 -822 -571 -788
rect -353 -822 -337 -788
rect -279 -822 -263 -788
rect -45 -822 -29 -788
rect 29 -822 45 -788
rect 263 -822 279 -788
rect 337 -822 353 -788
rect 571 -822 587 -788
rect 645 -822 661 -788
rect 879 -822 895 -788
rect 953 -822 969 -788
rect 1187 -822 1203 -788
rect 1261 -822 1277 -788
rect 1495 -822 1511 -788
rect 1569 -822 1585 -788
rect 1803 -822 1819 -788
rect 1877 -822 1893 -788
rect 2111 -822 2127 -788
rect 2185 -822 2201 -788
rect 2419 -822 2435 -788
rect -2615 -926 -2581 -864
rect 2581 -926 2615 -864
rect -2615 -960 -2519 -926
rect 2519 -960 2615 -926
<< viali >>
rect -2419 788 -2201 822
rect -2111 788 -1893 822
rect -1803 788 -1585 822
rect -1495 788 -1277 822
rect -1187 788 -969 822
rect -879 788 -661 822
rect -571 788 -353 822
rect -263 788 -45 822
rect 45 788 263 822
rect 353 788 571 822
rect 661 788 879 822
rect 969 788 1187 822
rect 1277 788 1495 822
rect 1585 788 1803 822
rect 1893 788 2111 822
rect 2201 788 2419 822
rect -2481 -738 -2447 738
rect -2173 -738 -2139 738
rect -1865 -738 -1831 738
rect -1557 -738 -1523 738
rect -1249 -738 -1215 738
rect -941 -738 -907 738
rect -633 -738 -599 738
rect -325 -738 -291 738
rect -17 -738 17 738
rect 291 -738 325 738
rect 599 -738 633 738
rect 907 -738 941 738
rect 1215 -738 1249 738
rect 1523 -738 1557 738
rect 1831 -738 1865 738
rect 2139 -738 2173 738
rect 2447 -738 2481 738
rect -2419 -822 -2201 -788
rect -2111 -822 -1893 -788
rect -1803 -822 -1585 -788
rect -1495 -822 -1277 -788
rect -1187 -822 -969 -788
rect -879 -822 -661 -788
rect -571 -822 -353 -788
rect -263 -822 -45 -788
rect 45 -822 263 -788
rect 353 -822 571 -788
rect 661 -822 879 -788
rect 969 -822 1187 -788
rect 1277 -822 1495 -788
rect 1585 -822 1803 -788
rect 1893 -822 2111 -788
rect 2201 -822 2419 -788
<< metal1 >>
rect -2431 822 -2189 828
rect -2431 788 -2419 822
rect -2201 788 -2189 822
rect -2431 782 -2189 788
rect -2123 822 -1881 828
rect -2123 788 -2111 822
rect -1893 788 -1881 822
rect -2123 782 -1881 788
rect -1815 822 -1573 828
rect -1815 788 -1803 822
rect -1585 788 -1573 822
rect -1815 782 -1573 788
rect -1507 822 -1265 828
rect -1507 788 -1495 822
rect -1277 788 -1265 822
rect -1507 782 -1265 788
rect -1199 822 -957 828
rect -1199 788 -1187 822
rect -969 788 -957 822
rect -1199 782 -957 788
rect -891 822 -649 828
rect -891 788 -879 822
rect -661 788 -649 822
rect -891 782 -649 788
rect -583 822 -341 828
rect -583 788 -571 822
rect -353 788 -341 822
rect -583 782 -341 788
rect -275 822 -33 828
rect -275 788 -263 822
rect -45 788 -33 822
rect -275 782 -33 788
rect 33 822 275 828
rect 33 788 45 822
rect 263 788 275 822
rect 33 782 275 788
rect 341 822 583 828
rect 341 788 353 822
rect 571 788 583 822
rect 341 782 583 788
rect 649 822 891 828
rect 649 788 661 822
rect 879 788 891 822
rect 649 782 891 788
rect 957 822 1199 828
rect 957 788 969 822
rect 1187 788 1199 822
rect 957 782 1199 788
rect 1265 822 1507 828
rect 1265 788 1277 822
rect 1495 788 1507 822
rect 1265 782 1507 788
rect 1573 822 1815 828
rect 1573 788 1585 822
rect 1803 788 1815 822
rect 1573 782 1815 788
rect 1881 822 2123 828
rect 1881 788 1893 822
rect 2111 788 2123 822
rect 1881 782 2123 788
rect 2189 822 2431 828
rect 2189 788 2201 822
rect 2419 788 2431 822
rect 2189 782 2431 788
rect -2487 738 -2441 750
rect -2487 -738 -2481 738
rect -2447 -738 -2441 738
rect -2487 -750 -2441 -738
rect -2179 738 -2133 750
rect -2179 -738 -2173 738
rect -2139 -738 -2133 738
rect -2179 -750 -2133 -738
rect -1871 738 -1825 750
rect -1871 -738 -1865 738
rect -1831 -738 -1825 738
rect -1871 -750 -1825 -738
rect -1563 738 -1517 750
rect -1563 -738 -1557 738
rect -1523 -738 -1517 738
rect -1563 -750 -1517 -738
rect -1255 738 -1209 750
rect -1255 -738 -1249 738
rect -1215 -738 -1209 738
rect -1255 -750 -1209 -738
rect -947 738 -901 750
rect -947 -738 -941 738
rect -907 -738 -901 738
rect -947 -750 -901 -738
rect -639 738 -593 750
rect -639 -738 -633 738
rect -599 -738 -593 738
rect -639 -750 -593 -738
rect -331 738 -285 750
rect -331 -738 -325 738
rect -291 -738 -285 738
rect -331 -750 -285 -738
rect -23 738 23 750
rect -23 -738 -17 738
rect 17 -738 23 738
rect -23 -750 23 -738
rect 285 738 331 750
rect 285 -738 291 738
rect 325 -738 331 738
rect 285 -750 331 -738
rect 593 738 639 750
rect 593 -738 599 738
rect 633 -738 639 738
rect 593 -750 639 -738
rect 901 738 947 750
rect 901 -738 907 738
rect 941 -738 947 738
rect 901 -750 947 -738
rect 1209 738 1255 750
rect 1209 -738 1215 738
rect 1249 -738 1255 738
rect 1209 -750 1255 -738
rect 1517 738 1563 750
rect 1517 -738 1523 738
rect 1557 -738 1563 738
rect 1517 -750 1563 -738
rect 1825 738 1871 750
rect 1825 -738 1831 738
rect 1865 -738 1871 738
rect 1825 -750 1871 -738
rect 2133 738 2179 750
rect 2133 -738 2139 738
rect 2173 -738 2179 738
rect 2133 -750 2179 -738
rect 2441 738 2487 750
rect 2441 -738 2447 738
rect 2481 -738 2487 738
rect 2441 -750 2487 -738
rect -2431 -788 -2189 -782
rect -2431 -822 -2419 -788
rect -2201 -822 -2189 -788
rect -2431 -828 -2189 -822
rect -2123 -788 -1881 -782
rect -2123 -822 -2111 -788
rect -1893 -822 -1881 -788
rect -2123 -828 -1881 -822
rect -1815 -788 -1573 -782
rect -1815 -822 -1803 -788
rect -1585 -822 -1573 -788
rect -1815 -828 -1573 -822
rect -1507 -788 -1265 -782
rect -1507 -822 -1495 -788
rect -1277 -822 -1265 -788
rect -1507 -828 -1265 -822
rect -1199 -788 -957 -782
rect -1199 -822 -1187 -788
rect -969 -822 -957 -788
rect -1199 -828 -957 -822
rect -891 -788 -649 -782
rect -891 -822 -879 -788
rect -661 -822 -649 -788
rect -891 -828 -649 -822
rect -583 -788 -341 -782
rect -583 -822 -571 -788
rect -353 -822 -341 -788
rect -583 -828 -341 -822
rect -275 -788 -33 -782
rect -275 -822 -263 -788
rect -45 -822 -33 -788
rect -275 -828 -33 -822
rect 33 -788 275 -782
rect 33 -822 45 -788
rect 263 -822 275 -788
rect 33 -828 275 -822
rect 341 -788 583 -782
rect 341 -822 353 -788
rect 571 -822 583 -788
rect 341 -828 583 -822
rect 649 -788 891 -782
rect 649 -822 661 -788
rect 879 -822 891 -788
rect 649 -828 891 -822
rect 957 -788 1199 -782
rect 957 -822 969 -788
rect 1187 -822 1199 -788
rect 957 -828 1199 -822
rect 1265 -788 1507 -782
rect 1265 -822 1277 -788
rect 1495 -822 1507 -788
rect 1265 -828 1507 -822
rect 1573 -788 1815 -782
rect 1573 -822 1585 -788
rect 1803 -822 1815 -788
rect 1573 -828 1815 -822
rect 1881 -788 2123 -782
rect 1881 -822 1893 -788
rect 2111 -822 2123 -788
rect 1881 -828 2123 -822
rect 2189 -788 2431 -782
rect 2189 -822 2201 -788
rect 2419 -822 2431 -788
rect 2189 -828 2431 -822
<< properties >>
string FIXED_BBOX -2598 -943 2598 943
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
