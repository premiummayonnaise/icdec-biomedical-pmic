magic
tech sky130A
magscale 1 2
timestamp 1769400417
<< metal3 >>
rect -4492 4172 -120 4200
rect -4492 148 -204 4172
rect -140 148 -120 4172
rect -4492 120 -120 148
rect 120 4172 4492 4200
rect 120 148 4408 4172
rect 4472 148 4492 4172
rect 120 120 4492 148
rect -4492 -148 -120 -120
rect -4492 -4172 -204 -148
rect -140 -4172 -120 -148
rect -4492 -4200 -120 -4172
rect 120 -148 4492 -120
rect 120 -4172 4408 -148
rect 4472 -4172 4492 -148
rect 120 -4200 4492 -4172
<< via3 >>
rect -204 148 -140 4172
rect 4408 148 4472 4172
rect -204 -4172 -140 -148
rect 4408 -4172 4472 -148
<< mimcap >>
rect -4452 4120 -452 4160
rect -4452 200 -4412 4120
rect -492 200 -452 4120
rect -4452 160 -452 200
rect 160 4120 4160 4160
rect 160 200 200 4120
rect 4120 200 4160 4120
rect 160 160 4160 200
rect -4452 -200 -452 -160
rect -4452 -4120 -4412 -200
rect -492 -4120 -452 -200
rect -4452 -4160 -452 -4120
rect 160 -200 4160 -160
rect 160 -4120 200 -200
rect 4120 -4120 4160 -200
rect 160 -4160 4160 -4120
<< mimcapcontact >>
rect -4412 200 -492 4120
rect 200 200 4120 4120
rect -4412 -4120 -492 -200
rect 200 -4120 4120 -200
<< metal4 >>
rect -2504 4121 -2400 4320
rect -224 4172 -120 4320
rect -4413 4120 -491 4121
rect -4413 200 -4412 4120
rect -492 200 -491 4120
rect -4413 199 -491 200
rect -2504 -199 -2400 199
rect -224 148 -204 4172
rect -140 148 -120 4172
rect 2108 4121 2212 4320
rect 4388 4172 4492 4320
rect 199 4120 4121 4121
rect 199 200 200 4120
rect 4120 200 4121 4120
rect 199 199 4121 200
rect -224 -148 -120 148
rect -4413 -200 -491 -199
rect -4413 -4120 -4412 -200
rect -492 -4120 -491 -200
rect -4413 -4121 -491 -4120
rect -2504 -4320 -2400 -4121
rect -224 -4172 -204 -148
rect -140 -4172 -120 -148
rect 2108 -199 2212 199
rect 4388 148 4408 4172
rect 4472 148 4492 4172
rect 4388 -148 4492 148
rect 199 -200 4121 -199
rect 199 -4120 200 -200
rect 4120 -4120 4121 -200
rect 199 -4121 4121 -4120
rect -224 -4320 -120 -4172
rect 2108 -4320 2212 -4121
rect 4388 -4172 4408 -148
rect 4472 -4172 4492 -148
rect 4388 -4320 4492 -4172
<< properties >>
string FIXED_BBOX 120 120 4200 4200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20.0 l 20.0 val 815.2 carea 2.00 cperi 0.19 class capacitor nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
