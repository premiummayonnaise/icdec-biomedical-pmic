magic
tech sky130A
magscale 1 2
timestamp 1769436194
<< metal3 >>
rect -5492 10492 -120 10520
rect -5492 5468 -204 10492
rect -140 5468 -120 10492
rect -5492 5440 -120 5468
rect 120 10492 5492 10520
rect 120 5468 5408 10492
rect 5472 5468 5492 10492
rect 120 5440 5492 5468
rect -5492 5172 -120 5200
rect -5492 148 -204 5172
rect -140 148 -120 5172
rect -5492 120 -120 148
rect 120 5172 5492 5200
rect 120 148 5408 5172
rect 5472 148 5492 5172
rect 120 120 5492 148
rect -5492 -148 -120 -120
rect -5492 -5172 -204 -148
rect -140 -5172 -120 -148
rect -5492 -5200 -120 -5172
rect 120 -148 5492 -120
rect 120 -5172 5408 -148
rect 5472 -5172 5492 -148
rect 120 -5200 5492 -5172
rect -5492 -5468 -120 -5440
rect -5492 -10492 -204 -5468
rect -140 -10492 -120 -5468
rect -5492 -10520 -120 -10492
rect 120 -5468 5492 -5440
rect 120 -10492 5408 -5468
rect 5472 -10492 5492 -5468
rect 120 -10520 5492 -10492
<< via3 >>
rect -204 5468 -140 10492
rect 5408 5468 5472 10492
rect -204 148 -140 5172
rect 5408 148 5472 5172
rect -204 -5172 -140 -148
rect 5408 -5172 5472 -148
rect -204 -10492 -140 -5468
rect 5408 -10492 5472 -5468
<< mimcap >>
rect -5452 10440 -452 10480
rect -5452 5520 -5412 10440
rect -492 5520 -452 10440
rect -5452 5480 -452 5520
rect 160 10440 5160 10480
rect 160 5520 200 10440
rect 5120 5520 5160 10440
rect 160 5480 5160 5520
rect -5452 5120 -452 5160
rect -5452 200 -5412 5120
rect -492 200 -452 5120
rect -5452 160 -452 200
rect 160 5120 5160 5160
rect 160 200 200 5120
rect 5120 200 5160 5120
rect 160 160 5160 200
rect -5452 -200 -452 -160
rect -5452 -5120 -5412 -200
rect -492 -5120 -452 -200
rect -5452 -5160 -452 -5120
rect 160 -200 5160 -160
rect 160 -5120 200 -200
rect 5120 -5120 5160 -200
rect 160 -5160 5160 -5120
rect -5452 -5520 -452 -5480
rect -5452 -10440 -5412 -5520
rect -492 -10440 -452 -5520
rect -5452 -10480 -452 -10440
rect 160 -5520 5160 -5480
rect 160 -10440 200 -5520
rect 5120 -10440 5160 -5520
rect 160 -10480 5160 -10440
<< mimcapcontact >>
rect -5412 5520 -492 10440
rect 200 5520 5120 10440
rect -5412 200 -492 5120
rect 200 200 5120 5120
rect -5412 -5120 -492 -200
rect 200 -5120 5120 -200
rect -5412 -10440 -492 -5520
rect 200 -10440 5120 -5520
<< metal4 >>
rect -3004 10441 -2900 10640
rect -224 10492 -120 10640
rect -5413 10440 -491 10441
rect -5413 5520 -5412 10440
rect -492 5520 -491 10440
rect -5413 5519 -491 5520
rect -3004 5121 -2900 5519
rect -224 5468 -204 10492
rect -140 5468 -120 10492
rect 2608 10441 2712 10640
rect 5388 10492 5492 10640
rect 199 10440 5121 10441
rect 199 5520 200 10440
rect 5120 5520 5121 10440
rect 199 5519 5121 5520
rect -224 5172 -120 5468
rect -5413 5120 -491 5121
rect -5413 200 -5412 5120
rect -492 200 -491 5120
rect -5413 199 -491 200
rect -3004 -199 -2900 199
rect -224 148 -204 5172
rect -140 148 -120 5172
rect 2608 5121 2712 5519
rect 5388 5468 5408 10492
rect 5472 5468 5492 10492
rect 5388 5172 5492 5468
rect 199 5120 5121 5121
rect 199 200 200 5120
rect 5120 200 5121 5120
rect 199 199 5121 200
rect -224 -148 -120 148
rect -5413 -200 -491 -199
rect -5413 -5120 -5412 -200
rect -492 -5120 -491 -200
rect -5413 -5121 -491 -5120
rect -3004 -5519 -2900 -5121
rect -224 -5172 -204 -148
rect -140 -5172 -120 -148
rect 2608 -199 2712 199
rect 5388 148 5408 5172
rect 5472 148 5492 5172
rect 5388 -148 5492 148
rect 199 -200 5121 -199
rect 199 -5120 200 -200
rect 5120 -5120 5121 -200
rect 199 -5121 5121 -5120
rect -224 -5468 -120 -5172
rect -5413 -5520 -491 -5519
rect -5413 -10440 -5412 -5520
rect -492 -10440 -491 -5520
rect -5413 -10441 -491 -10440
rect -3004 -10640 -2900 -10441
rect -224 -10492 -204 -5468
rect -140 -10492 -120 -5468
rect 2608 -5519 2712 -5121
rect 5388 -5172 5408 -148
rect 5472 -5172 5492 -148
rect 5388 -5468 5492 -5172
rect 199 -5520 5121 -5519
rect 199 -10440 200 -5520
rect 5120 -10440 5121 -5520
rect 199 -10441 5121 -10440
rect -224 -10640 -120 -10492
rect 2608 -10640 2712 -10441
rect 5388 -10492 5408 -5468
rect 5472 -10492 5492 -5468
rect 5388 -10640 5492 -10492
<< properties >>
string FIXED_BBOX 120 5440 5200 10520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 25.0 val 1.269k carea 2.00 cperi 0.19 class capacitor nx 2 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
