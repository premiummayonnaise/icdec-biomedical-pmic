* SPICE3 file created from two-stage-miller.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_V6JW4R a_n267_n536# a_29_n562# a_209_n536# a_n29_n536#
+ w_n467_n762# a_n209_n562# VSUBS
X0 a_n29_n536# a_n209_n562# a_n267_n536# w_n467_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.9
X1 a_209_n536# a_29_n562# a_n29_n536# w_n467_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.9
C0 a_n209_n562# w_n467_n762# 0.19926f
C1 a_n29_n536# a_209_n536# 0.29682f
C2 a_29_n562# a_209_n536# 0.10455f
C3 a_n267_n536# a_n29_n536# 0.29682f
C4 w_n467_n762# a_209_n536# 0.08941f
C5 a_29_n562# a_n29_n536# 0.10455f
C6 a_n267_n536# a_n209_n562# 0.10455f
C7 a_n209_n562# a_n29_n536# 0.10455f
C8 a_n267_n536# w_n467_n762# 0.08941f
C9 w_n467_n762# a_n29_n536# 0.01994f
C10 a_n209_n562# a_29_n562# 0.0619f
C11 a_29_n562# w_n467_n762# 0.19926f
C12 a_209_n536# VSUBS 0.41875f
C13 a_n29_n536# VSUBS 0.13822f
C14 a_n267_n536# VSUBS 0.41875f
C15 a_29_n562# VSUBS 0.23237f
C16 a_n209_n562# VSUBS 0.23237f
C17 w_n467_n762# VSUBS 4.49444f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_RFPNS8 a_587_n964# a_1203_n964# a_337_n1061#
+ a_n279_n1061# a_953_n1061# a_n895_n1061# a_n1203_n1061# a_n337_n964# a_n953_n964#
+ a_29_n1061# a_279_n964# a_895_n964# w_n1461_n1262# a_n1261_n964# a_645_n1061# a_n587_n1061#
+ a_n645_n964# a_n29_n964# VSUBS
X0 a_895_n964# a_645_n1061# a_587_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X1 a_n645_n964# a_n895_n1061# a_n953_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X2 a_n29_n964# a_n279_n1061# a_n337_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X3 a_n953_n964# a_n1203_n1061# a_n1261_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1.25
X4 a_1203_n964# a_953_n1061# a_895_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1.25
X5 a_587_n964# a_337_n1061# a_279_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X6 a_n337_n964# a_n587_n1061# a_n645_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X7 a_279_n964# a_29_n1061# a_n29_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
C0 a_1203_n964# a_895_n964# 0.45807f
C1 a_645_n1061# a_895_n964# 0.25181f
C2 a_n645_n964# a_n587_n1061# 0.25181f
C3 a_n645_n964# a_n337_n964# 0.45807f
C4 a_n1203_n1061# w_n1461_n1262# 0.2506f
C5 a_n279_n1061# a_29_n1061# 0.0619f
C6 a_n953_n964# a_n895_n1061# 0.25181f
C7 a_587_n964# a_279_n964# 0.45807f
C8 a_n29_n964# w_n1461_n1262# 0.01993f
C9 a_279_n964# a_29_n1061# 0.25181f
C10 a_n953_n964# a_n1203_n1061# 0.25181f
C11 a_n645_n964# a_n895_n1061# 0.25181f
C12 w_n1461_n1262# a_953_n1061# 0.2506f
C13 a_337_n1061# a_279_n964# 0.25181f
C14 a_n953_n964# w_n1461_n1262# 0.01993f
C15 a_n587_n1061# a_n337_n964# 0.25181f
C16 a_587_n964# w_n1461_n1262# 0.01993f
C17 a_n29_n964# a_29_n1061# 0.25181f
C18 a_n1203_n1061# a_n1261_n964# 0.25181f
C19 a_n587_n1061# a_n279_n1061# 0.0619f
C20 w_n1461_n1262# a_29_n1061# 0.23077f
C21 a_n279_n1061# a_n337_n964# 0.25181f
C22 a_n645_n964# w_n1461_n1262# 0.01993f
C23 w_n1461_n1262# a_n1261_n964# 0.15606f
C24 a_337_n1061# w_n1461_n1262# 0.23077f
C25 a_n587_n1061# a_n895_n1061# 0.0619f
C26 w_n1461_n1262# a_1203_n964# 0.15606f
C27 w_n1461_n1262# a_645_n1061# 0.23077f
C28 a_n645_n964# a_n953_n964# 0.45807f
C29 w_n1461_n1262# a_895_n964# 0.01993f
C30 a_n953_n964# a_n1261_n964# 0.45807f
C31 a_587_n964# a_337_n1061# 0.25181f
C32 a_953_n1061# a_1203_n964# 0.25181f
C33 a_953_n1061# a_645_n1061# 0.0619f
C34 a_953_n1061# a_895_n964# 0.25181f
C35 a_n29_n964# a_n337_n964# 0.45807f
C36 a_n587_n1061# w_n1461_n1262# 0.23077f
C37 a_337_n1061# a_29_n1061# 0.0619f
C38 a_587_n964# a_645_n1061# 0.25181f
C39 w_n1461_n1262# a_n337_n964# 0.01993f
C40 a_587_n964# a_895_n964# 0.45807f
C41 a_n29_n964# a_n279_n1061# 0.25181f
C42 w_n1461_n1262# a_n279_n1061# 0.23077f
C43 a_n1203_n1061# a_n895_n1061# 0.0619f
C44 a_n29_n964# a_279_n964# 0.45807f
C45 a_337_n1061# a_645_n1061# 0.0619f
C46 a_279_n964# w_n1461_n1262# 0.01993f
C47 a_n895_n1061# w_n1461_n1262# 0.23077f
C48 a_1203_n964# VSUBS 0.85861f
C49 a_895_n964# VSUBS 0.33133f
C50 a_587_n964# VSUBS 0.33133f
C51 a_279_n964# VSUBS 0.33133f
C52 a_n29_n964# VSUBS 0.33133f
C53 a_n337_n964# VSUBS 0.33133f
C54 a_n645_n964# VSUBS 0.33133f
C55 a_n953_n964# VSUBS 0.33133f
C56 a_n1261_n964# VSUBS 0.85861f
C57 a_953_n1061# VSUBS 0.32776f
C58 a_645_n1061# VSUBS 0.31082f
C59 a_337_n1061# VSUBS 0.31082f
C60 a_29_n1061# VSUBS 0.31082f
C61 a_n279_n1061# VSUBS 0.31082f
C62 a_n587_n1061# VSUBS 0.31082f
C63 a_n895_n1061# VSUBS 0.31082f
C64 a_n1203_n1061# VSUBS 0.32776f
C65 w_n1461_n1262# VSUBS 23.138f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_S5VYLR a_n337_n904# a_n587_n968# a_n953_n904#
+ a_645_n968# a_29_n968# a_1261_n968# a_1569_n968# a_n2185_n904# a_2435_n904# a_n2435_n968#
+ a_279_n904# a_895_n904# a_1511_n904# a_n1261_n904# a_n1569_n904# a_n1511_n968# a_1819_n904#
+ a_n1819_n968# a_n279_n968# a_n29_n904# a_n645_n904# a_n895_n968# a_337_n968# a_953_n968#
+ w_n2693_n1202# a_2127_n904# a_1877_n968# a_n2493_n904# a_n2127_n968# a_587_n904#
+ a_1203_n904# a_n1203_n968# a_n1877_n904# a_2185_n968# VSUBS
X0 a_n1877_n904# a_n2127_n968# a_n2185_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X1 a_895_n904# a_645_n968# a_587_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X2 a_n1569_n904# a_n1819_n968# a_n1877_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X3 a_n645_n904# a_n895_n968# a_n953_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X4 a_1819_n904# a_1569_n968# a_1511_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X5 a_n29_n904# a_n279_n968# a_n337_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X6 a_n2185_n904# a_n2435_n968# a_n2493_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=2.726 ps=19.38 w=9.4 l=1.25
X7 a_n953_n904# a_n1203_n968# a_n1261_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X8 a_1203_n904# a_953_n968# a_895_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X9 a_2435_n904# a_2185_n968# a_2127_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=2.726 pd=19.38 as=1.363 ps=9.69 w=9.4 l=1.25
X10 a_587_n904# a_337_n968# a_279_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X11 a_2127_n904# a_1877_n968# a_1819_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X12 a_n337_n904# a_n587_n968# a_n645_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X13 a_279_n904# a_29_n968# a_n29_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X14 a_n1261_n904# a_n1511_n968# a_n1569_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X15 a_1511_n904# a_1261_n968# a_1203_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
C0 a_n1261_n904# a_n1511_n968# 0.23705f
C1 a_953_n968# w_n2693_n1202# 0.21732f
C2 a_n1203_n968# a_n1511_n968# 0.04019f
C3 a_n1569_n904# a_n1877_n904# 0.43064f
C4 a_n1877_n904# a_n2185_n904# 0.43064f
C5 a_n29_n904# a_n279_n968# 0.23705f
C6 a_n279_n968# a_n337_n904# 0.23705f
C7 a_n279_n968# a_n587_n968# 0.04019f
C8 a_n1877_n904# w_n2693_n1202# 0.01993f
C9 a_645_n968# a_953_n968# 0.04019f
C10 a_29_n968# a_279_n904# 0.23705f
C11 a_n1261_n904# a_n1569_n904# 0.43064f
C12 a_1261_n968# w_n2693_n1202# 0.21732f
C13 a_895_n904# a_953_n968# 0.23705f
C14 a_n1261_n904# a_n953_n904# 0.43064f
C15 a_n1819_n968# a_n2127_n968# 0.04019f
C16 a_2435_n904# w_n2693_n1202# 0.14807f
C17 a_n1203_n968# a_n953_n904# 0.23705f
C18 a_n1569_n904# a_n1511_n968# 0.23705f
C19 a_n1261_n904# w_n2693_n1202# 0.01993f
C20 a_n29_n904# a_n337_n904# 0.43064f
C21 w_n2693_n1202# a_n1203_n968# 0.21732f
C22 a_n587_n968# a_n337_n904# 0.23705f
C23 a_1511_n904# w_n2693_n1202# 0.01993f
C24 w_n2693_n1202# a_n1511_n968# 0.21732f
C25 a_1569_n968# a_1819_n904# 0.23705f
C26 a_2435_n904# a_2185_n968# 0.23705f
C27 a_n1877_n904# a_n2127_n968# 0.23705f
C28 a_n645_n904# a_n337_n904# 0.43064f
C29 a_n29_n904# a_279_n904# 0.43064f
C30 a_n645_n904# a_n587_n968# 0.23705f
C31 w_n2693_n1202# a_n2185_n904# 0.01993f
C32 a_n1569_n904# w_n2693_n1202# 0.01993f
C33 w_n2693_n1202# a_n953_n904# 0.01993f
C34 a_n895_n968# a_n587_n968# 0.04019f
C35 a_337_n968# w_n2693_n1202# 0.21732f
C36 a_2127_n904# a_1819_n904# 0.43064f
C37 a_337_n968# a_587_n904# 0.23705f
C38 a_1877_n968# w_n2693_n1202# 0.21732f
C39 a_587_n904# w_n2693_n1202# 0.01993f
C40 a_337_n968# a_645_n968# 0.04019f
C41 a_645_n968# w_n2693_n1202# 0.21732f
C42 a_n2493_n904# a_n2185_n904# 0.43064f
C43 a_n895_n968# a_n645_n904# 0.23705f
C44 a_1261_n968# a_1569_n968# 0.04019f
C45 a_587_n904# a_645_n968# 0.23705f
C46 a_895_n904# w_n2693_n1202# 0.01993f
C47 a_2185_n968# w_n2693_n1202# 0.2317f
C48 a_953_n968# a_1203_n904# 0.23705f
C49 a_n2493_n904# w_n2693_n1202# 0.14807f
C50 a_n2127_n968# a_n2185_n904# 0.23705f
C51 a_2185_n968# a_1877_n968# 0.04019f
C52 a_587_n904# a_895_n904# 0.43064f
C53 a_1511_n904# a_1569_n968# 0.23705f
C54 a_337_n968# a_29_n968# 0.04019f
C55 a_895_n904# a_645_n968# 0.23705f
C56 a_n2127_n968# w_n2693_n1202# 0.21732f
C57 a_29_n968# w_n2693_n1202# 0.21732f
C58 a_2127_n904# a_2435_n904# 0.43064f
C59 a_1261_n968# a_1203_n904# 0.23705f
C60 a_n1819_n968# a_n1877_n904# 0.23705f
C61 a_n279_n968# w_n2693_n1202# 0.21732f
C62 a_n2435_n968# a_n2185_n904# 0.23705f
C63 a_1511_n904# a_1203_n904# 0.43064f
C64 a_1569_n968# w_n2693_n1202# 0.21732f
C65 a_n2435_n968# w_n2693_n1202# 0.2317f
C66 a_1569_n968# a_1877_n968# 0.04019f
C67 a_n895_n968# a_n1203_n968# 0.04019f
C68 a_1511_n904# a_1819_n904# 0.43064f
C69 a_1261_n968# a_953_n968# 0.04019f
C70 a_n29_n904# w_n2693_n1202# 0.01993f
C71 a_n337_n904# w_n2693_n1202# 0.01993f
C72 a_n587_n968# w_n2693_n1202# 0.21732f
C73 a_n1819_n968# a_n1511_n968# 0.04019f
C74 a_2127_n904# w_n2693_n1202# 0.01993f
C75 a_1203_n904# w_n2693_n1202# 0.01993f
C76 a_2127_n904# a_1877_n968# 0.23705f
C77 a_n279_n968# a_29_n968# 0.04019f
C78 a_n645_n904# a_n953_n904# 0.43064f
C79 a_n2435_n968# a_n2493_n904# 0.23705f
C80 a_337_n968# a_279_n904# 0.23705f
C81 a_n645_n904# w_n2693_n1202# 0.01993f
C82 a_n1569_n904# a_n1819_n968# 0.23705f
C83 a_279_n904# w_n2693_n1202# 0.01993f
C84 a_n895_n968# a_n953_n904# 0.23705f
C85 w_n2693_n1202# a_1819_n904# 0.01993f
C86 a_n2435_n968# a_n2127_n968# 0.04019f
C87 a_n895_n968# w_n2693_n1202# 0.21732f
C88 a_587_n904# a_279_n904# 0.43064f
C89 a_1877_n968# a_1819_n904# 0.23705f
C90 a_n1819_n968# w_n2693_n1202# 0.21732f
C91 a_2127_n904# a_2185_n968# 0.23705f
C92 a_1511_n904# a_1261_n968# 0.23705f
C93 a_895_n904# a_1203_n904# 0.43064f
C94 a_n29_n904# a_29_n968# 0.23705f
C95 a_n1261_n904# a_n1203_n968# 0.23705f
C96 a_2435_n904# VSUBS 0.80781f
C97 a_2127_n904# VSUBS 0.31212f
C98 a_1819_n904# VSUBS 0.31212f
C99 a_1511_n904# VSUBS 0.31212f
C100 a_1203_n904# VSUBS 0.31212f
C101 a_895_n904# VSUBS 0.31212f
C102 a_587_n904# VSUBS 0.31212f
C103 a_279_n904# VSUBS 0.31212f
C104 a_n29_n904# VSUBS 0.31212f
C105 a_n337_n904# VSUBS 0.31212f
C106 a_n645_n904# VSUBS 0.31212f
C107 a_n953_n904# VSUBS 0.31212f
C108 a_n1261_n904# VSUBS 0.31212f
C109 a_n1569_n904# VSUBS 0.31212f
C110 a_n1877_n904# VSUBS 0.31212f
C111 a_n2185_n904# VSUBS 0.31212f
C112 a_n2493_n904# VSUBS 0.80781f
C113 a_2185_n968# VSUBS 0.22385f
C114 a_1877_n968# VSUBS 0.20885f
C115 a_1569_n968# VSUBS 0.20885f
C116 a_1261_n968# VSUBS 0.20885f
C117 a_953_n968# VSUBS 0.20885f
C118 a_645_n968# VSUBS 0.20885f
C119 a_337_n968# VSUBS 0.20885f
C120 a_29_n968# VSUBS 0.20885f
C121 a_n279_n968# VSUBS 0.20885f
C122 a_n587_n968# VSUBS 0.20885f
C123 a_n895_n968# VSUBS 0.20885f
C124 a_n1203_n968# VSUBS 0.20885f
C125 a_n1511_n968# VSUBS 0.20885f
C126 a_n1819_n968# VSUBS 0.20885f
C127 a_n2127_n968# VSUBS 0.20885f
C128 a_n2435_n968# VSUBS 0.22385f
C129 w_n2693_n1202# VSUBS 40.8176f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DC2CKB a_n29_n440# a_29_n495# a_n187_n440# a_n129_n495#
+ a_187_n495# a_n287_n495# a_n345_n440# a_129_n440# a_287_n440# a_n479_n662#
X0 a_n187_n440# a_n287_n495# a_n345_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=1.3659 ps=10 w=4.71 l=0.5
X1 a_287_n440# a_187_n495# a_129_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3659 pd=10 as=0.68295 ps=5 w=4.71 l=0.5
X2 a_129_n440# a_29_n495# a_n29_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X3 a_n29_n440# a_n129_n495# a_n187_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
C0 a_n187_n440# a_n287_n495# 0.06224f
C1 a_287_n440# a_129_n440# 0.42026f
C2 a_n29_n440# a_n129_n495# 0.06224f
C3 a_n345_n440# a_n187_n440# 0.42026f
C4 a_129_n440# a_n29_n440# 0.42026f
C5 a_n129_n495# a_n187_n440# 0.06224f
C6 a_187_n495# a_29_n495# 0.05012f
C7 a_n29_n440# a_n187_n440# 0.42026f
C8 a_n345_n440# a_n287_n495# 0.06224f
C9 a_287_n440# a_187_n495# 0.06224f
C10 a_n129_n495# a_n287_n495# 0.05012f
C11 a_n129_n495# a_29_n495# 0.05012f
C12 a_129_n440# a_187_n495# 0.06224f
C13 a_129_n440# a_29_n495# 0.06224f
C14 a_n29_n440# a_29_n495# 0.06224f
C15 a_287_n440# a_n479_n662# 0.45374f
C16 a_129_n440# a_n479_n662# 0.1076f
C17 a_n29_n440# a_n479_n662# 0.1076f
C18 a_n187_n440# a_n479_n662# 0.1076f
C19 a_n345_n440# a_n479_n662# 0.49789f
C20 a_187_n495# a_n479_n662# 0.23558f
C21 a_29_n495# a_n479_n662# 0.20272f
C22 a_n129_n495# a_n479_n662# 0.20272f
C23 a_n287_n495# a_n479_n662# 0.23657f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2899RY a_n953_n781# a_2185_n807# a_n587_n807#
+ a_645_n807# a_29_n807# a_2435_n781# a_n2185_n781# a_1261_n807# a_1569_n807# a_279_n781#
+ a_895_n781# a_n2435_n807# a_n1261_n781# a_1511_n781# a_1819_n781# a_n1569_n781#
+ a_n29_n781# a_n645_n781# a_n1511_n807# a_n279_n807# a_n1819_n807# a_n895_n807# a_337_n807#
+ a_953_n807# a_2127_n781# a_n2493_n781# a_587_n781# a_1877_n807# a_n2627_n941# a_n2127_n807#
+ a_1203_n781# a_n1877_n781# a_n337_n781# a_n1203_n807#
X0 a_1511_n781# a_1261_n807# a_1203_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X1 a_n1261_n781# a_n1511_n807# a_n1569_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X2 a_n1877_n781# a_n2127_n807# a_n2185_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X3 a_895_n781# a_645_n807# a_587_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X4 a_n1569_n781# a_n1819_n807# a_n1877_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X5 a_n645_n781# a_n895_n807# a_n953_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X6 a_1819_n781# a_1569_n807# a_1511_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X7 a_n29_n781# a_n279_n807# a_n337_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X8 a_n953_n781# a_n1203_n807# a_n1261_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X9 a_2435_n781# a_2185_n807# a_2127_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=1.25
X10 a_n2185_n781# a_n2435_n807# a_n2493_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=1.25
X11 a_1203_n781# a_953_n807# a_895_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X12 a_587_n781# a_337_n807# a_279_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X13 a_2127_n781# a_1877_n807# a_1819_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X14 a_n337_n781# a_n587_n807# a_n645_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X15 a_279_n781# a_29_n807# a_n29_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
C0 a_2127_n781# a_1819_n781# 0.34377f
C1 a_587_n781# a_895_n781# 0.34377f
C2 a_n1569_n781# a_n1511_n807# 0.19032f
C3 a_n1569_n781# a_n1877_n781# 0.34377f
C4 a_587_n781# a_645_n807# 0.19032f
C5 a_587_n781# a_279_n781# 0.34377f
C6 a_1511_n781# a_1819_n781# 0.34377f
C7 a_n2435_n807# a_n2127_n807# 0.02909f
C8 a_279_n781# a_29_n807# 0.19032f
C9 a_279_n781# a_n29_n781# 0.34377f
C10 a_n1203_n807# a_n1511_n807# 0.02909f
C11 a_n1569_n781# a_n1819_n807# 0.19032f
C12 a_1877_n807# a_2185_n807# 0.02909f
C13 a_n1819_n807# a_n1511_n807# 0.02909f
C14 a_n1203_n807# a_n895_n807# 0.02909f
C15 a_n1819_n807# a_n1877_n781# 0.19032f
C16 a_2127_n781# a_2185_n807# 0.19032f
C17 a_n2185_n781# a_n1877_n781# 0.34377f
C18 a_1877_n807# a_1569_n807# 0.02909f
C19 a_645_n807# a_895_n781# 0.19032f
C20 a_587_n781# a_337_n807# 0.19032f
C21 a_n645_n781# a_n337_n781# 0.34377f
C22 a_1261_n807# a_1569_n807# 0.02909f
C23 a_29_n807# a_337_n807# 0.02909f
C24 a_n645_n781# a_n895_n807# 0.19032f
C25 a_n337_n781# a_n279_n807# 0.19032f
C26 a_953_n807# a_895_n781# 0.19032f
C27 a_1511_n781# a_1569_n807# 0.19032f
C28 a_953_n807# a_645_n807# 0.02909f
C29 a_n587_n807# a_n337_n781# 0.19032f
C30 a_n953_n781# a_n1261_n781# 0.34377f
C31 a_2127_n781# a_1877_n807# 0.19032f
C32 a_n337_n781# a_n29_n781# 0.34377f
C33 a_n587_n807# a_n895_n807# 0.02909f
C34 a_1261_n807# a_953_n807# 0.02909f
C35 a_n645_n781# a_n587_n807# 0.19032f
C36 a_2435_n781# a_2185_n807# 0.19032f
C37 a_1511_n781# a_1261_n807# 0.19032f
C38 a_n2435_n807# a_n2185_n781# 0.19032f
C39 a_n587_n807# a_n279_n807# 0.02909f
C40 a_1203_n781# a_895_n781# 0.34377f
C41 a_337_n807# a_645_n807# 0.02909f
C42 a_n2185_n781# a_n2493_n781# 0.34377f
C43 a_279_n781# a_337_n807# 0.19032f
C44 a_n953_n781# a_n1203_n807# 0.19032f
C45 a_n1877_n781# a_n2127_n807# 0.19032f
C46 a_29_n807# a_n279_n807# 0.02909f
C47 a_n29_n781# a_n279_n807# 0.19032f
C48 a_1203_n781# a_953_n807# 0.19032f
C49 a_n1569_n781# a_n1261_n781# 0.34377f
C50 a_n1819_n807# a_n2127_n807# 0.02909f
C51 a_1203_n781# a_1261_n807# 0.19032f
C52 a_1819_n781# a_1569_n807# 0.19032f
C53 a_n953_n781# a_n895_n807# 0.19032f
C54 a_n29_n781# a_29_n807# 0.19032f
C55 a_n2185_n781# a_n2127_n807# 0.19032f
C56 a_1203_n781# a_1511_n781# 0.34377f
C57 a_n953_n781# a_n645_n781# 0.34377f
C58 a_2127_n781# a_2435_n781# 0.34377f
C59 a_n1203_n807# a_n1261_n781# 0.19032f
C60 a_n1261_n781# a_n1511_n807# 0.19032f
C61 a_n2435_n807# a_n2493_n781# 0.19032f
C62 a_1877_n807# a_1819_n781# 0.19032f
C63 a_2435_n781# a_n2627_n941# 0.76245f
C64 a_2127_n781# a_n2627_n941# 0.27094f
C65 a_1819_n781# a_n2627_n941# 0.27094f
C66 a_1511_n781# a_n2627_n941# 0.27094f
C67 a_1203_n781# a_n2627_n941# 0.27094f
C68 a_895_n781# a_n2627_n941# 0.27094f
C69 a_587_n781# a_n2627_n941# 0.27094f
C70 a_279_n781# a_n2627_n941# 0.27094f
C71 a_n29_n781# a_n2627_n941# 0.27094f
C72 a_n337_n781# a_n2627_n941# 0.27094f
C73 a_n645_n781# a_n2627_n941# 0.27094f
C74 a_n953_n781# a_n2627_n941# 0.27094f
C75 a_n1261_n781# a_n2627_n941# 0.27094f
C76 a_n1569_n781# a_n2627_n941# 0.27094f
C77 a_n1877_n781# a_n2627_n941# 0.27094f
C78 a_n2185_n781# a_n2627_n941# 0.27094f
C79 a_n2493_n781# a_n2627_n941# 0.76245f
C80 a_2185_n807# a_n2627_n941# 0.41942f
C81 a_1877_n807# a_n2627_n941# 0.39834f
C82 a_1569_n807# a_n2627_n941# 0.39834f
C83 a_1261_n807# a_n2627_n941# 0.39834f
C84 a_953_n807# a_n2627_n941# 0.39834f
C85 a_645_n807# a_n2627_n941# 0.39834f
C86 a_337_n807# a_n2627_n941# 0.39834f
C87 a_29_n807# a_n2627_n941# 0.39834f
C88 a_n279_n807# a_n2627_n941# 0.39834f
C89 a_n587_n807# a_n2627_n941# 0.39834f
C90 a_n895_n807# a_n2627_n941# 0.39834f
C91 a_n1203_n807# a_n2627_n941# 0.39834f
C92 a_n1511_n807# a_n2627_n941# 0.39834f
C93 a_n1819_n807# a_n2627_n941# 0.39834f
C94 a_n2127_n807# a_n2627_n941# 0.39834f
C95 a_n2435_n807# a_n2627_n941# 0.41942f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_A8KA9K a_n29_n440# a_29_n495# a_n187_n440# a_n129_n495#
+ a_187_n495# a_n287_n495# a_n345_n440# a_129_n440# a_287_n440# a_n479_n662#
X0 a_n187_n440# a_n287_n495# a_n345_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=1.3659 ps=10 w=4.71 l=0.5
X1 a_287_n440# a_187_n495# a_129_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3659 pd=10 as=0.68295 ps=5 w=4.71 l=0.5
X2 a_129_n440# a_29_n495# a_n29_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X3 a_n29_n440# a_n129_n495# a_n187_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
C0 a_187_n495# a_29_n495# 0.03586f
C1 a_n129_n495# a_29_n495# 0.03586f
C2 a_n287_n495# a_n345_n440# 0.06224f
C3 a_129_n440# a_29_n495# 0.06224f
C4 a_n29_n440# a_n129_n495# 0.06224f
C5 a_n29_n440# a_129_n440# 0.42026f
C6 a_n187_n440# a_n129_n495# 0.06224f
C7 a_n187_n440# a_n287_n495# 0.06224f
C8 a_n29_n440# a_29_n495# 0.06224f
C9 a_n187_n440# a_n345_n440# 0.42026f
C10 a_287_n440# a_187_n495# 0.06224f
C11 a_129_n440# a_187_n495# 0.06224f
C12 a_129_n440# a_287_n440# 0.42026f
C13 a_n29_n440# a_n187_n440# 0.42026f
C14 a_n287_n495# a_n129_n495# 0.03586f
C15 a_287_n440# a_n479_n662# 0.49789f
C16 a_129_n440# a_n479_n662# 0.1076f
C17 a_n29_n440# a_n479_n662# 0.1076f
C18 a_n187_n440# a_n479_n662# 0.1076f
C19 a_n345_n440# a_n479_n662# 0.45374f
C20 a_187_n495# a_n479_n662# 0.21175f
C21 a_29_n495# a_n479_n662# 0.18614f
C22 a_n129_n495# a_n479_n662# 0.18614f
C23 a_n287_n495# a_n479_n662# 0.21095f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_N5GNFR a_n587_n807# a_29_n807# a_279_n781# a_n29_n781#
+ a_n645_n781# a_n779_n941# a_n279_n807# a_337_n807# a_587_n781# a_n337_n781#
X0 a_n29_n781# a_n279_n807# a_n337_n781# a_n779_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X1 a_587_n781# a_337_n807# a_279_n781# a_n779_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=1.25
X2 a_n337_n781# a_n587_n807# a_n645_n781# a_n779_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=1.25
X3 a_279_n781# a_29_n807# a_n29_n781# a_n779_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
C0 a_29_n807# a_279_n781# 0.19032f
C1 a_n337_n781# a_n645_n781# 0.34377f
C2 a_n645_n781# a_n587_n807# 0.19032f
C3 a_29_n807# a_n29_n781# 0.19032f
C4 a_n279_n807# a_n337_n781# 0.19032f
C5 a_29_n807# a_337_n807# 0.05942f
C6 a_n279_n807# a_n587_n807# 0.05942f
C7 a_n337_n781# a_n587_n807# 0.19032f
C8 a_587_n781# a_279_n781# 0.34377f
C9 a_n279_n807# a_n29_n781# 0.19032f
C10 a_n337_n781# a_n29_n781# 0.34377f
C11 a_n29_n781# a_279_n781# 0.34377f
C12 a_n279_n807# a_29_n807# 0.05942f
C13 a_337_n807# a_279_n781# 0.19032f
C14 a_337_n807# a_587_n781# 0.19032f
C15 a_587_n781# a_n779_n941# 0.76245f
C16 a_279_n781# a_n779_n941# 0.27094f
C17 a_n29_n781# a_n779_n941# 0.27094f
C18 a_n337_n781# a_n779_n941# 0.27094f
C19 a_n645_n781# a_n779_n941# 0.76245f
C20 a_337_n807# a_n779_n941# 0.56775f
C21 a_29_n807# a_n779_n941# 0.53283f
C22 a_n279_n807# a_n779_n941# 0.53283f
C23 a_n587_n807# a_n779_n941# 0.56775f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_X6KG9Z a_n345_n502# a_129_n502# a_29_n528# a_n129_n528#
+ a_287_n502# a_187_n528# a_n287_n528# a_n29_n502# a_n479_n662# a_n187_n502#
X0 a_287_n502# a_187_n528# a_129_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3659 pd=10 as=0.68295 ps=5 w=4.71 l=0.5
X1 a_129_n502# a_29_n528# a_n29_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X2 a_n29_n502# a_n129_n528# a_n187_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X3 a_n187_n502# a_n287_n528# a_n345_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=1.3659 ps=10 w=4.71 l=0.5
C0 a_n187_n502# a_n287_n528# 0.06224f
C1 a_287_n502# a_129_n502# 0.42026f
C2 a_29_n528# a_187_n528# 0.05012f
C3 a_n287_n528# a_n345_n502# 0.06224f
C4 a_n29_n502# a_n129_n528# 0.06224f
C5 a_29_n528# a_n129_n528# 0.05012f
C6 a_n287_n528# a_n129_n528# 0.05012f
C7 a_29_n528# a_n29_n502# 0.06224f
C8 a_287_n502# a_187_n528# 0.06224f
C9 a_129_n502# a_187_n528# 0.06224f
C10 a_n187_n502# a_n345_n502# 0.42026f
C11 a_129_n502# a_n29_n502# 0.42026f
C12 a_29_n528# a_129_n502# 0.06224f
C13 a_n187_n502# a_n129_n528# 0.06224f
C14 a_n187_n502# a_n29_n502# 0.42026f
C15 a_287_n502# a_n479_n662# 0.49789f
C16 a_129_n502# a_n479_n662# 0.1076f
C17 a_n29_n502# a_n479_n662# 0.1076f
C18 a_n187_n502# a_n479_n662# 0.1076f
C19 a_n345_n502# a_n479_n662# 0.45374f
C20 a_187_n528# a_n479_n662# 0.23657f
C21 a_29_n528# a_n479_n662# 0.20272f
C22 a_n129_n528# a_n479_n662# 0.20272f
C23 a_n287_n528# a_n479_n662# 0.23558f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_R7S84X m3_n2686_n21160# c1_n2646_n21120# VSUBS
X0 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X1 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X2 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X3 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X4 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X5 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X6 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X7 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
C0 m3_n2686_n21160# c1_n2646_n21120# 0.44473p
C1 c1_n2646_n21120# VSUBS 11.1251f
C2 m3_n2686_n21160# VSUBS 97.539f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PBQQNH a_n345_n502# a_129_n502# a_29_n528# a_n129_n528#
+ a_287_n502# a_187_n528# a_n287_n528# a_n29_n502# a_n479_n662# a_n187_n502#
X0 a_287_n502# a_187_n528# a_129_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3659 pd=10 as=0.68295 ps=5 w=4.71 l=0.5
X1 a_129_n502# a_29_n528# a_n29_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X2 a_n29_n502# a_n129_n528# a_n187_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X3 a_n187_n502# a_n287_n528# a_n345_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=1.3659 ps=10 w=4.71 l=0.5
C0 a_n29_n502# a_129_n502# 0.42026f
C1 a_n287_n528# a_n187_n502# 0.06224f
C2 a_129_n502# a_187_n528# 0.06224f
C3 a_29_n528# a_129_n502# 0.06224f
C4 a_n29_n502# a_n187_n502# 0.42026f
C5 a_n187_n502# a_n129_n528# 0.06224f
C6 a_n287_n528# a_n129_n528# 0.03586f
C7 a_n29_n502# a_n129_n528# 0.06224f
C8 a_n345_n502# a_n187_n502# 0.42026f
C9 a_187_n528# a_287_n502# 0.06224f
C10 a_n287_n528# a_n345_n502# 0.06224f
C11 a_29_n528# a_n29_n502# 0.06224f
C12 a_29_n528# a_n129_n528# 0.03586f
C13 a_29_n528# a_187_n528# 0.03586f
C14 a_129_n502# a_287_n502# 0.42026f
C15 a_287_n502# a_n479_n662# 0.45374f
C16 a_129_n502# a_n479_n662# 0.1076f
C17 a_n29_n502# a_n479_n662# 0.1076f
C18 a_n187_n502# a_n479_n662# 0.1076f
C19 a_n345_n502# a_n479_n662# 0.49789f
C20 a_187_n528# a_n479_n662# 0.21095f
C21 a_29_n528# a_n479_n662# 0.18614f
C22 a_n129_n528# a_n479_n662# 0.18614f
C23 a_n287_n528# a_n479_n662# 0.21175f
.ends

.subckt two-stage-miller VDD OUT VP VN IBIAS VSS
Xsky130_fd_pr__pfet_g5v0d10v5_V6JW4R_1 OUT VSS OUT m1_n2200_3200# VDD VSS VSS sky130_fd_pr__pfet_g5v0d10v5_V6JW4R
Xsky130_fd_pr__pfet_g5v0d10v5_RFPNS8_0 OUT OUT m1_n1120_1120# m1_n1120_1120# m1_n1120_1120#
+ m1_n1120_1120# m1_n1120_1120# VDD VDD m1_n1120_1120# VDD VDD VDD OUT m1_n1120_1120#
+ m1_n1120_1120# OUT OUT VSS sky130_fd_pr__pfet_g5v0d10v5_RFPNS8
XXM2 VDD m1_2160_1440# VDD m1_2160_1440# m1_2160_1440# m1_2160_1440# m1_2160_1440#
+ VDD m1_2160_1440# m1_2160_1440# VDD VDD VDD m1_2160_1440# VDD m1_2160_1440# m1_n1120_1120#
+ m1_2160_1440# m1_2160_1440# m1_2160_1440# m1_n1120_1120# m1_2160_1440# m1_2160_1440#
+ m1_2160_1440# VDD VDD m1_2160_1440# m1_2160_1440# m1_2160_1440# m1_n1120_1120# m1_2160_1440#
+ m1_2160_1440# m1_n1120_1120# m1_2160_1440# VSS sky130_fd_pr__pfet_g5v0d10v5_S5VYLR
XXM3 m1_2160_1440# VP m1_2740_n3440# VP VP VP m1_2160_1440# m1_2740_n3440# m1_2160_1440#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_DC2CKB
XXM5 VSS IBIAS IBIAS IBIAS IBIAS IBIAS VSS IBIAS IBIAS VSS VSS IBIAS IBIAS VSS m1_2740_n3440#
+ VSS IBIAS m1_2740_n3440# IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS VSS IBIAS m1_2740_n3440#
+ IBIAS VSS IBIAS IBIAS m1_2740_n3440# VSS IBIAS sky130_fd_pr__nfet_g5v0d10v5_2899RY
Xsky130_fd_pr__nfet_g5v0d10v5_A8KA9K_0 m1_n1120_1120# VN m1_2740_n3440# VN VN VN m1_n1120_1120#
+ m1_2740_n3440# m1_n1120_1120# VSS sky130_fd_pr__nfet_g5v0d10v5_A8KA9K
XXM7 OUT OUT m1_n1120_1120# m1_n1120_1120# m1_n1120_1120# m1_n1120_1120# m1_n1120_1120#
+ VDD VDD m1_n1120_1120# VDD VDD VDD OUT m1_n1120_1120# m1_n1120_1120# OUT OUT VSS
+ sky130_fd_pr__pfet_g5v0d10v5_RFPNS8
XXM8 IBIAS IBIAS VSS OUT OUT VSS IBIAS IBIAS OUT VSS sky130_fd_pr__nfet_g5v0d10v5_N5GNFR
Xsky130_fd_pr__nfet_g5v0d10v5_X6KG9Z_0 m1_2160_1440# m1_2740_n3440# VP VP m1_2160_1440#
+ VP VP m1_2160_1440# VSS m1_2740_n3440# sky130_fd_pr__nfet_g5v0d10v5_X6KG9Z
Xsky130_fd_pr__cap_mim_m3_1_R7S84X_0 m1_n1120_1120# m1_n2200_3200# VSS sky130_fd_pr__cap_mim_m3_1_R7S84X
Xsky130_fd_pr__nfet_g5v0d10v5_N5GNFR_0 IBIAS IBIAS VSS OUT OUT VSS IBIAS IBIAS OUT
+ VSS sky130_fd_pr__nfet_g5v0d10v5_N5GNFR
Xsky130_fd_pr__nfet_g5v0d10v5_PBQQNH_0 m1_n1120_1120# m1_2740_n3440# VN VN m1_n1120_1120#
+ VN VN m1_n1120_1120# VSS m1_2740_n3440# sky130_fd_pr__nfet_g5v0d10v5_PBQQNH
Xsky130_fd_pr__pfet_g5v0d10v5_V6JW4R_0 OUT VSS OUT m1_n2200_3200# VDD VSS VSS sky130_fd_pr__pfet_g5v0d10v5_V6JW4R
C0 m1_n1120_1120# OUT 2.31052f
C1 VDD m1_2160_1440# 9.96962f
C2 OUT IBIAS 1.15932f
C3 OUT VP 0.09958f
C4 m1_n1120_1120# VDD 19.54036f
C5 VN m1_2740_n3440# 0.66005f
C6 VN VSS 1.58934f
C7 VDD VP 0.01582f
C8 VN m1_2160_1440# 1.16845f
C9 m1_n1120_1120# VN 2.95636f
C10 m1_2740_n3440# VSS 1.40409f
C11 m1_n2200_3200# VSS 2.97735f
C12 VN IBIAS 0.47606f
C13 VDD OUT 6.46108f
C14 VN VP 0.3521f
C15 m1_2160_1440# m1_2740_n3440# 4.90242f
C16 m1_2160_1440# VSS 2.31782f
C17 m1_n1120_1120# m1_2740_n3440# 3.65355f
C18 m1_n1120_1120# m1_n2200_3200# 1.4767f
C19 m1_n1120_1120# VSS 1.06936f
C20 IBIAS m1_2740_n3440# 2.03627f
C21 IBIAS m1_n2200_3200# 0.19595f
C22 VN OUT 0.08699f
C23 IBIAS VSS 12.9339f
C24 VP m1_2740_n3440# 0.80903f
C25 VP VSS 1.56228f
C26 m1_n1120_1120# m1_2160_1440# 14.16827f
C27 VDD VN 0.01778f
C28 m1_2160_1440# IBIAS 0.58216f
C29 m1_2160_1440# VP 1.2916f
C30 m1_n1120_1120# IBIAS 0.58047f
C31 OUT m1_n2200_3200# 6.50839f
C32 OUT VSS 4.857f
C33 m1_n1120_1120# VP 3.39887f
C34 IBIAS VP 0.44611f
C35 VDD m1_2740_n3440# 0.14829f
C36 VDD m1_n2200_3200# 1.86773f
C37 VDD VSS 1.58824f
C38 OUT m1_2160_1440# 0.3293f
C39 m1_n2200_3200# 0 31.55975f
C40 m1_n1120_1120# 0 0.11133p
C41 VN 0 4.40862f
C42 VSS 0 22.34968f
C43 OUT 0 23.03029f
C44 m1_2160_1440# 0 11.22809f
C45 m1_2740_n3440# 0 3.88057f
C46 IBIAS 0 14.08802f
C47 VP 0 3.26044f
C48 VDD 0 0.10583p
.ends

