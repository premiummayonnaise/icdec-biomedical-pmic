magic
tech sky130A
magscale 1 2
timestamp 1768990256
<< mvnmos >>
rect -467 -440 -367 502
rect -189 -440 -89 502
rect 89 -440 189 502
rect 367 -440 467 502
<< mvndiff >>
rect -525 490 -467 502
rect -525 -428 -513 490
rect -479 -428 -467 490
rect -525 -440 -467 -428
rect -367 490 -309 502
rect -367 -428 -355 490
rect -321 -428 -309 490
rect -367 -440 -309 -428
rect -247 490 -189 502
rect -247 -428 -235 490
rect -201 -428 -189 490
rect -247 -440 -189 -428
rect -89 490 -31 502
rect -89 -428 -77 490
rect -43 -428 -31 490
rect -89 -440 -31 -428
rect 31 490 89 502
rect 31 -428 43 490
rect 77 -428 89 490
rect 31 -440 89 -428
rect 189 490 247 502
rect 189 -428 201 490
rect 235 -428 247 490
rect 189 -440 247 -428
rect 309 490 367 502
rect 309 -428 321 490
rect 355 -428 367 490
rect 309 -440 367 -428
rect 467 490 525 502
rect 467 -428 479 490
rect 513 -428 525 490
rect 467 -440 525 -428
<< mvndiffc >>
rect -513 -428 -479 490
rect -355 -428 -321 490
rect -235 -428 -201 490
rect -77 -428 -43 490
rect 43 -428 77 490
rect 201 -428 235 490
rect 321 -428 355 490
rect 479 -428 513 490
<< poly >>
rect -467 502 -367 528
rect -189 502 -89 528
rect 89 502 189 528
rect 367 502 467 528
rect -467 -478 -367 -440
rect -467 -512 -451 -478
rect -383 -512 -367 -478
rect -467 -528 -367 -512
rect -189 -478 -89 -440
rect -189 -512 -173 -478
rect -105 -512 -89 -478
rect -189 -528 -89 -512
rect 89 -478 189 -440
rect 89 -512 105 -478
rect 173 -512 189 -478
rect 89 -528 189 -512
rect 367 -478 467 -440
rect 367 -512 383 -478
rect 451 -512 467 -478
rect 367 -528 467 -512
<< polycont >>
rect -451 -512 -383 -478
rect -173 -512 -105 -478
rect 105 -512 173 -478
rect 383 -512 451 -478
<< locali >>
rect -513 490 -479 506
rect -513 -444 -479 -428
rect -355 490 -321 506
rect -355 -444 -321 -428
rect -235 490 -201 506
rect -235 -444 -201 -428
rect -77 490 -43 506
rect -77 -444 -43 -428
rect 43 490 77 506
rect 43 -444 77 -428
rect 201 490 235 506
rect 201 -444 235 -428
rect 321 490 355 506
rect 321 -444 355 -428
rect 479 490 513 506
rect 479 -444 513 -428
rect -467 -512 -451 -478
rect -383 -512 -367 -478
rect -189 -512 -173 -478
rect -105 -512 -89 -478
rect 89 -512 105 -478
rect 173 -512 189 -478
rect 367 -512 383 -478
rect 451 -512 467 -478
<< viali >>
rect -513 -428 -479 490
rect -355 -428 -321 490
rect -235 -428 -201 490
rect -77 -428 -43 490
rect 43 -428 77 490
rect 201 -428 235 490
rect 321 -428 355 490
rect 479 -428 513 490
rect -451 -512 -383 -478
rect -173 -512 -105 -478
rect 105 -512 173 -478
rect 383 -512 451 -478
<< metal1 >>
rect -519 490 -473 502
rect -519 -428 -513 490
rect -479 -428 -473 490
rect -519 -440 -473 -428
rect -361 490 -315 502
rect -361 -428 -355 490
rect -321 -428 -315 490
rect -361 -440 -315 -428
rect -241 490 -195 502
rect -241 -428 -235 490
rect -201 -428 -195 490
rect -241 -440 -195 -428
rect -83 490 -37 502
rect -83 -428 -77 490
rect -43 -428 -37 490
rect -83 -440 -37 -428
rect 37 490 83 502
rect 37 -428 43 490
rect 77 -428 83 490
rect 37 -440 83 -428
rect 195 490 241 502
rect 195 -428 201 490
rect 235 -428 241 490
rect 195 -440 241 -428
rect 315 490 361 502
rect 315 -428 321 490
rect 355 -428 361 490
rect 315 -440 361 -428
rect 473 490 519 502
rect 473 -428 479 490
rect 513 -428 519 490
rect 473 -440 519 -428
rect -463 -478 -371 -472
rect -463 -512 -451 -478
rect -383 -512 -371 -478
rect -463 -518 -371 -512
rect -185 -478 -93 -472
rect -185 -512 -173 -478
rect -105 -512 -93 -478
rect -185 -518 -93 -512
rect 93 -478 185 -472
rect 93 -512 105 -478
rect 173 -512 185 -478
rect 93 -518 185 -512
rect 371 -478 463 -472
rect 371 -512 383 -478
rect 451 -512 463 -478
rect 371 -518 463 -512
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.7125 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
