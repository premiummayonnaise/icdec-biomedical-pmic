magic
tech sky130A
magscale 1 2
timestamp 1769135993
<< pwell >>
rect -791 -315 791 315
<< nmos >>
rect -595 -105 -445 105
rect -387 -105 -237 105
rect -179 -105 -29 105
rect 29 -105 179 105
rect 237 -105 387 105
rect 445 -105 595 105
<< ndiff >>
rect -653 93 -595 105
rect -653 -93 -641 93
rect -607 -93 -595 93
rect -653 -105 -595 -93
rect -445 93 -387 105
rect -445 -93 -433 93
rect -399 -93 -387 93
rect -445 -105 -387 -93
rect -237 93 -179 105
rect -237 -93 -225 93
rect -191 -93 -179 93
rect -237 -105 -179 -93
rect -29 93 29 105
rect -29 -93 -17 93
rect 17 -93 29 93
rect -29 -105 29 -93
rect 179 93 237 105
rect 179 -93 191 93
rect 225 -93 237 93
rect 179 -105 237 -93
rect 387 93 445 105
rect 387 -93 399 93
rect 433 -93 445 93
rect 387 -105 445 -93
rect 595 93 653 105
rect 595 -93 607 93
rect 641 -93 653 93
rect 595 -105 653 -93
<< ndiffc >>
rect -641 -93 -607 93
rect -433 -93 -399 93
rect -225 -93 -191 93
rect -17 -93 17 93
rect 191 -93 225 93
rect 399 -93 433 93
rect 607 -93 641 93
<< psubdiff >>
rect -755 245 -659 279
rect 659 245 755 279
rect -755 183 -721 245
rect 721 183 755 245
rect -755 -245 -721 -183
rect 721 -245 755 -183
rect -755 -279 -659 -245
rect 659 -279 755 -245
<< psubdiffcont >>
rect -659 245 659 279
rect -755 -183 -721 183
rect 721 -183 755 183
rect -659 -279 659 -245
<< poly >>
rect -595 177 -445 193
rect -595 143 -579 177
rect -461 143 -445 177
rect -595 105 -445 143
rect -387 177 -237 193
rect -387 143 -371 177
rect -253 143 -237 177
rect -387 105 -237 143
rect -179 177 -29 193
rect -179 143 -163 177
rect -45 143 -29 177
rect -179 105 -29 143
rect 29 177 179 193
rect 29 143 45 177
rect 163 143 179 177
rect 29 105 179 143
rect 237 177 387 193
rect 237 143 253 177
rect 371 143 387 177
rect 237 105 387 143
rect 445 177 595 193
rect 445 143 461 177
rect 579 143 595 177
rect 445 105 595 143
rect -595 -143 -445 -105
rect -595 -177 -579 -143
rect -461 -177 -445 -143
rect -595 -193 -445 -177
rect -387 -143 -237 -105
rect -387 -177 -371 -143
rect -253 -177 -237 -143
rect -387 -193 -237 -177
rect -179 -143 -29 -105
rect -179 -177 -163 -143
rect -45 -177 -29 -143
rect -179 -193 -29 -177
rect 29 -143 179 -105
rect 29 -177 45 -143
rect 163 -177 179 -143
rect 29 -193 179 -177
rect 237 -143 387 -105
rect 237 -177 253 -143
rect 371 -177 387 -143
rect 237 -193 387 -177
rect 445 -143 595 -105
rect 445 -177 461 -143
rect 579 -177 595 -143
rect 445 -193 595 -177
<< polycont >>
rect -579 143 -461 177
rect -371 143 -253 177
rect -163 143 -45 177
rect 45 143 163 177
rect 253 143 371 177
rect 461 143 579 177
rect -579 -177 -461 -143
rect -371 -177 -253 -143
rect -163 -177 -45 -143
rect 45 -177 163 -143
rect 253 -177 371 -143
rect 461 -177 579 -143
<< locali >>
rect -755 245 -659 279
rect 659 245 755 279
rect -755 183 -721 245
rect 721 183 755 245
rect -595 143 -579 177
rect -461 143 -445 177
rect -387 143 -371 177
rect -253 143 -237 177
rect -179 143 -163 177
rect -45 143 -29 177
rect 29 143 45 177
rect 163 143 179 177
rect 237 143 253 177
rect 371 143 387 177
rect 445 143 461 177
rect 579 143 595 177
rect -641 93 -607 109
rect -641 -109 -607 -93
rect -433 93 -399 109
rect -433 -109 -399 -93
rect -225 93 -191 109
rect -225 -109 -191 -93
rect -17 93 17 109
rect -17 -109 17 -93
rect 191 93 225 109
rect 191 -109 225 -93
rect 399 93 433 109
rect 399 -109 433 -93
rect 607 93 641 109
rect 607 -109 641 -93
rect -595 -177 -579 -143
rect -461 -177 -445 -143
rect -387 -177 -371 -143
rect -253 -177 -237 -143
rect -179 -177 -163 -143
rect -45 -177 -29 -143
rect 29 -177 45 -143
rect 163 -177 179 -143
rect 237 -177 253 -143
rect 371 -177 387 -143
rect 445 -177 461 -143
rect 579 -177 595 -143
rect -755 -245 -721 -183
rect 721 -245 755 -183
rect -755 -279 -659 -245
rect 659 -279 755 -245
<< viali >>
rect -579 143 -461 177
rect -371 143 -253 177
rect -163 143 -45 177
rect 45 143 163 177
rect 253 143 371 177
rect 461 143 579 177
rect -641 -93 -607 93
rect -433 -93 -399 93
rect -225 -93 -191 93
rect -17 -93 17 93
rect 191 -93 225 93
rect 399 -93 433 93
rect 607 -93 641 93
rect -579 -177 -461 -143
rect -371 -177 -253 -143
rect -163 -177 -45 -143
rect 45 -177 163 -143
rect 253 -177 371 -143
rect 461 -177 579 -143
<< metal1 >>
rect -591 177 -449 183
rect -591 143 -579 177
rect -461 143 -449 177
rect -591 137 -449 143
rect -383 177 -241 183
rect -383 143 -371 177
rect -253 143 -241 177
rect -383 137 -241 143
rect -175 177 -33 183
rect -175 143 -163 177
rect -45 143 -33 177
rect -175 137 -33 143
rect 33 177 175 183
rect 33 143 45 177
rect 163 143 175 177
rect 33 137 175 143
rect 241 177 383 183
rect 241 143 253 177
rect 371 143 383 177
rect 241 137 383 143
rect 449 177 591 183
rect 449 143 461 177
rect 579 143 591 177
rect 449 137 591 143
rect -647 93 -601 105
rect -647 -93 -641 93
rect -607 -93 -601 93
rect -647 -105 -601 -93
rect -439 93 -393 105
rect -439 -93 -433 93
rect -399 -93 -393 93
rect -439 -105 -393 -93
rect -231 93 -185 105
rect -231 -93 -225 93
rect -191 -93 -185 93
rect -231 -105 -185 -93
rect -23 93 23 105
rect -23 -93 -17 93
rect 17 -93 23 93
rect -23 -105 23 -93
rect 185 93 231 105
rect 185 -93 191 93
rect 225 -93 231 93
rect 185 -105 231 -93
rect 393 93 439 105
rect 393 -93 399 93
rect 433 -93 439 93
rect 393 -105 439 -93
rect 601 93 647 105
rect 601 -93 607 93
rect 641 -93 647 93
rect 601 -105 647 -93
rect -591 -143 -449 -137
rect -591 -177 -579 -143
rect -461 -177 -449 -143
rect -591 -183 -449 -177
rect -383 -143 -241 -137
rect -383 -177 -371 -143
rect -253 -177 -241 -143
rect -383 -183 -241 -177
rect -175 -143 -33 -137
rect -175 -177 -163 -143
rect -45 -177 -33 -143
rect -175 -183 -33 -177
rect 33 -143 175 -137
rect 33 -177 45 -143
rect 163 -177 175 -143
rect 33 -183 175 -177
rect 241 -143 383 -137
rect 241 -177 253 -143
rect 371 -177 383 -143
rect 241 -183 383 -177
rect 449 -143 591 -137
rect 449 -177 461 -143
rect 579 -177 591 -143
rect 449 -183 591 -177
<< properties >>
string FIXED_BBOX -738 -262 738 262
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.05 l 0.75 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
