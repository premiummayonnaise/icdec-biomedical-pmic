magic
tech sky130A
magscale 1 2
timestamp 1768990256
<< mvnmos >>
rect -467 -502 -367 440
rect -189 -502 -89 440
rect 89 -502 189 440
rect 367 -502 467 440
<< mvndiff >>
rect -525 428 -467 440
rect -525 -490 -513 428
rect -479 -490 -467 428
rect -525 -502 -467 -490
rect -367 428 -309 440
rect -367 -490 -355 428
rect -321 -490 -309 428
rect -367 -502 -309 -490
rect -247 428 -189 440
rect -247 -490 -235 428
rect -201 -490 -189 428
rect -247 -502 -189 -490
rect -89 428 -31 440
rect -89 -490 -77 428
rect -43 -490 -31 428
rect -89 -502 -31 -490
rect 31 428 89 440
rect 31 -490 43 428
rect 77 -490 89 428
rect 31 -502 89 -490
rect 189 428 247 440
rect 189 -490 201 428
rect 235 -490 247 428
rect 189 -502 247 -490
rect 309 428 367 440
rect 309 -490 321 428
rect 355 -490 367 428
rect 309 -502 367 -490
rect 467 428 525 440
rect 467 -490 479 428
rect 513 -490 525 428
rect 467 -502 525 -490
<< mvndiffc >>
rect -513 -490 -479 428
rect -355 -490 -321 428
rect -235 -490 -201 428
rect -77 -490 -43 428
rect 43 -490 77 428
rect 201 -490 235 428
rect 321 -490 355 428
rect 479 -490 513 428
<< poly >>
rect -467 512 -367 528
rect -467 478 -451 512
rect -383 478 -367 512
rect -467 440 -367 478
rect -189 512 -89 528
rect -189 478 -173 512
rect -105 478 -89 512
rect -189 440 -89 478
rect 89 512 189 528
rect 89 478 105 512
rect 173 478 189 512
rect 89 440 189 478
rect 367 512 467 528
rect 367 478 383 512
rect 451 478 467 512
rect 367 440 467 478
rect -467 -528 -367 -502
rect -189 -528 -89 -502
rect 89 -528 189 -502
rect 367 -528 467 -502
<< polycont >>
rect -451 478 -383 512
rect -173 478 -105 512
rect 105 478 173 512
rect 383 478 451 512
<< locali >>
rect -467 478 -451 512
rect -383 478 -367 512
rect -189 478 -173 512
rect -105 478 -89 512
rect 89 478 105 512
rect 173 478 189 512
rect 367 478 383 512
rect 451 478 467 512
rect -513 428 -479 444
rect -513 -506 -479 -490
rect -355 428 -321 444
rect -355 -506 -321 -490
rect -235 428 -201 444
rect -235 -506 -201 -490
rect -77 428 -43 444
rect -77 -506 -43 -490
rect 43 428 77 444
rect 43 -506 77 -490
rect 201 428 235 444
rect 201 -506 235 -490
rect 321 428 355 444
rect 321 -506 355 -490
rect 479 428 513 444
rect 479 -506 513 -490
<< viali >>
rect -451 478 -383 512
rect -173 478 -105 512
rect 105 478 173 512
rect 383 478 451 512
rect -513 -490 -479 428
rect -355 -490 -321 428
rect -235 -490 -201 428
rect -77 -490 -43 428
rect 43 -490 77 428
rect 201 -490 235 428
rect 321 -490 355 428
rect 479 -490 513 428
<< metal1 >>
rect -463 512 -371 518
rect -463 478 -451 512
rect -383 478 -371 512
rect -463 472 -371 478
rect -185 512 -93 518
rect -185 478 -173 512
rect -105 478 -93 512
rect -185 472 -93 478
rect 93 512 185 518
rect 93 478 105 512
rect 173 478 185 512
rect 93 472 185 478
rect 371 512 463 518
rect 371 478 383 512
rect 451 478 463 512
rect 371 472 463 478
rect -519 428 -473 440
rect -519 -490 -513 428
rect -479 -490 -473 428
rect -519 -502 -473 -490
rect -361 428 -315 440
rect -361 -490 -355 428
rect -321 -490 -315 428
rect -361 -502 -315 -490
rect -241 428 -195 440
rect -241 -490 -235 428
rect -201 -490 -195 428
rect -241 -502 -195 -490
rect -83 428 -37 440
rect -83 -490 -77 428
rect -43 -490 -37 428
rect -83 -502 -37 -490
rect 37 428 83 440
rect 37 -490 43 428
rect 77 -490 83 428
rect 37 -502 83 -490
rect 195 428 241 440
rect 195 -490 201 428
rect 235 -490 241 428
rect 195 -502 241 -490
rect 315 428 361 440
rect 315 -490 321 428
rect 355 -490 361 428
rect 315 -502 361 -490
rect 473 428 519 440
rect 473 -490 479 428
rect 513 -490 519 428
rect 473 -502 519 -490
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.7125 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
