magic
tech sky130A
magscale 1 2
timestamp 1770083657
<< pwell >>
rect -371 -532 371 470
<< mvnmos >>
rect -287 -506 -187 444
rect -129 -506 -29 444
rect 29 -506 129 444
rect 187 -506 287 444
<< mvndiff >>
rect -345 326 -287 444
rect -345 292 -333 326
rect -299 292 -287 326
rect -345 258 -287 292
rect -345 224 -333 258
rect -299 224 -287 258
rect -345 190 -287 224
rect -345 156 -333 190
rect -299 156 -287 190
rect -345 122 -287 156
rect -345 88 -333 122
rect -299 88 -287 122
rect -345 54 -287 88
rect -345 20 -333 54
rect -299 20 -287 54
rect -345 -14 -287 20
rect -345 -48 -333 -14
rect -299 -48 -287 -14
rect -345 -82 -287 -48
rect -345 -116 -333 -82
rect -299 -116 -287 -82
rect -345 -150 -287 -116
rect -345 -184 -333 -150
rect -299 -184 -287 -150
rect -345 -218 -287 -184
rect -345 -252 -333 -218
rect -299 -252 -287 -218
rect -345 -286 -287 -252
rect -345 -320 -333 -286
rect -299 -320 -287 -286
rect -345 -354 -287 -320
rect -345 -388 -333 -354
rect -299 -388 -287 -354
rect -345 -506 -287 -388
rect -187 326 -129 444
rect -187 292 -175 326
rect -141 292 -129 326
rect -187 258 -129 292
rect -187 224 -175 258
rect -141 224 -129 258
rect -187 190 -129 224
rect -187 156 -175 190
rect -141 156 -129 190
rect -187 122 -129 156
rect -187 88 -175 122
rect -141 88 -129 122
rect -187 54 -129 88
rect -187 20 -175 54
rect -141 20 -129 54
rect -187 -14 -129 20
rect -187 -48 -175 -14
rect -141 -48 -129 -14
rect -187 -82 -129 -48
rect -187 -116 -175 -82
rect -141 -116 -129 -82
rect -187 -150 -129 -116
rect -187 -184 -175 -150
rect -141 -184 -129 -150
rect -187 -218 -129 -184
rect -187 -252 -175 -218
rect -141 -252 -129 -218
rect -187 -286 -129 -252
rect -187 -320 -175 -286
rect -141 -320 -129 -286
rect -187 -354 -129 -320
rect -187 -388 -175 -354
rect -141 -388 -129 -354
rect -187 -506 -129 -388
rect -29 326 29 444
rect -29 292 -17 326
rect 17 292 29 326
rect -29 258 29 292
rect -29 224 -17 258
rect 17 224 29 258
rect -29 190 29 224
rect -29 156 -17 190
rect 17 156 29 190
rect -29 122 29 156
rect -29 88 -17 122
rect 17 88 29 122
rect -29 54 29 88
rect -29 20 -17 54
rect 17 20 29 54
rect -29 -14 29 20
rect -29 -48 -17 -14
rect 17 -48 29 -14
rect -29 -82 29 -48
rect -29 -116 -17 -82
rect 17 -116 29 -82
rect -29 -150 29 -116
rect -29 -184 -17 -150
rect 17 -184 29 -150
rect -29 -218 29 -184
rect -29 -252 -17 -218
rect 17 -252 29 -218
rect -29 -286 29 -252
rect -29 -320 -17 -286
rect 17 -320 29 -286
rect -29 -354 29 -320
rect -29 -388 -17 -354
rect 17 -388 29 -354
rect -29 -506 29 -388
rect 129 326 187 444
rect 129 292 141 326
rect 175 292 187 326
rect 129 258 187 292
rect 129 224 141 258
rect 175 224 187 258
rect 129 190 187 224
rect 129 156 141 190
rect 175 156 187 190
rect 129 122 187 156
rect 129 88 141 122
rect 175 88 187 122
rect 129 54 187 88
rect 129 20 141 54
rect 175 20 187 54
rect 129 -14 187 20
rect 129 -48 141 -14
rect 175 -48 187 -14
rect 129 -82 187 -48
rect 129 -116 141 -82
rect 175 -116 187 -82
rect 129 -150 187 -116
rect 129 -184 141 -150
rect 175 -184 187 -150
rect 129 -218 187 -184
rect 129 -252 141 -218
rect 175 -252 187 -218
rect 129 -286 187 -252
rect 129 -320 141 -286
rect 175 -320 187 -286
rect 129 -354 187 -320
rect 129 -388 141 -354
rect 175 -388 187 -354
rect 129 -506 187 -388
rect 287 326 345 444
rect 287 292 299 326
rect 333 292 345 326
rect 287 258 345 292
rect 287 224 299 258
rect 333 224 345 258
rect 287 190 345 224
rect 287 156 299 190
rect 333 156 345 190
rect 287 122 345 156
rect 287 88 299 122
rect 333 88 345 122
rect 287 54 345 88
rect 287 20 299 54
rect 333 20 345 54
rect 287 -14 345 20
rect 287 -48 299 -14
rect 333 -48 345 -14
rect 287 -82 345 -48
rect 287 -116 299 -82
rect 333 -116 345 -82
rect 287 -150 345 -116
rect 287 -184 299 -150
rect 333 -184 345 -150
rect 287 -218 345 -184
rect 287 -252 299 -218
rect 333 -252 345 -218
rect 287 -286 345 -252
rect 287 -320 299 -286
rect 333 -320 345 -286
rect 287 -354 345 -320
rect 287 -388 299 -354
rect 333 -388 345 -354
rect 287 -506 345 -388
<< mvndiffc >>
rect -333 292 -299 326
rect -333 224 -299 258
rect -333 156 -299 190
rect -333 88 -299 122
rect -333 20 -299 54
rect -333 -48 -299 -14
rect -333 -116 -299 -82
rect -333 -184 -299 -150
rect -333 -252 -299 -218
rect -333 -320 -299 -286
rect -333 -388 -299 -354
rect -175 292 -141 326
rect -175 224 -141 258
rect -175 156 -141 190
rect -175 88 -141 122
rect -175 20 -141 54
rect -175 -48 -141 -14
rect -175 -116 -141 -82
rect -175 -184 -141 -150
rect -175 -252 -141 -218
rect -175 -320 -141 -286
rect -175 -388 -141 -354
rect -17 292 17 326
rect -17 224 17 258
rect -17 156 17 190
rect -17 88 17 122
rect -17 20 17 54
rect -17 -48 17 -14
rect -17 -116 17 -82
rect -17 -184 17 -150
rect -17 -252 17 -218
rect -17 -320 17 -286
rect -17 -388 17 -354
rect 141 292 175 326
rect 141 224 175 258
rect 141 156 175 190
rect 141 88 175 122
rect 141 20 175 54
rect 141 -48 175 -14
rect 141 -116 175 -82
rect 141 -184 175 -150
rect 141 -252 175 -218
rect 141 -320 175 -286
rect 141 -388 175 -354
rect 299 292 333 326
rect 299 224 333 258
rect 299 156 333 190
rect 299 88 333 122
rect 299 20 333 54
rect 299 -48 333 -14
rect 299 -116 333 -82
rect 299 -184 333 -150
rect 299 -252 333 -218
rect 299 -320 333 -286
rect 299 -388 333 -354
<< poly >>
rect -287 516 -187 532
rect -287 482 -254 516
rect -220 482 -187 516
rect -287 444 -187 482
rect -129 516 -29 532
rect -129 482 -96 516
rect -62 482 -29 516
rect -129 444 -29 482
rect 29 516 129 532
rect 29 482 62 516
rect 96 482 129 516
rect 29 444 129 482
rect 187 516 287 532
rect 187 482 220 516
rect 254 482 287 516
rect 187 444 287 482
rect -287 -532 -187 -506
rect -129 -532 -29 -506
rect 29 -532 129 -506
rect 187 -532 287 -506
<< polycont >>
rect -254 482 -220 516
rect -96 482 -62 516
rect 62 482 96 516
rect 220 482 254 516
<< locali >>
rect -287 482 -254 516
rect -220 482 -187 516
rect -129 482 -96 516
rect -62 482 -29 516
rect 29 482 62 516
rect 96 482 129 516
rect 187 482 220 516
rect 254 482 287 516
rect -333 326 -299 355
rect -333 258 -299 276
rect -333 190 -299 204
rect -333 122 -299 132
rect -333 54 -299 60
rect -333 -14 -299 -12
rect -333 -50 -299 -48
rect -333 -122 -299 -116
rect -333 -194 -299 -184
rect -333 -266 -299 -252
rect -333 -338 -299 -320
rect -333 -417 -299 -388
rect -175 326 -141 355
rect -175 258 -141 276
rect -175 190 -141 204
rect -175 122 -141 132
rect -175 54 -141 60
rect -175 -14 -141 -12
rect -175 -50 -141 -48
rect -175 -122 -141 -116
rect -175 -194 -141 -184
rect -175 -266 -141 -252
rect -175 -338 -141 -320
rect -175 -417 -141 -388
rect -17 326 17 355
rect -17 258 17 276
rect -17 190 17 204
rect -17 122 17 132
rect -17 54 17 60
rect -17 -14 17 -12
rect -17 -50 17 -48
rect -17 -122 17 -116
rect -17 -194 17 -184
rect -17 -266 17 -252
rect -17 -338 17 -320
rect -17 -417 17 -388
rect 141 326 175 355
rect 141 258 175 276
rect 141 190 175 204
rect 141 122 175 132
rect 141 54 175 60
rect 141 -14 175 -12
rect 141 -50 175 -48
rect 141 -122 175 -116
rect 141 -194 175 -184
rect 141 -266 175 -252
rect 141 -338 175 -320
rect 141 -417 175 -388
rect 299 326 333 355
rect 299 258 333 276
rect 299 190 333 204
rect 299 122 333 132
rect 299 54 333 60
rect 299 -14 333 -12
rect 299 -50 333 -48
rect 299 -122 333 -116
rect 299 -194 333 -184
rect 299 -266 333 -252
rect 299 -338 333 -320
rect 299 -417 333 -388
<< viali >>
rect -254 482 -220 516
rect -96 482 -62 516
rect 62 482 96 516
rect 220 482 254 516
rect -333 292 -299 310
rect -333 276 -299 292
rect -333 224 -299 238
rect -333 204 -299 224
rect -333 156 -299 166
rect -333 132 -299 156
rect -333 88 -299 94
rect -333 60 -299 88
rect -333 20 -299 22
rect -333 -12 -299 20
rect -333 -82 -299 -50
rect -333 -84 -299 -82
rect -333 -150 -299 -122
rect -333 -156 -299 -150
rect -333 -218 -299 -194
rect -333 -228 -299 -218
rect -333 -286 -299 -266
rect -333 -300 -299 -286
rect -333 -354 -299 -338
rect -333 -372 -299 -354
rect -175 292 -141 310
rect -175 276 -141 292
rect -175 224 -141 238
rect -175 204 -141 224
rect -175 156 -141 166
rect -175 132 -141 156
rect -175 88 -141 94
rect -175 60 -141 88
rect -175 20 -141 22
rect -175 -12 -141 20
rect -175 -82 -141 -50
rect -175 -84 -141 -82
rect -175 -150 -141 -122
rect -175 -156 -141 -150
rect -175 -218 -141 -194
rect -175 -228 -141 -218
rect -175 -286 -141 -266
rect -175 -300 -141 -286
rect -175 -354 -141 -338
rect -175 -372 -141 -354
rect -17 292 17 310
rect -17 276 17 292
rect -17 224 17 238
rect -17 204 17 224
rect -17 156 17 166
rect -17 132 17 156
rect -17 88 17 94
rect -17 60 17 88
rect -17 20 17 22
rect -17 -12 17 20
rect -17 -82 17 -50
rect -17 -84 17 -82
rect -17 -150 17 -122
rect -17 -156 17 -150
rect -17 -218 17 -194
rect -17 -228 17 -218
rect -17 -286 17 -266
rect -17 -300 17 -286
rect -17 -354 17 -338
rect -17 -372 17 -354
rect 141 292 175 310
rect 141 276 175 292
rect 141 224 175 238
rect 141 204 175 224
rect 141 156 175 166
rect 141 132 175 156
rect 141 88 175 94
rect 141 60 175 88
rect 141 20 175 22
rect 141 -12 175 20
rect 141 -82 175 -50
rect 141 -84 175 -82
rect 141 -150 175 -122
rect 141 -156 175 -150
rect 141 -218 175 -194
rect 141 -228 175 -218
rect 141 -286 175 -266
rect 141 -300 175 -286
rect 141 -354 175 -338
rect 141 -372 175 -354
rect 299 292 333 310
rect 299 276 333 292
rect 299 224 333 238
rect 299 204 333 224
rect 299 156 333 166
rect 299 132 333 156
rect 299 88 333 94
rect 299 60 333 88
rect 299 20 333 22
rect 299 -12 333 20
rect 299 -82 333 -50
rect 299 -84 333 -82
rect 299 -150 333 -122
rect 299 -156 333 -150
rect 299 -218 333 -194
rect 299 -228 333 -218
rect 299 -286 333 -266
rect 299 -300 333 -286
rect 299 -354 333 -338
rect 299 -372 333 -354
<< metal1 >>
rect -283 516 -191 522
rect -283 482 -254 516
rect -220 482 -191 516
rect -283 476 -191 482
rect -125 516 -33 522
rect -125 482 -96 516
rect -62 482 -33 516
rect -125 476 -33 482
rect 33 516 125 522
rect 33 482 62 516
rect 96 482 125 516
rect 33 476 125 482
rect 191 516 283 522
rect 191 482 220 516
rect 254 482 283 516
rect 191 476 283 482
rect -339 310 -293 351
rect -339 276 -333 310
rect -299 276 -293 310
rect -339 238 -293 276
rect -339 204 -333 238
rect -299 204 -293 238
rect -339 166 -293 204
rect -339 132 -333 166
rect -299 132 -293 166
rect -339 94 -293 132
rect -339 60 -333 94
rect -299 60 -293 94
rect -339 22 -293 60
rect -339 -12 -333 22
rect -299 -12 -293 22
rect -339 -50 -293 -12
rect -339 -84 -333 -50
rect -299 -84 -293 -50
rect -339 -122 -293 -84
rect -339 -156 -333 -122
rect -299 -156 -293 -122
rect -339 -194 -293 -156
rect -339 -228 -333 -194
rect -299 -228 -293 -194
rect -339 -266 -293 -228
rect -339 -300 -333 -266
rect -299 -300 -293 -266
rect -339 -338 -293 -300
rect -339 -372 -333 -338
rect -299 -372 -293 -338
rect -339 -413 -293 -372
rect -181 310 -135 351
rect -181 276 -175 310
rect -141 276 -135 310
rect -181 238 -135 276
rect -181 204 -175 238
rect -141 204 -135 238
rect -181 166 -135 204
rect -181 132 -175 166
rect -141 132 -135 166
rect -181 94 -135 132
rect -181 60 -175 94
rect -141 60 -135 94
rect -181 22 -135 60
rect -181 -12 -175 22
rect -141 -12 -135 22
rect -181 -50 -135 -12
rect -181 -84 -175 -50
rect -141 -84 -135 -50
rect -181 -122 -135 -84
rect -181 -156 -175 -122
rect -141 -156 -135 -122
rect -181 -194 -135 -156
rect -181 -228 -175 -194
rect -141 -228 -135 -194
rect -181 -266 -135 -228
rect -181 -300 -175 -266
rect -141 -300 -135 -266
rect -181 -338 -135 -300
rect -181 -372 -175 -338
rect -141 -372 -135 -338
rect -181 -413 -135 -372
rect -23 310 23 351
rect -23 276 -17 310
rect 17 276 23 310
rect -23 238 23 276
rect -23 204 -17 238
rect 17 204 23 238
rect -23 166 23 204
rect -23 132 -17 166
rect 17 132 23 166
rect -23 94 23 132
rect -23 60 -17 94
rect 17 60 23 94
rect -23 22 23 60
rect -23 -12 -17 22
rect 17 -12 23 22
rect -23 -50 23 -12
rect -23 -84 -17 -50
rect 17 -84 23 -50
rect -23 -122 23 -84
rect -23 -156 -17 -122
rect 17 -156 23 -122
rect -23 -194 23 -156
rect -23 -228 -17 -194
rect 17 -228 23 -194
rect -23 -266 23 -228
rect -23 -300 -17 -266
rect 17 -300 23 -266
rect -23 -338 23 -300
rect -23 -372 -17 -338
rect 17 -372 23 -338
rect -23 -413 23 -372
rect 135 310 181 351
rect 135 276 141 310
rect 175 276 181 310
rect 135 238 181 276
rect 135 204 141 238
rect 175 204 181 238
rect 135 166 181 204
rect 135 132 141 166
rect 175 132 181 166
rect 135 94 181 132
rect 135 60 141 94
rect 175 60 181 94
rect 135 22 181 60
rect 135 -12 141 22
rect 175 -12 181 22
rect 135 -50 181 -12
rect 135 -84 141 -50
rect 175 -84 181 -50
rect 135 -122 181 -84
rect 135 -156 141 -122
rect 175 -156 181 -122
rect 135 -194 181 -156
rect 135 -228 141 -194
rect 175 -228 181 -194
rect 135 -266 181 -228
rect 135 -300 141 -266
rect 175 -300 181 -266
rect 135 -338 181 -300
rect 135 -372 141 -338
rect 175 -372 181 -338
rect 135 -413 181 -372
rect 293 310 339 351
rect 293 276 299 310
rect 333 276 339 310
rect 293 238 339 276
rect 293 204 299 238
rect 333 204 339 238
rect 293 166 339 204
rect 293 132 299 166
rect 333 132 339 166
rect 293 94 339 132
rect 293 60 299 94
rect 333 60 339 94
rect 293 22 339 60
rect 293 -12 299 22
rect 333 -12 339 22
rect 293 -50 339 -12
rect 293 -84 299 -50
rect 333 -84 339 -50
rect 293 -122 339 -84
rect 293 -156 299 -122
rect 333 -156 339 -122
rect 293 -194 339 -156
rect 293 -228 299 -194
rect 333 -228 339 -194
rect 293 -266 339 -228
rect 293 -300 299 -266
rect 333 -300 339 -266
rect 293 -338 339 -300
rect 293 -372 299 -338
rect 333 -372 339 -338
rect 293 -413 339 -372
<< end >>
