magic
tech sky130A
magscale 1 2
timestamp 1769409653
<< pwell >>
rect -451 -1647 451 1647
<< psubdiff >>
rect -415 1577 -319 1611
rect 319 1577 415 1611
rect -415 -1577 -381 1577
rect 381 -1577 415 1577
rect -415 -1611 415 -1577
<< psubdiffcont >>
rect -319 1577 319 1611
<< xpolycontact >>
rect -285 1049 285 1481
rect -285 -1481 285 -1049
<< xpolyres >>
rect -285 -1049 285 1049
<< locali >>
rect -415 1577 -319 1611
rect 319 1577 415 1611
rect -415 -1577 -381 1577
rect 381 -1577 415 1577
rect -415 -1611 415 -1577
<< viali >>
rect -269 1066 269 1463
rect -269 -1463 269 -1066
<< metal1 >>
rect -281 1463 281 1469
rect -281 1066 -269 1463
rect 269 1066 281 1463
rect -281 1060 281 1066
rect -281 -1066 281 -1060
rect -281 -1463 -269 -1066
rect 269 -1463 281 -1066
rect -281 -1469 281 -1463
<< labels >>
rlabel psubdiff 0 -1594 0 -1594 0 B
port 1 nsew
rlabel xpolycontact 0 1446 0 1446 0 R1
port 2 nsew
rlabel xpolycontact 0 -1446 0 -1446 0 R2
port 3 nsew
<< properties >>
string FIXED_BBOX -398 -1594 398 1594
string gencell sky130_fd_pr__res_xhigh_po_2p85
string library sky130
string parameters w 2.850 l 10.65 m 1 nx 1 wmin 2.850 lmin 0.50 class resistor rho 2000 val 7.605k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 2.850 guard 1 glc 0 grc 0 gtc 1 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 doports 1
<< end >>
