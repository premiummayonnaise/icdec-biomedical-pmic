magic
tech sky130A
magscale 1 2
timestamp 1769400417
<< error_p >>
rect -29 -92 29 -86
rect -29 -126 -17 -92
rect -29 -132 29 -126
<< nmos >>
rect -15 -54 15 116
<< ndiff >>
rect -73 104 -15 116
rect -73 -42 -61 104
rect -27 -42 -15 104
rect -73 -54 -15 -42
rect 15 104 73 116
rect 15 -42 27 104
rect 61 -42 73 104
rect 15 -54 73 -42
<< ndiffc >>
rect -61 -42 -27 104
rect 27 -42 61 104
<< poly >>
rect -15 116 15 142
rect -15 -76 15 -54
rect -33 -92 33 -76
rect -33 -126 -17 -92
rect 17 -126 33 -92
rect -33 -142 33 -126
<< polycont >>
rect -17 -126 17 -92
<< locali >>
rect -61 104 -27 120
rect -61 -58 -27 -42
rect 27 104 61 120
rect 27 -58 61 -42
rect -33 -126 -17 -92
rect 17 -126 33 -92
<< viali >>
rect -61 -42 -27 104
rect 27 -42 61 104
rect -17 -126 17 -92
<< metal1 >>
rect -67 104 -21 116
rect -67 -42 -61 104
rect -27 -42 -21 104
rect -67 -54 -21 -42
rect 21 104 67 116
rect 21 -42 27 104
rect 61 -42 67 104
rect 21 -54 67 -42
rect -29 -92 29 -86
rect -29 -126 -17 -92
rect 17 -126 29 -92
rect -29 -132 29 -126
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.85 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
