* SPICE3 file created from 1st-stage.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7 a_n29_n444# a_n187_n444# a_29_n532# a_n129_n532#
+ a_129_n444# VSUBS
X0 a_129_n444# a_29_n532# a_n29_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.3775 pd=10.08 as=0.68875 ps=5.04 w=4.75 l=0.5
X1 a_n29_n444# a_n129_n532# a_n187_n444# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=1.3775 ps=10.08 w=4.75 l=0.5
C0 a_n29_n444# a_129_n444# 0.42382f
C1 a_29_n532# a_129_n444# 0.06273f
C2 a_n187_n444# a_n29_n444# 0.42382f
C3 a_29_n532# a_n29_n444# 0.06273f
C4 a_n129_n532# a_n29_n444# 0.06273f
C5 a_n129_n532# a_n187_n444# 0.06273f
C6 a_n129_n532# a_29_n532# 0.05942f
C7 a_129_n444# VSUBS 0.45597f
C8 a_n29_n444# VSUBS 0.10803f
C9 a_n187_n444# VSUBS 0.45597f
C10 a_29_n532# VSUBS 0.25901f
C11 a_n129_n532# VSUBS 0.25901f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_838SN6 a_n187_n506# a_129_n506# a_29_n532# a_n129_n532#
+ a_n29_n506# VSUBS
X0 a_129_n506# a_29_n532# a_n29_n506# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.3775 pd=10.08 as=0.68875 ps=5.04 w=4.75 l=0.5
X1 a_n29_n506# a_n129_n532# a_n187_n506# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.68875 pd=5.04 as=1.3775 ps=10.08 w=4.75 l=0.5
C0 a_n29_n506# a_129_n506# 0.42382f
C1 a_29_n532# a_129_n506# 0.06273f
C2 a_n187_n506# a_n29_n506# 0.42382f
C3 a_29_n532# a_n29_n506# 0.06273f
C4 a_n129_n532# a_n29_n506# 0.06273f
C5 a_n129_n532# a_n187_n506# 0.06273f
C6 a_n129_n532# a_29_n532# 0.05942f
C7 a_129_n506# VSUBS 0.45597f
C8 a_n29_n506# VSUBS 0.10803f
C9 a_n187_n506# VSUBS 0.45597f
C10 a_29_n532# VSUBS 0.25901f
C11 a_n129_n532# VSUBS 0.25901f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_RKS84X m3_n2686_n5200# c1_n2646_n5160# VSUBS
X0 c1_n2646_n5160# m3_n2686_n5200# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X1 c1_n2646_n5160# m3_n2686_n5200# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
C0 m3_n2686_n5200# c1_n2646_n5160# 0.11107p
C1 c1_n2646_n5160# VSUBS 3.9139f
C2 m3_n2686_n5200# VSUBS 25.7614f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DQUD5W a_n953_n781# a_2185_n807# a_n587_n807#
+ a_645_n807# a_29_n807# a_2435_n781# a_n2185_n781# a_1261_n807# a_1569_n807# a_279_n781#
+ a_895_n781# a_n2435_n807# a_n1261_n781# a_1511_n781# a_1819_n781# a_n1569_n781#
+ a_n29_n781# a_n645_n781# a_n1511_n807# a_n279_n807# a_n1819_n807# a_n895_n807# a_337_n807#
+ a_953_n807# a_2127_n781# a_n2493_n781# a_587_n781# a_1877_n807# a_n2127_n807# a_1203_n781#
+ a_n1877_n781# a_n337_n781# a_n1203_n807# VSUBS
X0 a_1511_n781# a_1261_n807# a_1203_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X1 a_n1261_n781# a_n1511_n807# a_n1569_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X2 a_n1877_n781# a_n2127_n807# a_n2185_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X3 a_895_n781# a_645_n807# a_587_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X4 a_n1569_n781# a_n1819_n807# a_n1877_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X5 a_n645_n781# a_n895_n807# a_n953_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X6 a_1819_n781# a_1569_n807# a_1511_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X7 a_n29_n781# a_n279_n807# a_n337_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X8 a_n953_n781# a_n1203_n807# a_n1261_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X9 a_2435_n781# a_2185_n807# a_2127_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=1.25
X10 a_n2185_n781# a_n2435_n807# a_n2493_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=1.25
X11 a_1203_n781# a_953_n807# a_895_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X12 a_587_n781# a_337_n807# a_279_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X13 a_2127_n781# a_1877_n807# a_1819_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X14 a_n337_n781# a_n587_n807# a_n645_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X15 a_279_n781# a_29_n807# a_n29_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
C0 a_29_n807# a_337_n807# 0.05942f
C1 a_n279_n807# a_29_n807# 0.05942f
C2 a_n587_n807# a_n279_n807# 0.05942f
C3 a_n895_n807# a_n587_n807# 0.05942f
C4 a_n1203_n807# a_n895_n807# 0.05942f
C5 a_n1511_n807# a_n1203_n807# 0.05942f
C6 a_n1819_n807# a_n1511_n807# 0.05942f
C7 a_2127_n781# a_2435_n781# 0.34377f
C8 a_n2127_n807# a_n1819_n807# 0.05942f
C9 a_1819_n781# a_2127_n781# 0.34377f
C10 a_n2435_n807# a_n2127_n807# 0.05942f
C11 a_1511_n781# a_1819_n781# 0.34377f
C12 a_1203_n781# a_1511_n781# 0.34377f
C13 a_895_n781# a_1203_n781# 0.34377f
C14 a_587_n781# a_895_n781# 0.34377f
C15 a_279_n781# a_587_n781# 0.34377f
C16 a_n29_n781# a_279_n781# 0.34377f
C17 a_n337_n781# a_n29_n781# 0.34377f
C18 a_2185_n807# a_2435_n781# 0.19032f
C19 a_2185_n807# a_2127_n781# 0.19032f
C20 a_1877_n807# a_2127_n781# 0.19032f
C21 a_n645_n781# a_n337_n781# 0.34377f
C22 a_1877_n807# a_1819_n781# 0.19032f
C23 a_1569_n807# a_1819_n781# 0.19032f
C24 a_n953_n781# a_n645_n781# 0.34377f
C25 a_1569_n807# a_1511_n781# 0.19032f
C26 a_n1261_n781# a_n953_n781# 0.34377f
C27 a_n1569_n781# a_n1261_n781# 0.34377f
C28 a_n1877_n781# a_n1569_n781# 0.34377f
C29 a_1261_n807# a_1511_n781# 0.19032f
C30 a_n2185_n781# a_n1877_n781# 0.34377f
C31 a_1261_n807# a_1203_n781# 0.19032f
C32 a_953_n807# a_1203_n781# 0.19032f
C33 a_n2493_n781# a_n2185_n781# 0.34377f
C34 a_953_n807# a_895_n781# 0.19032f
C35 a_645_n807# a_895_n781# 0.19032f
C36 a_645_n807# a_587_n781# 0.19032f
C37 a_337_n807# a_587_n781# 0.19032f
C38 a_1877_n807# a_2185_n807# 0.05942f
C39 a_337_n807# a_279_n781# 0.19032f
C40 a_29_n807# a_279_n781# 0.19032f
C41 a_1569_n807# a_1877_n807# 0.05942f
C42 a_29_n807# a_n29_n781# 0.19032f
C43 a_n279_n807# a_n29_n781# 0.19032f
C44 a_n279_n807# a_n337_n781# 0.19032f
C45 a_n587_n807# a_n337_n781# 0.19032f
C46 a_n587_n807# a_n645_n781# 0.19032f
C47 a_n895_n807# a_n645_n781# 0.19032f
C48 a_n895_n807# a_n953_n781# 0.19032f
C49 a_n1203_n807# a_n953_n781# 0.19032f
C50 a_1261_n807# a_1569_n807# 0.05942f
C51 a_n1203_n807# a_n1261_n781# 0.19032f
C52 a_n1511_n807# a_n1261_n781# 0.19032f
C53 a_n1511_n807# a_n1569_n781# 0.19032f
C54 a_n1819_n807# a_n1569_n781# 0.19032f
C55 a_n1819_n807# a_n1877_n781# 0.19032f
C56 a_n2127_n807# a_n1877_n781# 0.19032f
C57 a_n2127_n807# a_n2185_n781# 0.19032f
C58 a_953_n807# a_1261_n807# 0.05942f
C59 a_n2435_n807# a_n2185_n781# 0.19032f
C60 a_n2435_n807# a_n2493_n781# 0.19032f
C61 a_645_n807# a_953_n807# 0.05942f
C62 a_337_n807# a_645_n807# 0.05942f
C63 a_2435_n781# VSUBS 0.75893f
C64 a_2127_n781# VSUBS 0.26915f
C65 a_1819_n781# VSUBS 0.26915f
C66 a_1511_n781# VSUBS 0.26915f
C67 a_1203_n781# VSUBS 0.26915f
C68 a_895_n781# VSUBS 0.26915f
C69 a_587_n781# VSUBS 0.26915f
C70 a_279_n781# VSUBS 0.26915f
C71 a_n29_n781# VSUBS 0.26915f
C72 a_n337_n781# VSUBS 0.26915f
C73 a_n645_n781# VSUBS 0.26915f
C74 a_n953_n781# VSUBS 0.26915f
C75 a_n1261_n781# VSUBS 0.26915f
C76 a_n1569_n781# VSUBS 0.26915f
C77 a_n1877_n781# VSUBS 0.26915f
C78 a_n2185_n781# VSUBS 0.26915f
C79 a_n2493_n781# VSUBS 0.75893f
C80 a_2185_n807# VSUBS 0.56406f
C81 a_1877_n807# VSUBS 0.52924f
C82 a_1569_n807# VSUBS 0.52924f
C83 a_1261_n807# VSUBS 0.52924f
C84 a_953_n807# VSUBS 0.52924f
C85 a_645_n807# VSUBS 0.52924f
C86 a_337_n807# VSUBS 0.52924f
C87 a_29_n807# VSUBS 0.52924f
C88 a_n279_n807# VSUBS 0.52924f
C89 a_n587_n807# VSUBS 0.52924f
C90 a_n895_n807# VSUBS 0.52924f
C91 a_n1203_n807# VSUBS 0.52924f
C92 a_n1511_n807# VSUBS 0.52924f
C93 a_n1819_n807# VSUBS 0.52924f
C94 a_n2127_n807# VSUBS 0.52924f
C95 a_n2435_n807# VSUBS 0.56406f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DNNC3W a_29_n807# a_n129_n807# a_n29_n781# a_n187_n781#
+ a_129_n781# VSUBS
X0 a_n29_n781# a_n129_n807# a_n187_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=0.5
X1 a_129_n781# a_29_n807# a_n29_n781# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=0.5
C0 a_n29_n781# a_129_n781# 0.66815f
C1 a_n187_n781# a_n29_n781# 0.66815f
C2 a_29_n807# a_129_n781# 0.0968f
C3 a_29_n807# a_n29_n781# 0.0968f
C4 a_n129_n807# a_n29_n781# 0.0968f
C5 a_n129_n807# a_n187_n781# 0.0968f
C6 a_n129_n807# a_29_n807# 0.05942f
C7 a_129_n781# VSUBS 0.7007f
C8 a_n29_n781# VSUBS 0.1527f
C9 a_n187_n781# VSUBS 0.7007f
C10 a_29_n807# VSUBS 0.25717f
C11 a_n129_n807# VSUBS 0.25717f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_DETAA8 a_587_n964# a_1203_n964# a_337_n1061#
+ a_n279_n1061# a_953_n1061# a_n895_n1061# a_n1203_n1061# a_n337_n964# a_n953_n964#
+ a_29_n1061# w_n1297_n1064# a_279_n964# a_895_n964# a_n1261_n964# a_645_n1061# a_n587_n1061#
+ a_n645_n964# a_n29_n964# VSUBS
X0 a_895_n964# a_645_n1061# a_587_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X1 a_n645_n964# a_n895_n1061# a_n953_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X2 a_n29_n964# a_n279_n1061# a_n337_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X3 a_n953_n964# a_n1203_n1061# a_n1261_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1.25
X4 a_1203_n964# a_953_n1061# a_895_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1.25
X5 a_587_n964# a_337_n1061# a_279_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X6 a_n337_n964# a_n587_n1061# a_n645_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X7 a_279_n964# a_29_n1061# a_n29_n964# w_n1297_n1064# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
C0 a_n279_n1061# a_29_n1061# 0.0619f
C1 a_n587_n1061# a_n279_n1061# 0.0619f
C2 w_n1297_n1064# a_29_n1061# 0.12683f
C3 a_n895_n1061# a_n587_n1061# 0.0619f
C4 w_n1297_n1064# a_n279_n1061# 0.12683f
C5 w_n1297_n1064# a_n587_n1061# 0.12683f
C6 a_n1203_n1061# a_n895_n1061# 0.0619f
C7 w_n1297_n1064# a_n895_n1061# 0.12683f
C8 w_n1297_n1064# a_n1203_n1061# 0.13293f
C9 a_279_n964# a_29_n1061# 0.25181f
C10 a_n29_n964# a_29_n1061# 0.25181f
C11 a_n29_n964# a_n279_n1061# 0.25181f
C12 a_1203_n964# w_n1297_n1064# 0.02956f
C13 a_n337_n964# a_n279_n1061# 0.25181f
C14 a_895_n964# w_n1297_n1064# 0.00517f
C15 a_587_n964# w_n1297_n1064# 0.00517f
C16 a_n337_n964# a_n587_n1061# 0.25181f
C17 a_n645_n964# a_n587_n1061# 0.25181f
C18 a_279_n964# w_n1297_n1064# 0.00517f
C19 a_n29_n964# w_n1297_n1064# 0.00517f
C20 a_n645_n964# a_n895_n1061# 0.25181f
C21 a_895_n964# a_1203_n964# 0.45807f
C22 a_n953_n964# a_n895_n1061# 0.25181f
C23 a_n337_n964# w_n1297_n1064# 0.00517f
C24 a_n645_n964# w_n1297_n1064# 0.00517f
C25 a_n953_n964# a_n1203_n1061# 0.25181f
C26 a_337_n1061# a_29_n1061# 0.0619f
C27 a_n953_n964# w_n1297_n1064# 0.00517f
C28 a_n1261_n964# a_n1203_n1061# 0.25181f
C29 a_587_n964# a_895_n964# 0.45807f
C30 a_n1261_n964# w_n1297_n1064# 0.02956f
C31 a_953_n1061# w_n1297_n1064# 0.13293f
C32 a_279_n964# a_587_n964# 0.45807f
C33 a_645_n1061# w_n1297_n1064# 0.12683f
C34 a_337_n1061# w_n1297_n1064# 0.12683f
C35 a_n29_n964# a_279_n964# 0.45807f
C36 a_n337_n964# a_n29_n964# 0.45807f
C37 a_953_n1061# a_1203_n964# 0.25181f
C38 a_953_n1061# a_895_n964# 0.25181f
C39 a_n645_n964# a_n337_n964# 0.45807f
C40 a_645_n1061# a_895_n964# 0.25181f
C41 a_645_n1061# a_587_n964# 0.25181f
C42 a_n953_n964# a_n645_n964# 0.45807f
C43 a_337_n1061# a_587_n964# 0.25181f
C44 a_337_n1061# a_279_n964# 0.25181f
C45 a_n1261_n964# a_n953_n964# 0.45807f
C46 a_645_n1061# a_953_n1061# 0.0619f
C47 a_337_n1061# a_645_n1061# 0.0619f
C48 a_1203_n964# VSUBS 0.97158f
C49 a_895_n964# VSUBS 0.34405f
C50 a_587_n964# VSUBS 0.34405f
C51 a_279_n964# VSUBS 0.34405f
C52 a_n29_n964# VSUBS 0.34405f
C53 a_n337_n964# VSUBS 0.34405f
C54 a_n645_n964# VSUBS 0.34405f
C55 a_n953_n964# VSUBS 0.34405f
C56 a_n1261_n964# VSUBS 0.97158f
C57 a_953_n1061# VSUBS 0.44026f
C58 a_645_n1061# VSUBS 0.40993f
C59 a_337_n1061# VSUBS 0.40993f
C60 a_29_n1061# VSUBS 0.40993f
C61 a_n279_n1061# VSUBS 0.40993f
C62 a_n587_n1061# VSUBS 0.40993f
C63 a_n895_n1061# VSUBS 0.40993f
C64 a_n1203_n1061# VSUBS 0.44026f
C65 w_n1297_n1064# VSUBS 16.8247f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_686LYQ a_n587_n807# a_587_n719# a_29_n807# a_n337_n719#
+ a_n279_n807# a_337_n807# a_279_n719# a_n29_n719# a_n645_n719# VSUBS
X0 a_n29_n719# a_n279_n807# a_n337_n719# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X1 a_587_n719# a_337_n807# a_279_n719# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=1.25
X2 a_n337_n719# a_n587_n807# a_n645_n719# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=1.25
X3 a_279_n719# a_29_n807# a_n29_n719# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
C0 a_n645_n719# a_n337_n719# 0.34377f
C1 a_n279_n807# a_n337_n719# 0.19032f
C2 a_29_n807# a_337_n807# 0.05942f
C3 a_n587_n807# a_n337_n719# 0.19032f
C4 a_n587_n807# a_n645_n719# 0.19032f
C5 a_n279_n807# a_29_n807# 0.05942f
C6 a_n587_n807# a_n279_n807# 0.05942f
C7 a_n29_n719# a_n337_n719# 0.34377f
C8 a_587_n719# a_337_n807# 0.19032f
C9 a_279_n719# a_337_n807# 0.19032f
C10 a_279_n719# a_29_n807# 0.19032f
C11 a_n29_n719# a_29_n807# 0.19032f
C12 a_n29_n719# a_n279_n807# 0.19032f
C13 a_279_n719# a_587_n719# 0.34377f
C14 a_n29_n719# a_279_n719# 0.34377f
C15 a_587_n719# VSUBS 0.75893f
C16 a_279_n719# VSUBS 0.26915f
C17 a_n29_n719# VSUBS 0.26915f
C18 a_n337_n719# VSUBS 0.26915f
C19 a_n645_n719# VSUBS 0.75893f
C20 a_337_n807# VSUBS 0.56406f
C21 a_29_n807# VSUBS 0.52924f
C22 a_n279_n807# VSUBS 0.52924f
C23 a_n587_n807# VSUBS 0.56406f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y a_29_n1001# w_n223_n1004# a_n129_n1001#
+ a_n29_n904# a_n187_n904# a_129_n904# VSUBS
X0 a_129_n904# a_29_n1001# a_n29_n904# w_n223_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=2.726 pd=19.38 as=1.363 ps=9.69 w=9.4 l=0.5
X1 a_n29_n904# a_n129_n1001# a_n187_n904# w_n223_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=2.726 ps=19.38 w=9.4 l=0.5
C0 a_n129_n1001# a_29_n1001# 0.0619f
C1 w_n223_n1004# a_29_n1001# 0.07336f
C2 w_n223_n1004# a_n129_n1001# 0.07336f
C3 a_129_n904# a_29_n1001# 0.12034f
C4 a_n29_n904# a_29_n1001# 0.12034f
C5 a_129_n904# w_n223_n1004# 0.02814f
C6 a_n29_n904# a_n129_n1001# 0.12034f
C7 a_n29_n904# w_n223_n1004# 0.0052f
C8 a_n187_n904# a_n129_n1001# 0.12034f
C9 a_n187_n904# w_n223_n1004# 0.02814f
C10 a_n29_n904# a_129_n904# 0.83696f
C11 a_n187_n904# a_n29_n904# 0.83696f
C12 a_129_n904# VSUBS 0.84164f
C13 a_n29_n904# VSUBS 0.17835f
C14 a_n187_n904# VSUBS 0.84164f
C15 a_29_n1001# VSUBS 0.18948f
C16 a_n129_n1001# VSUBS 0.18948f
C17 w_n223_n1004# VSUBS 2.7322f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Y7F49Y a_n337_n904# a_n1203_n1001# a_n953_n904#
+ a_2185_n1001# a_29_n1001# w_n2529_n1004# a_n2185_n904# a_2435_n904# a_n2435_n1001#
+ a_279_n904# a_1877_n1001# a_895_n904# a_1261_n1001# a_1511_n904# a_n1261_n904# a_n1569_n904#
+ a_1819_n904# a_645_n1001# a_n587_n1001# a_n1511_n1001# a_n29_n904# a_n645_n904#
+ a_2127_n904# a_n2493_n904# a_n2127_n1001# a_1569_n1001# a_587_n904# a_1203_n904#
+ a_n1877_n904# a_953_n1001# a_337_n1001# a_n279_n1001# a_n895_n1001# a_n1819_n1001#
+ VSUBS
X0 a_n1877_n904# a_n2127_n1001# a_n2185_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X1 a_895_n904# a_645_n1001# a_587_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X2 a_n1569_n904# a_n1819_n1001# a_n1877_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X3 a_n645_n904# a_n895_n1001# a_n953_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X4 a_1819_n904# a_1569_n1001# a_1511_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X5 a_n29_n904# a_n279_n1001# a_n337_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X6 a_n2185_n904# a_n2435_n1001# a_n2493_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=2.726 ps=19.38 w=9.4 l=1.25
X7 a_n953_n904# a_n1203_n1001# a_n1261_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X8 a_1203_n904# a_953_n1001# a_895_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X9 a_2435_n904# a_2185_n1001# a_2127_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=2.726 pd=19.38 as=1.363 ps=9.69 w=9.4 l=1.25
X10 a_587_n904# a_337_n1001# a_279_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X11 a_2127_n904# a_1877_n1001# a_1819_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X12 a_n337_n904# a_n587_n1001# a_n645_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X13 a_279_n904# a_29_n1001# a_n29_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X14 a_n1261_n904# a_n1511_n1001# a_n1569_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X15 a_1511_n904# a_1261_n1001# a_1203_n904# w_n2529_n1004# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
C0 a_n1569_n904# a_n1261_n904# 0.34564f
C1 a_n1877_n904# a_n1569_n904# 0.34564f
C2 a_n2185_n904# a_n1877_n904# 0.34564f
C3 a_n2493_n904# a_n2185_n904# 0.34564f
C4 a_1877_n1001# a_2185_n1001# 0.0619f
C5 a_2127_n904# a_2435_n904# 0.34564f
C6 a_1569_n1001# a_1877_n1001# 0.0619f
C7 a_1819_n904# a_2127_n904# 0.34564f
C8 a_1261_n1001# a_1569_n1001# 0.0619f
C9 a_1511_n904# a_1819_n904# 0.34564f
C10 a_953_n1001# a_1261_n1001# 0.0619f
C11 a_1203_n904# a_1511_n904# 0.34564f
C12 a_645_n1001# a_953_n1001# 0.0619f
C13 a_895_n904# a_1203_n904# 0.34564f
C14 a_587_n904# a_895_n904# 0.34564f
C15 w_n2529_n1004# a_2435_n904# 0.02194f
C16 w_n2529_n1004# a_2127_n904# 0.00341f
C17 a_279_n904# a_587_n904# 0.34564f
C18 w_n2529_n1004# a_1819_n904# 0.00341f
C19 w_n2529_n1004# a_1511_n904# 0.00341f
C20 w_n2529_n1004# a_1203_n904# 0.00341f
C21 a_n29_n904# a_279_n904# 0.34564f
C22 w_n2529_n1004# a_895_n904# 0.00341f
C23 w_n2529_n1004# a_587_n904# 0.00341f
C24 w_n2529_n1004# a_279_n904# 0.00341f
C25 w_n2529_n1004# a_n29_n904# 0.00341f
C26 a_n2435_n1001# a_n2127_n1001# 0.0619f
C27 a_337_n1001# a_587_n904# 0.19111f
C28 a_337_n1001# a_279_n904# 0.19111f
C29 w_n2529_n1004# a_n2127_n1001# 0.12683f
C30 w_n2529_n1004# a_n2435_n1001# 0.13293f
C31 a_29_n1001# a_279_n904# 0.19111f
C32 a_29_n1001# a_n29_n904# 0.19111f
C33 a_n279_n1001# a_n29_n904# 0.19111f
C34 a_337_n1001# w_n2529_n1004# 0.12683f
C35 a_29_n1001# w_n2529_n1004# 0.12683f
C36 a_n279_n1001# w_n2529_n1004# 0.12683f
C37 a_n587_n1001# w_n2529_n1004# 0.12683f
C38 a_29_n1001# a_337_n1001# 0.0619f
C39 a_n895_n1001# w_n2529_n1004# 0.12683f
C40 a_n1203_n1001# w_n2529_n1004# 0.12683f
C41 a_n1819_n1001# a_n2127_n1001# 0.0619f
C42 a_n279_n1001# a_29_n1001# 0.0619f
C43 a_n1511_n1001# w_n2529_n1004# 0.12683f
C44 a_n1819_n1001# w_n2529_n1004# 0.12683f
C45 a_n587_n1001# a_n279_n1001# 0.0619f
C46 a_n895_n1001# a_n587_n1001# 0.0619f
C47 a_2185_n1001# a_2435_n904# 0.19111f
C48 a_n337_n904# a_n29_n904# 0.34564f
C49 a_n1203_n1001# a_n895_n1001# 0.0619f
C50 a_2185_n1001# a_2127_n904# 0.19111f
C51 a_1877_n1001# a_2127_n904# 0.19111f
C52 a_n1511_n1001# a_n1203_n1001# 0.0619f
C53 a_1877_n1001# a_1819_n904# 0.19111f
C54 a_n337_n904# w_n2529_n1004# 0.00341f
C55 a_1569_n1001# a_1819_n904# 0.19111f
C56 a_n645_n904# w_n2529_n1004# 0.00341f
C57 a_n1819_n1001# a_n1511_n1001# 0.0619f
C58 a_n953_n904# w_n2529_n1004# 0.00341f
C59 a_1569_n1001# a_1511_n904# 0.19111f
C60 a_1261_n1001# a_1511_n904# 0.19111f
C61 a_n1877_n904# a_n2127_n1001# 0.19111f
C62 a_n1261_n904# w_n2529_n1004# 0.00341f
C63 a_n2185_n904# a_n2127_n1001# 0.19111f
C64 a_n1569_n904# w_n2529_n1004# 0.00341f
C65 a_n337_n904# a_n279_n1001# 0.19111f
C66 a_1261_n1001# a_1203_n904# 0.19111f
C67 a_n2185_n904# a_n2435_n1001# 0.19111f
C68 a_n337_n904# a_n587_n1001# 0.19111f
C69 a_953_n1001# a_1203_n904# 0.19111f
C70 a_n1877_n904# w_n2529_n1004# 0.00341f
C71 a_953_n1001# a_895_n904# 0.19111f
C72 a_n2185_n904# w_n2529_n1004# 0.00341f
C73 a_n2493_n904# a_n2435_n1001# 0.19111f
C74 a_n645_n904# a_n587_n1001# 0.19111f
C75 a_n645_n904# a_n895_n1001# 0.19111f
C76 a_645_n1001# a_895_n904# 0.19111f
C77 a_n2493_n904# w_n2529_n1004# 0.02194f
C78 a_645_n1001# a_587_n904# 0.19111f
C79 a_n953_n904# a_n895_n1001# 0.19111f
C80 a_2185_n1001# w_n2529_n1004# 0.13293f
C81 a_n953_n904# a_n1203_n1001# 0.19111f
C82 a_1877_n1001# w_n2529_n1004# 0.12683f
C83 a_n1261_n904# a_n1203_n1001# 0.19111f
C84 a_1569_n1001# w_n2529_n1004# 0.12683f
C85 a_n1261_n904# a_n1511_n1001# 0.19111f
C86 a_1261_n1001# w_n2529_n1004# 0.12683f
C87 a_n1569_n904# a_n1511_n1001# 0.19111f
C88 a_953_n1001# w_n2529_n1004# 0.12683f
C89 a_n1569_n904# a_n1819_n1001# 0.19111f
C90 a_645_n1001# w_n2529_n1004# 0.12683f
C91 a_n1877_n904# a_n1819_n1001# 0.19111f
C92 a_645_n1001# a_337_n1001# 0.0619f
C93 a_n645_n904# a_n337_n904# 0.34564f
C94 a_n953_n904# a_n645_n904# 0.34564f
C95 a_n1261_n904# a_n953_n904# 0.34564f
C96 a_2435_n904# VSUBS 0.72996f
C97 a_2127_n904# VSUBS 0.25611f
C98 a_1819_n904# VSUBS 0.25611f
C99 a_1511_n904# VSUBS 0.25611f
C100 a_1203_n904# VSUBS 0.25611f
C101 a_895_n904# VSUBS 0.25611f
C102 a_587_n904# VSUBS 0.25611f
C103 a_279_n904# VSUBS 0.25611f
C104 a_n29_n904# VSUBS 0.25611f
C105 a_n337_n904# VSUBS 0.25611f
C106 a_n645_n904# VSUBS 0.25611f
C107 a_n953_n904# VSUBS 0.25611f
C108 a_n1261_n904# VSUBS 0.25611f
C109 a_n1569_n904# VSUBS 0.25611f
C110 a_n1877_n904# VSUBS 0.25611f
C111 a_n2185_n904# VSUBS 0.25611f
C112 a_n2493_n904# VSUBS 0.72996f
C113 a_2185_n1001# VSUBS 0.44026f
C114 a_1877_n1001# VSUBS 0.40993f
C115 a_1569_n1001# VSUBS 0.40993f
C116 a_1261_n1001# VSUBS 0.40993f
C117 a_953_n1001# VSUBS 0.40993f
C118 a_645_n1001# VSUBS 0.40993f
C119 a_337_n1001# VSUBS 0.40993f
C120 a_29_n1001# VSUBS 0.40993f
C121 a_n279_n1001# VSUBS 0.40993f
C122 a_n587_n1001# VSUBS 0.40993f
C123 a_n895_n1001# VSUBS 0.40993f
C124 a_n1203_n1001# VSUBS 0.40993f
C125 a_n1511_n1001# VSUBS 0.40993f
C126 a_n1819_n1001# VSUBS 0.40993f
C127 a_n2127_n1001# VSUBS 0.40993f
C128 a_n2435_n1001# VSUBS 0.44026f
C129 w_n2529_n1004# VSUBS 30.9853f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AXYYHE w_n303_n564# a_n267_n464# a_29_n561# a_209_n464#
+ a_n29_n464# a_n209_n561# VSUBS
X0 a_n29_n464# a_n209_n561# a_n267_n464# w_n303_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.9
X1 a_209_n464# a_29_n561# a_n29_n464# w_n303_n564# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.9
C0 a_n29_n464# a_209_n464# 0.29682f
C1 a_n267_n464# a_n29_n464# 0.29682f
C2 a_29_n561# a_209_n464# 0.10455f
C3 a_29_n561# a_n29_n464# 0.10455f
C4 w_n303_n564# a_209_n464# 0.01763f
C5 a_n209_n561# a_n29_n464# 0.10455f
C6 a_n209_n561# a_n267_n464# 0.10455f
C7 w_n303_n564# a_n29_n464# 0.00519f
C8 a_n209_n561# a_29_n561# 0.0619f
C9 w_n303_n564# a_n267_n464# 0.01763f
C10 w_n303_n564# a_29_n561# 0.10539f
C11 w_n303_n564# a_n209_n561# 0.10539f
C12 a_209_n464# VSUBS 0.4826f
C13 a_n29_n464# VSUBS 0.15094f
C14 a_n267_n464# VSUBS 0.4826f
C15 a_29_n561# VSUBS 0.32575f
C16 a_n209_n561# VSUBS 0.32575f
C17 w_n303_n564# VSUBS 2.11252f
.ends

.subckt x1st-stage VP VN IBIAS VSS OUT VDD
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_5 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_2 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506#
+ sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# m1_10360_n5790# m1_10360_n5790#
+ li_9700_n5600# VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__cap_mim_m3_1_RKS84X_0 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200#
+ sky130_fd_pr__cap_mim_m3_1_RKS84X_0/c1_n2646_n5160# VSS sky130_fd_pr__cap_mim_m3_1_RKS84X
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_6 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_3 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
XXM24 VSS m1_10880_n8480# m1_10880_n8480# m1_10880_n8480# m1_10880_n8480# m1_10880_n8480#
+ VSS m1_10880_n8480# m1_10880_n8480# VSS VSS m1_10880_n8480# m1_10880_n8480# VSS
+ li_9700_n5600# VSS m1_10880_n8480# li_9700_n5600# m1_10880_n8480# m1_10880_n8480#
+ m1_10880_n8480# m1_10880_n8480# m1_10880_n8480# m1_10880_n8480# VSS m1_10880_n8480#
+ li_9700_n5600# m1_10880_n8480# m1_10880_n8480# m1_10880_n8480# li_9700_n5600# VSS
+ m1_10880_n8480# VSS sky130_fd_pr__nfet_g5v0d10v5_DQUD5W
XXM25 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_DNNC3W
Xsky130_fd_pr__cap_mim_m3_1_RKS84X_1 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200#
+ sky130_fd_pr__cap_mim_m3_1_RKS84X_1/c1_n2646_n5160# VSS sky130_fd_pr__cap_mim_m3_1_RKS84X
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_8 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444#
+ m1_10360_n5790# m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_129_n444#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_4 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506#
+ sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# m1_10360_n5240# m1_10360_n5240#
+ li_9700_n5600# VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__cap_mim_m3_1_RKS84X_2 sky130_fd_pr__cap_mim_m3_1_RKS84X_2/m3_n2686_n5200#
+ sky130_fd_pr__cap_mim_m3_1_RKS84X_2/c1_n2646_n5160# VSS sky130_fd_pr__cap_mim_m3_1_RKS84X
XXM27 XM27/a_587_n964# XM27/a_1203_n964# XM27/a_337_n1061# XM27/a_n279_n1061# XM27/a_953_n1061#
+ XM27/a_n895_n1061# XM27/a_n1203_n1061# VDD VDD XM27/a_29_n1061# VDD VDD VDD XM27/a_n1261_n964#
+ XM27/a_645_n1061# XM27/a_n587_n1061# XM27/a_n645_n964# XM27/a_n29_n964# VSS sky130_fd_pr__pfet_g5v0d10v5_DETAA8
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_9 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_5 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__cap_mim_m3_1_RKS84X_3 sky130_fd_pr__cap_mim_m3_1_RKS84X_3/m3_n2686_n5200#
+ sky130_fd_pr__cap_mim_m3_1_RKS84X_3/c1_n2646_n5160# VSS sky130_fd_pr__cap_mim_m3_1_RKS84X
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_6 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
XXM28 XM28/a_n587_n807# XM28/a_587_n719# XM28/a_29_n807# VSS XM28/a_n279_n807# XM28/a_337_n807#
+ VSS XM28/a_n29_n719# XM28/a_n645_n719# VSS sky130_fd_pr__nfet_g5v0d10v5_686LYQ
Xsky130_fd_pr__nfet_g5v0d10v5_DNNC3W_0 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_DNNC3W
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_8 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_7 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506#
+ sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# m1_10360_n5240# m1_10360_n5240#
+ li_9700_n5600# VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__pfet_g5v0d10v5_DU7D3Y_0 VDD VDD VDD VDD VDD VDD VSS sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_9 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_686LYQ_0 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n587_n807#
+ sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n279_n807# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n645_n719#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_686LYQ
XXM2 VDD m1_10860_n2820# VDD m1_10860_n2820# m1_10860_n2820# VDD VDD m1_10860_n2820#
+ m1_10860_n2820# VDD m1_10860_n2820# VDD m1_10860_n2820# VDD m1_10860_n2820# VDD
+ XM2/a_1819_n904# m1_10860_n2820# m1_10860_n2820# m1_10860_n2820# m1_10860_n2820#
+ XM2/a_n645_n904# VDD m1_10860_n2820# m1_10860_n2820# m1_10860_n2820# XM2/a_587_n904#
+ m1_10860_n2820# XM2/a_n1877_n904# m1_10860_n2820# m1_10860_n2820# m1_10860_n2820#
+ m1_10860_n2820# m1_10860_n2820# VSS sky130_fd_pr__pfet_g5v0d10v5_Y7F49Y
XXM4 VDD VDD VDD VDD VDD VDD VSS sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y
Xsky130_fd_pr__pfet_g5v0d10v5_DETAA8_0 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_587_n964#
+ sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_1203_n964# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_337_n1061#
+ sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n279_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_953_n1061#
+ sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n895_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1203_n1061#
+ VDD VDD sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1261_n964#
+ sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_645_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n587_n1061#
+ sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n645_n964# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964#
+ VSS sky130_fd_pr__pfet_g5v0d10v5_DETAA8
Xsky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n267_n464#
+ sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_29_n561# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464#
+ sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n29_n464# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n209_n561#
+ VSS sky130_fd_pr__pfet_g5v0d10v5_AXYYHE
Xsky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464#
+ sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_29_n561# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_209_n464#
+ sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n29_n464# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561#
+ VSS sky130_fd_pr__pfet_g5v0d10v5_AXYYHE
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_n187_n444#
+ m1_10360_n5240# m1_10360_n5240# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_11 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_0 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_1 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444#
+ m1_10360_n5240# m1_10360_n5240# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_129_n444#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_10 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506#
+ sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# m1_10360_n5790# m1_10360_n5790#
+ li_9700_n5600# VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_3 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_0 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_11 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
Xsky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_n187_n444#
+ m1_10360_n5790# m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7
Xsky130_fd_pr__nfet_g5v0d10v5_838SN6_1 VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_838SN6
C0 XM28/a_29_n807# a_18500_n4990# 0
C1 m1_10860_n2820# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_1203_n964# 0.02398f
C2 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n645_n719# VDD 0.01115f
C3 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# a_8920_n5020# 0.04451f
C4 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_n187_n444# 0.1338f
C5 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444# m2_10300_n4700# 0.11389f
C6 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1203_n1061# 0.02752f
C7 XM28/a_n29_n719# a_18890_n7340# 0.00139f
C8 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# 0
C9 a_17900_n4990# m2_15700_n4700# 0
C10 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# XM27/a_1203_n964# 0.00488f
C11 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# m2_14700_n6200# 0.14275f
C12 XM27/a_645_n1061# VDD 0.86052f
C13 m2_10700_n6800# m3_9300_n10400# 0.00154f
C14 m2_14700_n6200# m3_17100_n10400# 0.00839f
C15 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_209_n464# 0.31561f
C16 XM27/a_n645_n964# m1_10860_n2820# 0
C17 XM27/a_n279_n1061# m1_10860_n2820# 0.00146f
C18 m1_10360_n5790# a_17500_n7340# 0
C19 XM28/a_n279_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n29_n464# 0
C20 m1_10860_n2820# m1_10880_n8480# 0.08148f
C21 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# 0
C22 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# 0
C23 sky130_fd_pr__cap_mim_m3_1_RKS84X_3/m3_n2686_n5200# m3_9300_n10400# 0.13182f
C24 XM28/a_n279_n807# m2_14700_n6200# 0
C25 m1_10360_n5240# m2_14700_n6200# 0.32196f
C26 li_9700_n5600# m2_10700_n6800# 1.20993f
C27 li_9700_n5600# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# 0.00398f
C28 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n29_n464# 0.02806f
C29 IBIAS OUT 0.0352f
C30 XM28/a_29_n807# m3_17100_n10400# 0.04632f
C31 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n587_n807# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n645_n719# -0.02312f
C32 m2_10860_n3800# m2_14300_n4700# 0.55606f
C33 m2_10300_n4700# m2_11700_n4700# 0.02273f
C34 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n645_n719# a_7840_n7320# 0.09425f
C35 VDD m2_10860_n3800# 1.11781f
C36 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# 0
C37 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n29_n464# a_17900_n4990# 0.00427f
C38 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# a_18500_n4990# 0.00145f
C39 li_9700_n5600# XM28/a_n645_n719# 0.00506f
C40 XM28/a_337_n807# VDD 0.01119f
C41 m1_10360_n5790# m2_14700_n6200# 0.25068f
C42 VDD sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444# 0
C43 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444# 0
C44 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n279_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n29_n464# 0.00222f
C45 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1203_n1061# VDD 0.84591f
C46 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_953_n1061# VDD 0.767f
C47 m1_10860_n2820# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# 0.00131f
C48 XM27/a_n645_n964# a_16800_n3320# 0.00188f
C49 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506# m2_14700_n6200# 0.00213f
C50 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# m2_14300_n6800# 0.06259f
C51 m2_14300_n6800# m3_17100_n10400# 0.00154f
C52 VDD a_18890_n7340# 0.01422f
C53 XM28/a_587_n719# VDD 0.01097f
C54 li_9700_n5600# a_8920_n5020# 0
C55 XM27/a_n279_n1061# XM27/a_n29_n964# -0.03407f
C56 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# m1_10360_n5240# -0.02285f
C57 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# XM27/a_29_n1061# 0.02855f
C58 m1_10860_n2820# m2_10300_n4700# 0.51222f
C59 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n279_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n267_n464# 0.00116f
C60 VDD a_19390_n3320# 1.61879f
C61 m1_10360_n5240# m2_14300_n6800# 0.06383f
C62 m1_10860_n2820# a_9230_n7320# 0
C63 li_9700_n5600# m3_9300_n10400# 0.02842f
C64 XM28/a_n587_n807# a_17500_n7340# 0.02643f
C65 XM27/a_645_n1061# XM27/a_587_n964# -0.04158f
C66 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# a_8320_n5020# 0.00147f
C67 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506# m1_10360_n5240# -0.00184f
C68 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# 0.00786f
C69 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444# m1_10360_n5240# -0.01855f
C70 m2_10860_n3800# m2_10300_n6200# 0.4584f
C71 m1_10880_n8480# m2_14700_n6200# 0
C72 XM28/a_n29_n719# a_17500_n7340# 0.00139f
C73 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# a_9950_n3320# 0
C74 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n587_n1061# a_8320_n5020# 0
C75 m1_10360_n5790# m2_14300_n6800# 0.01428f
C76 XM27/a_337_n1061# VDD 0.83963f
C77 XM27/a_n587_n1061# m1_10860_n2820# 0.00606f
C78 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506# m2_14300_n6800# 0.09708f
C79 XM28/a_n279_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# 0
C80 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_n187_n444# m2_10860_n3800# 0.03446f
C81 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# m3_17100_n10400# 0.002f
C82 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506# 0.0024f
C83 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# m1_10360_n5240# 0
C84 a_17900_n4990# a_18500_n4990# 0.02883f
C85 m1_10360_n5240# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444# 0.00698f
C86 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444# a_17900_n4990# 0
C87 XM28/a_n587_n807# m2_14700_n6200# 0.00192f
C88 XM28/a_n29_n719# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n29_n464# 0.00187f
C89 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# a_9230_n7320# 0.02643f
C90 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n267_n464# 0.20182f
C91 a_8320_n5020# a_8920_n5020# 0.02883f
C92 m1_10860_n2820# m2_14300_n4700# 0
C93 m1_10860_n2820# VDD 25.07858f
C94 XM28/a_n279_n807# m3_17100_n10400# 0.06989f
C95 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_1203_n964# a_9950_n3320# 0.08685f
C96 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_129_n444# m1_10360_n5240# 0.0024f
C97 m1_10360_n5240# m3_17100_n10400# 0.24047f
C98 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# m1_10880_n8480# 0
C99 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_29_n561# 0
C100 m1_10860_n2820# XM2/a_587_n904# -0.0062f
C101 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444# -0.02309f
C102 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# a_17900_n4990# 0.04527f
C103 m2_14300_n4700# m2_15700_n4700# 0.02273f
C104 m2_10860_n3800# m2_10700_n6800# 0.57208f
C105 m1_10880_n8480# m2_14300_n6800# 0.05301f
C106 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# a_9230_n7320# 0.09425f
C107 VDD m2_15700_n4700# 0.00966f
C108 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n279_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n267_n464# 0.00227f
C109 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_645_n1061# VDD 0.82988f
C110 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n645_n719# m3_9300_n10400# 0.00257f
C111 XM28/a_n645_n719# sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# 0
C112 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# -0.01775f
C113 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444# m1_10360_n5240# 0.00744f
C114 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# -0.02054f
C115 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_129_n444# -0.00664f
C116 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506# m1_10880_n8480# 0
C117 m1_10360_n5790# m3_17100_n10400# 0.34263f
C118 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444# 0
C119 m1_10860_n2820# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_129_n444# 0.02362f
C120 XM28/a_29_n807# XM28/a_n29_n719# -0.032f
C121 XM27/a_587_n964# a_19390_n3320# 0.00184f
C122 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_29_n561# 0.0073f
C123 VDD a_17500_n7340# 0
C124 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_n187_n444# m2_11700_n4700# 0.14734f
C125 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# XM27/a_n279_n1061# 0.02362f
C126 XM27/a_n279_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# 0.0025f
C127 m1_10860_n2820# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_n187_n444# 0.02918f
C128 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# VDD 0.01039f
C129 m1_10360_n5790# XM28/a_n279_n807# 0
C130 XM28/a_n587_n807# m2_14300_n6800# 0
C131 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n29_n464# a_8920_n5020# 0.00417f
C132 VDD a_16800_n3320# 1.57526f
C133 m1_10360_n5790# m1_10360_n5240# 6.90487f
C134 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# -0.01775f
C135 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444# -0.0206f
C136 m1_10860_n2820# m2_10300_n6200# 0.56833f
C137 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506# m1_10360_n5240# -0.02051f
C138 XM27/a_337_n1061# XM27/a_587_n964# -0.03703f
C139 XM27/a_n29_n964# VDD 0.18761f
C140 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_n187_n444# m2_15700_n4700# 0.14734f
C141 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n29_n464# 0.02336f
C142 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_337_n1061# 0
C143 XM28/a_n645_n719# a_18890_n7340# 0
C144 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# VDD 0.00127f
C145 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444# a_8920_n5020# 0
C146 XM28/a_29_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_29_n561# 0.00718f
C147 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# a_7360_n3320# 0
C148 m1_10860_n2820# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_n187_n444# 0
C149 m1_10880_n8480# m3_17100_n10400# 0.0227f
C150 XM27/a_n1261_n964# m1_10860_n2820# 0.02429f
C151 XM27/a_n895_n1061# m1_10860_n2820# 0.00926f
C152 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# 0
C153 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506# 0.00843f
C154 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# 0.12536f
C155 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561# m2_15700_n4700# 0
C156 XM27/a_1203_n964# VDD 0.85434f
C157 m1_10360_n5240# m1_10880_n8480# 0.02219f
C158 li_9700_n5600# m2_10860_n3800# 1.4509f
C159 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# m2_10300_n6200# 0.00181f
C160 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_29_n561# a_18500_n4990# 0.0269f
C161 XM28/a_n587_n807# m3_17100_n10400# 0.11447f
C162 XM28/a_29_n807# VDD 0.00719f
C163 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444# 0.10715f
C164 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_29_n561# 0.00879f
C165 m1_10860_n2820# m2_10700_n6800# 0.49752f
C166 XM27/a_n279_n1061# a_17900_n4990# 0.00198f
C167 XM28/a_n29_n719# m3_17100_n10400# 0.00742f
C168 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# a_7840_n7320# 0
C169 m1_10360_n5790# m1_10880_n8480# 0.00626f
C170 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_337_n1061# VDD 0.77317f
C171 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# m2_10300_n6200# 0
C172 XM27/a_n1261_n964# a_16800_n3320# 0.08908f
C173 XM27/a_953_n1061# a_19390_n3320# 0.02625f
C174 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506# m1_10880_n8480# 0.00241f
C175 XM27/a_n29_n964# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561# 0.00168f
C176 XM27/a_29_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_29_n561# 0.00906f
C177 XM28/a_n645_n719# m1_10860_n2820# 0
C178 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_29_n561# m2_10300_n4700# 0
C179 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# -0.04469f
C180 XM28/a_n279_n807# XM28/a_n29_n719# -0.02638f
C181 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# a_9230_n7320# 0
C182 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n209_n561# 0
C183 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# 0.15104f
C184 VDD a_18500_n4990# 0.80961f
C185 VDD sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444# 0
C186 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1203_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1261_n964# -0.03554f
C187 m1_10360_n5790# XM28/a_n587_n807# 0
C188 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n29_n464# a_8320_n5020# 0.00427f
C189 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n267_n464# a_8920_n5020# 0.00145f
C190 VDD a_9950_n3320# 1.58528f
C191 m1_10360_n5240# m2_10300_n4700# 0.11936f
C192 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/c1_n2646_n5160# VDD 0.03902f
C193 li_9700_n5600# m2_11700_n4700# 0.33582f
C194 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# 0.00488f
C195 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# m2_10700_n6800# 0
C196 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# a_9230_n7320# 0
C197 XM27/a_29_n1061# VDD 0.79651f
C198 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# VDD 0.58115f
C199 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# 0.25361f
C200 XM28/a_n645_n719# a_17500_n7340# 0.09425f
C201 m1_10860_n2820# m3_9300_n10400# 0.12513f
C202 VDD sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444# 0
C203 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# m2_10300_n6200# 0.0024f
C204 XM27/a_n1203_n1061# m1_10860_n2820# 0.02156f
C205 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# m2_10700_n6800# 0
C206 m1_10360_n5790# a_9230_n7320# 0
C207 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_129_n444# m2_14300_n4700# 0.14523f
C208 VDD m3_17100_n10400# 0.24025f
C209 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_29_n561# 0.18471f
C210 li_9700_n5600# m1_10860_n2820# 1.17961f
C211 XM2/a_n645_n904# VDD 0.12001f
C212 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# a_7360_n3320# 0.00296f
C213 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506# m2_10300_n6200# 0.06818f
C214 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# a_8920_n5020# 0
C215 m1_10860_n2820# XM2/a_n1877_n904# 0.00391f
C216 XM28/a_n645_n719# m2_14700_n6200# 0
C217 XM28/a_n279_n807# VDD 0.0071f
C218 m1_10360_n5240# m2_14300_n4700# 0.005f
C219 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444# m2_14300_n4700# 0.11389f
C220 VDD m1_10360_n5240# 0.04493f
C221 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444# VDD 0
C222 li_9700_n5600# m2_15700_n4700# 0.31472f
C223 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# VDD 0.22168f
C224 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# m3_9300_n10400# 0.10864f
C225 XM27/a_n1203_n1061# a_16800_n3320# 0.02831f
C226 m1_10860_n2820# XM2/a_1819_n904# 0.0046f
C227 a_9230_n7320# m1_10880_n8480# 0
C228 li_9700_n5600# a_17500_n7340# 0.00143f
C229 sky130_fd_pr__cap_mim_m3_1_RKS84X_2/c1_n2646_n5160# m3_17100_n10400# 0.00923f
C230 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# m2_10700_n6800# 0.10888f
C231 XM27/a_29_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561# 0.00293f
C232 m1_10360_n5790# m2_14300_n4700# 0.12654f
C233 m1_10360_n5790# VDD 0.01074f
C234 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n279_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# -0.03407f
C235 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# m3_9300_n10400# 0.13102f
C236 m1_10860_n2820# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_587_n964# 0
C237 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# VDD 0.00664f
C238 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n279_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n209_n561# 0.00514f
C239 VDD a_17900_n4990# 0.72625f
C240 XM27/a_n587_n1061# XM27/a_n645_n964# -0.0326f
C241 m1_10360_n5240# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_129_n444# -0.01853f
C242 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# m2_10300_n6200# 0.14065f
C243 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_1203_n964# VDD 0.80119f
C244 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n267_n464# a_8320_n5020# 0.04527f
C245 VDD a_7360_n3320# 1.62535f
C246 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# XM27/a_587_n964# 0.00488f
C247 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_n187_n444# m1_10360_n5240# -0.01579f
C248 XM27/a_337_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_209_n464# 0.00142f
C249 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506# m2_10700_n6800# 0.12787f
C250 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# 0.02577f
C251 XM28/a_337_n807# XM28/a_587_n719# -0.01788f
C252 XM28/a_337_n807# a_18890_n7340# 0.02643f
C253 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_645_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_587_n964# -0.04158f
C254 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# 0.0051f
C255 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# m2_10860_n3800# 0.02458f
C256 XM28/a_n645_n719# m2_14300_n6800# 0
C257 m1_10360_n5240# m2_10300_n6200# 0.32247f
C258 XM27/a_n645_n964# VDD 0.221f
C259 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# m2_10300_n6200# 0.10931f
C260 XM27/a_n279_n1061# VDD 0.82211f
C261 li_9700_n5600# m2_14700_n6200# 0.71432f
C262 XM27/a_953_n1061# XM27/a_1203_n964# -0.02548f
C263 XM28/a_n279_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561# 0.00761f
C264 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n645_n964# a_7360_n3320# 0.00188f
C265 XM2/a_1819_n904# a_16800_n3320# 0
C266 m2_10860_n3800# m2_11700_n4700# 0.55606f
C267 VDD m1_10880_n8480# 0.01299f
C268 XM28/a_587_n719# a_18890_n7340# 0.09425f
C269 m1_10360_n5240# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_n187_n444# 0.00234f
C270 XM28/a_n29_n719# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_29_n561# 0
C271 m1_10360_n5790# m2_10300_n6200# 0.25068f
C272 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n209_n561# 0.17929f
C273 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# m2_10300_n6200# 0
C274 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# -0.021f
C275 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# m2_10700_n6800# 0.04151f
C276 m1_10860_n2820# sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# 0.00819f
C277 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_n187_n444# -0.00384f
C278 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561# a_17900_n4990# 0.02831f
C279 XM28/a_n587_n807# VDD 0.01052f
C280 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# 0.12649f
C281 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n279_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n209_n561# 0.01101f
C282 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# VDD 0.86494f
C283 m1_10860_n2820# m2_10860_n3800# 3.97566f
C284 XM28/a_n645_n719# sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# 0
C285 XM28/a_n645_n719# m3_17100_n10400# 0.13475f
C286 XM28/a_n29_n719# VDD 0.00124f
C287 m1_10360_n5240# m2_10700_n6800# 0.06256f
C288 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# m2_10700_n6800# 0.00197f
C289 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# m1_10360_n5240# 0
C290 li_9700_n5600# m2_14300_n6800# 1.21451f
C291 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/c1_n2646_n5160# VDD 0.05954f
C292 m1_10860_n2820# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444# 0.00799f
C293 m1_10860_n2820# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_953_n1061# 0.02067f
C294 sky130_fd_pr__cap_mim_m3_1_RKS84X_2/m3_n2686_n5200# m3_17100_n10400# 0.12057f
C295 XM27/a_n279_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561# 0.00459f
C296 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506# 0.1326f
C297 m2_10860_n3800# m2_15700_n4700# 0.01364f
C298 m1_10880_n8480# m2_10300_n6200# 0
C299 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444# 0.12564f
C300 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# VDD 0.63662f
C301 VDD m2_10300_n4700# 0.00844f
C302 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# a_17500_n7340# 0
C303 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n279_n807# VDD 0.00724f
C304 VDD a_9230_n7320# 0.00137f
C305 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_29_n561# a_8920_n5020# 0.0269f
C306 XM27/a_n895_n1061# XM27/a_n645_n964# -0.04626f
C307 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# XM27/a_953_n1061# 0.02932f
C308 m1_10360_n5790# m2_10700_n6800# 0.01484f
C309 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n209_n561# 0.00321f
C310 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# m3_9300_n10400# 0.0021f
C311 XM2/a_n1877_n904# a_9950_n3320# 0
C312 li_9700_n5600# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# 0.00382f
C313 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_29_n561# 0.18888f
C314 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n645_n964# 0.00488f
C315 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n279_n1061# 0.02778f
C316 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_337_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_587_n964# -0.02272f
C317 m1_10360_n5790# XM28/a_n645_n719# 0
C318 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444# 0.1267f
C319 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_129_n444# m2_10300_n4700# 0.14523f
C320 XM27/a_n587_n1061# VDD 0.81793f
C321 m1_10860_n2820# m2_11700_n4700# 0
C322 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# m2_14700_n6200# 0.12214f
C323 m1_10360_n5240# m3_9300_n10400# 0.24047f
C324 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# m3_9300_n10400# 0.00401f
C325 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# 0.13202f
C326 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# li_9700_n5600# 0.15042f
C327 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_129_n444# 0.15232f
C328 li_9700_n5600# m3_17100_n10400# 0.02785f
C329 XM28/a_587_n719# a_17500_n7340# 0
C330 a_17500_n7340# a_18890_n7340# 0.01812f
C331 XM28/a_29_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_209_n464# 0
C332 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_587_n964# a_9950_n3320# 0.00184f
C333 m2_10860_n3800# m2_14700_n6200# 0.4584f
C334 m1_10880_n8480# m2_10700_n6800# 0.05125f
C335 a_7840_n7320# a_9230_n7320# 0.01812f
C336 a_9230_n7320# m2_10300_n6200# 0.00145f
C337 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n279_n807# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# -0.02638f
C338 m1_10360_n5790# m3_9300_n10400# 0.34346f
C339 li_9700_n5600# m1_10360_n5240# 7.49028f
C340 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# a_9230_n7320# 0.00139f
C341 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# li_9700_n5600# 0.10695f
C342 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444# 0.10827f
C343 XM2/a_587_n904# VDD 0.14329f
C344 VP VN 0.0352f
C345 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# m3_9300_n10400# 0.07275f
C346 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n645_n964# VDD 0.18806f
C347 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n279_n1061# VDD 0.81753f
C348 XM27/a_n29_n964# a_19390_n3320# 0
C349 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_209_n464# a_18500_n4990# 0.04451f
C350 sky130_fd_pr__cap_mim_m3_1_RKS84X_3/c1_n2646_n5160# VDD 0.00638f
C351 VDD sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_129_n444# 0
C352 m1_10360_n5790# li_9700_n5600# 7.23542f
C353 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# 0.00397f
C354 m1_10860_n2820# m2_15700_n4700# 0.51469f
C355 m1_10860_n2820# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_645_n1061# 0.00929f
C356 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# m2_14700_n6200# 0.04519f
C357 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506# 0.10819f
C358 li_9700_n5600# a_17900_n4990# 0
C359 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# m2_14300_n6800# 0.00222f
C360 sky130_fd_pr__cap_mim_m3_1_RKS84X_2/c1_n2646_n5160# VDD 0.00588f
C361 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# m2_10860_n3800# 0.00903f
C362 XM28/a_n587_n807# XM28/a_n645_n719# -0.02312f
C363 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n587_n807# VDD 0.01127f
C364 VDD a_7840_n7320# 0.01447f
C365 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# XM27/a_645_n1061# 0.02649f
C366 m1_10860_n2820# a_17500_n7340# 0
C367 m2_10860_n3800# m2_14300_n6800# 0.57208f
C368 m1_10880_n8480# m3_9300_n10400# 0.02215f
C369 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# m2_10300_n4700# 0
C370 XM27/a_1203_n964# a_19390_n3320# 0.08685f
C371 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# VDD 0
C372 a_9230_n7320# m2_10700_n6800# 0
C373 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506# m2_10860_n3800# 0.02794f
C374 m1_10860_n2820# a_16800_n3320# 0.00665f
C375 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561# 0.18569f
C376 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n587_n1061# 0.02803f
C377 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# a_8920_n5020# 0.00147f
C378 XM27/a_n1261_n964# VDD 0.81114f
C379 XM27/a_n895_n1061# VDD 0.8497f
C380 li_9700_n5600# m1_10880_n8480# 5.19572f
C381 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# m1_10860_n2820# 0
C382 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1261_n964# a_7360_n3320# 0.08908f
C383 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_953_n1061# a_9950_n3320# 0.02625f
C384 XM27/a_587_n964# VDD 0.22153f
C385 m1_10860_n2820# m2_14700_n6200# 0.56833f
C386 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# m2_14300_n6800# 0.12595f
C387 a_8920_n5020# m2_10300_n4700# 0
C388 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444# m2_10860_n3800# 0.01111f
C389 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# m3_17100_n10400# 0.00378f
C390 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n587_n807# a_7840_n7320# 0.02643f
C391 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_129_n444# m2_10860_n3800# 0.02901f
C392 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# a_7840_n7320# 0.00139f
C393 VDD sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# 0.31883f
C394 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n279_n807# m3_9300_n10400# 0.04772f
C395 a_9230_n7320# m3_9300_n10400# 0.02466f
C396 XM28/a_337_n807# m3_17100_n10400# 0.03269f
C397 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n29_n464# 0.00106f
C398 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n587_n1061# VDD 0.82209f
C399 XM27/a_337_n1061# a_18500_n4990# 0.00198f
C400 XM27/a_n29_n964# a_16800_n3320# 0
C401 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# a_19390_n3320# 0.00291f
C402 a_17500_n7340# m2_14700_n6200# 0.00152f
C403 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_209_n464# a_17900_n4990# 0.00147f
C404 XM28/a_n645_n719# VDD 0.00127f
C405 sky130_fd_pr__cap_mim_m3_1_RKS84X_3/m3_n2686_n5200# VDD 0.32519f
C406 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# -0.0286f
C407 m1_10360_n5240# m2_10860_n3800# 1.19867f
C408 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444# m2_10860_n3800# 0.01044f
C409 li_9700_n5600# m2_10300_n4700# 0.31451f
C410 m1_10860_n2820# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_337_n1061# 0.00555f
C411 a_18890_n7340# m3_17100_n10400# 0.00349f
C412 XM28/a_587_n719# m3_17100_n10400# 0.00261f
C413 li_9700_n5600# a_9230_n7320# 0.00143f
C414 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# -0.02054f
C415 m1_10360_n5240# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444# -0.01579f
C416 sky130_fd_pr__cap_mim_m3_1_RKS84X_2/m3_n2686_n5200# VDD 0.31878f
C417 m1_10860_n2820# m2_14300_n6800# 0.49752f
C418 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n587_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n645_n964# -0.0326f
C419 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n29_n464# 0.00116f
C420 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444# m2_11700_n4700# 0.12672f
C421 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n209_n561# a_8320_n5020# 0.02831f
C422 VDD a_8920_n5020# 0.75851f
C423 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# XM27/a_337_n1061# 0.02726f
C424 m1_10360_n5790# m2_10860_n3800# 1.6602f
C425 m1_10860_n2820# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444# 0.00866f
C426 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506# m2_10860_n3800# 0.00834f
C427 m1_10860_n2820# a_9950_n3320# 0.00677f
C428 m2_10300_n6200# m2_10700_n6800# 0.19444f
C429 VDD m3_9300_n10400# 0.24031f
C430 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1261_n964# 0.00488f
C431 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n895_n1061# 0.02829f
C432 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# m1_10360_n5240# -0.00464f
C433 XM27/a_n1203_n1061# VDD 0.74616f
C434 XM27/a_953_n1061# VDD 0.7994f
C435 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444# m2_15700_n4700# 0.12672f
C436 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_953_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_1203_n964# -0.02548f
C437 a_17500_n7340# m2_14300_n6800# 0
C438 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1203_n1061# a_7360_n3320# 0.02831f
C439 m1_10360_n5240# m2_11700_n4700# 0.00667f
C440 m1_10860_n2820# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444# 0.0027f
C441 li_9700_n5600# m2_14300_n4700# 0.33561f
C442 li_9700_n5600# VDD 0.10716f
C443 m1_10360_n5790# sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# 0.00246f
C444 sky130_fd_pr__cap_mim_m3_1_RKS84X_3/c1_n2646_n5160# m3_9300_n10400# 0.01044f
C445 m1_10880_n8480# m2_10860_n3800# 0.08357f
C446 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n279_n807# a_8320_n5020# 0
C447 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# m2_15700_n4700# 0
C448 m1_10860_n2820# sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# 0.02465f
C449 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# m1_10860_n2820# 0.02117f
C450 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_129_n444# m1_10860_n2820# 0
C451 m1_10860_n2820# m3_17100_n10400# 0.12513f
C452 XM2/a_n1877_n904# VDD 0.12135f
C453 m1_10860_n2820# XM2/a_n645_n904# 0.00442f
C454 m1_10360_n5790# m2_11700_n4700# 0.12434f
C455 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n645_n719# a_9230_n7320# 0
C456 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n587_n807# m3_9300_n10400# 0.03062f
C457 a_7840_n7320# m3_9300_n10400# 0.00345f
C458 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n29_n464# a_18500_n4990# 0.00417f
C459 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_129_n444# 0.15173f
C460 m2_14700_n6200# m2_14300_n6800# 0.19444f
C461 m2_10300_n6200# m3_9300_n10400# 0.00839f
C462 m1_10860_n2820# m1_10360_n5240# 1.42928f
C463 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# m1_10860_n2820# 0.00758f
C464 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444# m1_10860_n2820# 0.00272f
C465 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1261_n964# VDD 0.91243f
C466 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n895_n1061# VDD 0.81395f
C467 XM2/a_1819_n904# VDD 0.12027f
C468 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# m3_9300_n10400# 0.00726f
C469 li_9700_n5600# sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_n187_n444# 0.13324f
C470 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_587_n964# VDD 0.18868f
C471 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# a_17500_n7340# 0
C472 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# m1_10880_n8480# 0
C473 a_17500_n7340# m3_17100_n10400# 0.0247f
C474 XM27/a_29_n1061# XM27/a_n29_n964# -0.02972f
C475 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# XM27/a_n29_n964# 0.00488f
C476 m1_10360_n5240# m2_15700_n4700# 0.11934f
C477 XM27/a_29_n1061# sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n29_n464# 0.0025f
C478 li_9700_n5600# m2_10300_n6200# 0.71756f
C479 m1_10360_n5790# m1_10860_n2820# 0.84328f
C480 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n895_n1061# sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n645_n964# -0.03115f
C481 VDD a_8320_n5020# 0.77339f
C482 XM27/a_n1203_n1061# XM27/a_n1261_n964# -0.02136f
C483 m2_10860_n3800# m2_10300_n4700# 0.01818f
C484 OUT VSS 0.15979f
C485 IBIAS VSS 0.15979f
C486 VN VSS 0.15979f
C487 VP VSS 0.15979f
C488 m3_17100_n10400# VSS 3.18057f **FLOATING
C489 m3_9300_n10400# VSS 3.19623f **FLOATING
C490 m2_14300_n6800# VSS 1.69656f **FLOATING
C491 m2_10700_n6800# VSS 1.6971f **FLOATING
C492 m2_14700_n6200# VSS 1.67582f **FLOATING
C493 m2_10300_n6200# VSS 1.66931f **FLOATING
C494 m2_15700_n4700# VSS 0.84866f **FLOATING
C495 m2_14300_n4700# VSS 0.80379f **FLOATING
C496 m2_11700_n4700# VSS 0.80961f **FLOATING
C497 m2_10300_n4700# VSS 0.84137f **FLOATING
C498 m2_10860_n3800# VSS 4.8071f **FLOATING
C499 m1_10880_n8480# VSS 27.11354f
C500 a_18890_n7340# VSS 1.46233f **FLOATING
C501 a_17500_n7340# VSS 1.49112f **FLOATING
C502 a_18500_n4990# VSS 0.01533f **FLOATING
C503 a_17900_n4990# VSS 0.06911f **FLOATING
C504 a_9230_n7320# VSS 1.46962f **FLOATING
C505 a_7840_n7320# VSS 1.48112f **FLOATING
C506 a_8920_n5020# VSS 0.07896f **FLOATING
C507 a_8320_n5020# VSS 0.01465f **FLOATING
C508 a_19390_n3320# VSS 0.08083f **FLOATING
C509 a_16800_n3320# VSS 0.04815f **FLOATING
C510 a_9950_n3320# VSS 0.04836f **FLOATING
C511 a_7360_n3320# VSS 0.08311f **FLOATING
C512 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_129_n444# VSS 1.05043f
C513 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4/a_n187_n444# VSS 1.06835f
C514 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_129_n506# VSS 1.05107f
C515 sky130_fd_pr__nfet_g5v0d10v5_838SN6_10/a_n187_n506# VSS 1.06815f
C516 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_129_n444# VSS 1.04645f
C517 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2/a_n187_n444# VSS 1.07232f
C518 m1_10360_n5240# VSS 4.58803f
C519 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_129_n444# VSS 1.05043f
C520 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10/a_n187_n444# VSS 1.06835f
C521 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_209_n464# VSS 0.48356f
C522 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n29_n464# VSS 0.15151f
C523 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n267_n464# VSS 0.53681f
C524 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_29_n561# VSS 0.33043f
C525 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1/a_n209_n561# VSS 0.33311f
C526 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_209_n464# VSS 0.54505f
C527 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n29_n464# VSS 0.1516f
C528 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n267_n464# VSS 0.48326f
C529 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_29_n561# VSS 0.33483f
C530 sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0/a_n209_n561# VSS 0.33125f
C531 VDD VSS 0.20106p
C532 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_1203_n964# VSS 0.97448f
C533 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_587_n964# VSS 0.34423f
C534 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n29_n964# VSS 0.34405f
C535 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n645_n964# VSS 0.34405f
C536 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1261_n964# VSS 0.97158f
C537 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_953_n1061# VSS 0.45542f
C538 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_645_n1061# VSS 0.42534f
C539 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_337_n1061# VSS 0.40993f
C540 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_29_n1061# VSS 0.40993f
C541 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n279_n1061# VSS 0.40993f
C542 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n587_n1061# VSS 0.40993f
C543 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n895_n1061# VSS 0.40993f
C544 sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0/a_n1203_n1061# VSS 0.44026f
C545 XM2/a_1819_n904# VSS 0.25611f
C546 XM2/a_587_n904# VSS 0.25611f
C547 XM2/a_n645_n904# VSS 0.25611f
C548 XM2/a_n1877_n904# VSS 0.25611f
C549 m1_10860_n2820# VSS 5.9758f
C550 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_587_n719# VSS 1.33888f
C551 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n29_n719# VSS 0.41169f
C552 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n645_n719# VSS 1.29873f
C553 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_337_n807# VSS 1.15875f
C554 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_29_n807# VSS 1.07616f
C555 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n279_n807# VSS 1.10251f
C556 sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0/a_n587_n807# VSS 1.13254f
C557 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_129_n506# VSS 1.04625f
C558 sky130_fd_pr__nfet_g5v0d10v5_838SN6_7/a_n187_n506# VSS 1.07302f
C559 XM28/a_587_n719# VSS 1.25703f
C560 XM28/a_n29_n719# VSS 0.34908f
C561 XM28/a_n645_n719# VSS 1.35742f
C562 XM28/a_337_n807# VSS 1.12003f
C563 XM28/a_29_n807# VSS 1.14281f
C564 XM28/a_n279_n807# VSS 0.84888f
C565 XM28/a_n587_n807# VSS 1.14859f
C566 sky130_fd_pr__cap_mim_m3_1_RKS84X_3/c1_n2646_n5160# VSS 3.96799f
C567 sky130_fd_pr__cap_mim_m3_1_RKS84X_3/m3_n2686_n5200# VSS 26.11986f
C568 XM27/a_1203_n964# VSS 0.97158f
C569 XM27/a_587_n964# VSS 0.34405f
C570 XM27/a_n29_n964# VSS 0.34405f
C571 XM27/a_n645_n964# VSS 0.34502f
C572 XM27/a_n1261_n964# VSS 0.97452f
C573 XM27/a_953_n1061# VSS 0.44026f
C574 XM27/a_645_n1061# VSS 0.40993f
C575 XM27/a_337_n1061# VSS 0.40993f
C576 XM27/a_29_n1061# VSS 0.40993f
C577 XM27/a_n279_n1061# VSS 0.40993f
C578 XM27/a_n587_n1061# VSS 0.40993f
C579 XM27/a_n895_n1061# VSS 0.42534f
C580 XM27/a_n1203_n1061# VSS 0.45503f
C581 sky130_fd_pr__cap_mim_m3_1_RKS84X_2/c1_n2646_n5160# VSS 3.95199f
C582 sky130_fd_pr__cap_mim_m3_1_RKS84X_2/m3_n2686_n5200# VSS 26.09601f
C583 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_129_n506# VSS 1.05285f
C584 sky130_fd_pr__nfet_g5v0d10v5_838SN6_4/a_n187_n506# VSS 1.06815f
C585 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_129_n444# VSS 1.04645f
C586 sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7/a_n187_n444# VSS 1.07232f
C587 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/c1_n2646_n5160# VSS 3.9139f
C588 sky130_fd_pr__cap_mim_m3_1_RKS84X_1/m3_n2686_n5200# VSS 25.7614f
C589 li_9700_n5600# VSS 28.52663f
C590 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/c1_n2646_n5160# VSS 3.9139f
C591 sky130_fd_pr__cap_mim_m3_1_RKS84X_0/m3_n2686_n5200# VSS 25.7614f
C592 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_129_n506# VSS 1.0464f
C593 sky130_fd_pr__nfet_g5v0d10v5_838SN6_2/a_n187_n506# VSS 1.07167f
C594 m1_10360_n5790# VSS 4.66799f
.ends

