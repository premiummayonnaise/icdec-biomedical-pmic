magic
tech sky130A
timestamp 1769135993
<< pwell >>
rect -123 -275 123 275
<< nmos >>
rect -25 -170 25 170
<< ndiff >>
rect -54 164 -25 170
rect -54 -164 -48 164
rect -31 -164 -25 164
rect -54 -170 -25 -164
rect 25 164 54 170
rect 25 -164 31 164
rect 48 -164 54 164
rect 25 -170 54 -164
<< ndiffc >>
rect -48 -164 -31 164
rect 31 -164 48 164
<< psubdiff >>
rect -105 240 -57 257
rect 57 240 105 257
rect -105 209 -88 240
rect 88 209 105 240
rect -105 -240 -88 -209
rect 88 -240 105 -209
rect -105 -257 -57 -240
rect 57 -257 105 -240
<< psubdiffcont >>
rect -57 240 57 257
rect -105 -209 -88 209
rect 88 -209 105 209
rect -57 -257 57 -240
<< poly >>
rect -25 206 25 214
rect -25 189 -17 206
rect 17 189 25 206
rect -25 170 25 189
rect -25 -189 25 -170
rect -25 -206 -17 -189
rect 17 -206 25 -189
rect -25 -214 25 -206
<< polycont >>
rect -17 189 17 206
rect -17 -206 17 -189
<< locali >>
rect -105 240 -57 257
rect 57 240 105 257
rect -105 209 -88 240
rect 88 209 105 240
rect -25 189 -17 206
rect 17 189 25 206
rect -48 164 -31 172
rect -48 -172 -31 -164
rect 31 164 48 172
rect 31 -172 48 -164
rect -25 -206 -17 -189
rect 17 -206 25 -189
rect -105 -240 -88 -209
rect 88 -240 105 -209
rect -105 -257 -57 -240
rect 57 -257 105 -240
<< viali >>
rect -17 189 17 206
rect -48 -164 -31 164
rect 31 -164 48 164
rect -17 -206 17 -189
<< metal1 >>
rect -23 206 23 209
rect -23 189 -17 206
rect 17 189 23 206
rect -23 186 23 189
rect -51 164 -28 170
rect -51 -164 -48 164
rect -31 -164 -28 164
rect -51 -170 -28 -164
rect 28 164 51 170
rect 28 -164 31 164
rect 48 -164 51 164
rect 28 -170 51 -164
rect -23 -189 23 -186
rect -23 -206 -17 -189
rect 17 -206 23 -189
rect -23 -209 23 -206
<< properties >>
string FIXED_BBOX -96 -248 96 248
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.4 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
