magic
tech sky130A
magscale 1 2
timestamp 1769406237
<< nwell >>
rect -4993 -408 4993 442
<< pmos >>
rect -4899 -308 -4649 380
rect -4591 -308 -4341 380
rect -4283 -308 -4033 380
rect -3975 -308 -3725 380
rect -3667 -308 -3417 380
rect -3359 -308 -3109 380
rect -3051 -308 -2801 380
rect -2743 -308 -2493 380
rect -2435 -308 -2185 380
rect -2127 -308 -1877 380
rect -1819 -308 -1569 380
rect -1511 -308 -1261 380
rect -1203 -308 -953 380
rect -895 -308 -645 380
rect -587 -308 -337 380
rect -279 -308 -29 380
rect 29 -308 279 380
rect 337 -308 587 380
rect 645 -308 895 380
rect 953 -308 1203 380
rect 1261 -308 1511 380
rect 1569 -308 1819 380
rect 1877 -308 2127 380
rect 2185 -308 2435 380
rect 2493 -308 2743 380
rect 2801 -308 3051 380
rect 3109 -308 3359 380
rect 3417 -308 3667 380
rect 3725 -308 3975 380
rect 4033 -308 4283 380
rect 4341 -308 4591 380
rect 4649 -308 4899 380
<< pdiff >>
rect -4957 368 -4899 380
rect -4957 -296 -4945 368
rect -4911 -296 -4899 368
rect -4957 -308 -4899 -296
rect -4649 368 -4591 380
rect -4649 -296 -4637 368
rect -4603 -296 -4591 368
rect -4649 -308 -4591 -296
rect -4341 368 -4283 380
rect -4341 -296 -4329 368
rect -4295 -296 -4283 368
rect -4341 -308 -4283 -296
rect -4033 368 -3975 380
rect -4033 -296 -4021 368
rect -3987 -296 -3975 368
rect -4033 -308 -3975 -296
rect -3725 368 -3667 380
rect -3725 -296 -3713 368
rect -3679 -296 -3667 368
rect -3725 -308 -3667 -296
rect -3417 368 -3359 380
rect -3417 -296 -3405 368
rect -3371 -296 -3359 368
rect -3417 -308 -3359 -296
rect -3109 368 -3051 380
rect -3109 -296 -3097 368
rect -3063 -296 -3051 368
rect -3109 -308 -3051 -296
rect -2801 368 -2743 380
rect -2801 -296 -2789 368
rect -2755 -296 -2743 368
rect -2801 -308 -2743 -296
rect -2493 368 -2435 380
rect -2493 -296 -2481 368
rect -2447 -296 -2435 368
rect -2493 -308 -2435 -296
rect -2185 368 -2127 380
rect -2185 -296 -2173 368
rect -2139 -296 -2127 368
rect -2185 -308 -2127 -296
rect -1877 368 -1819 380
rect -1877 -296 -1865 368
rect -1831 -296 -1819 368
rect -1877 -308 -1819 -296
rect -1569 368 -1511 380
rect -1569 -296 -1557 368
rect -1523 -296 -1511 368
rect -1569 -308 -1511 -296
rect -1261 368 -1203 380
rect -1261 -296 -1249 368
rect -1215 -296 -1203 368
rect -1261 -308 -1203 -296
rect -953 368 -895 380
rect -953 -296 -941 368
rect -907 -296 -895 368
rect -953 -308 -895 -296
rect -645 368 -587 380
rect -645 -296 -633 368
rect -599 -296 -587 368
rect -645 -308 -587 -296
rect -337 368 -279 380
rect -337 -296 -325 368
rect -291 -296 -279 368
rect -337 -308 -279 -296
rect -29 368 29 380
rect -29 -296 -17 368
rect 17 -296 29 368
rect -29 -308 29 -296
rect 279 368 337 380
rect 279 -296 291 368
rect 325 -296 337 368
rect 279 -308 337 -296
rect 587 368 645 380
rect 587 -296 599 368
rect 633 -296 645 368
rect 587 -308 645 -296
rect 895 368 953 380
rect 895 -296 907 368
rect 941 -296 953 368
rect 895 -308 953 -296
rect 1203 368 1261 380
rect 1203 -296 1215 368
rect 1249 -296 1261 368
rect 1203 -308 1261 -296
rect 1511 368 1569 380
rect 1511 -296 1523 368
rect 1557 -296 1569 368
rect 1511 -308 1569 -296
rect 1819 368 1877 380
rect 1819 -296 1831 368
rect 1865 -296 1877 368
rect 1819 -308 1877 -296
rect 2127 368 2185 380
rect 2127 -296 2139 368
rect 2173 -296 2185 368
rect 2127 -308 2185 -296
rect 2435 368 2493 380
rect 2435 -296 2447 368
rect 2481 -296 2493 368
rect 2435 -308 2493 -296
rect 2743 368 2801 380
rect 2743 -296 2755 368
rect 2789 -296 2801 368
rect 2743 -308 2801 -296
rect 3051 368 3109 380
rect 3051 -296 3063 368
rect 3097 -296 3109 368
rect 3051 -308 3109 -296
rect 3359 368 3417 380
rect 3359 -296 3371 368
rect 3405 -296 3417 368
rect 3359 -308 3417 -296
rect 3667 368 3725 380
rect 3667 -296 3679 368
rect 3713 -296 3725 368
rect 3667 -308 3725 -296
rect 3975 368 4033 380
rect 3975 -296 3987 368
rect 4021 -296 4033 368
rect 3975 -308 4033 -296
rect 4283 368 4341 380
rect 4283 -296 4295 368
rect 4329 -296 4341 368
rect 4283 -308 4341 -296
rect 4591 368 4649 380
rect 4591 -296 4603 368
rect 4637 -296 4649 368
rect 4591 -308 4649 -296
rect 4899 368 4957 380
rect 4899 -296 4911 368
rect 4945 -296 4957 368
rect 4899 -308 4957 -296
<< pdiffc >>
rect -4945 -296 -4911 368
rect -4637 -296 -4603 368
rect -4329 -296 -4295 368
rect -4021 -296 -3987 368
rect -3713 -296 -3679 368
rect -3405 -296 -3371 368
rect -3097 -296 -3063 368
rect -2789 -296 -2755 368
rect -2481 -296 -2447 368
rect -2173 -296 -2139 368
rect -1865 -296 -1831 368
rect -1557 -296 -1523 368
rect -1249 -296 -1215 368
rect -941 -296 -907 368
rect -633 -296 -599 368
rect -325 -296 -291 368
rect -17 -296 17 368
rect 291 -296 325 368
rect 599 -296 633 368
rect 907 -296 941 368
rect 1215 -296 1249 368
rect 1523 -296 1557 368
rect 1831 -296 1865 368
rect 2139 -296 2173 368
rect 2447 -296 2481 368
rect 2755 -296 2789 368
rect 3063 -296 3097 368
rect 3371 -296 3405 368
rect 3679 -296 3713 368
rect 3987 -296 4021 368
rect 4295 -296 4329 368
rect 4603 -296 4637 368
rect 4911 -296 4945 368
<< poly >>
rect -4899 380 -4649 406
rect -4591 380 -4341 406
rect -4283 380 -4033 406
rect -3975 380 -3725 406
rect -3667 380 -3417 406
rect -3359 380 -3109 406
rect -3051 380 -2801 406
rect -2743 380 -2493 406
rect -2435 380 -2185 406
rect -2127 380 -1877 406
rect -1819 380 -1569 406
rect -1511 380 -1261 406
rect -1203 380 -953 406
rect -895 380 -645 406
rect -587 380 -337 406
rect -279 380 -29 406
rect 29 380 279 406
rect 337 380 587 406
rect 645 380 895 406
rect 953 380 1203 406
rect 1261 380 1511 406
rect 1569 380 1819 406
rect 1877 380 2127 406
rect 2185 380 2435 406
rect 2493 380 2743 406
rect 2801 380 3051 406
rect 3109 380 3359 406
rect 3417 380 3667 406
rect 3725 380 3975 406
rect 4033 380 4283 406
rect 4341 380 4591 406
rect 4649 380 4899 406
rect -4899 -355 -4649 -308
rect -4899 -372 -4829 -355
rect -4845 -389 -4829 -372
rect -4719 -372 -4649 -355
rect -4591 -355 -4341 -308
rect -4591 -372 -4521 -355
rect -4719 -389 -4703 -372
rect -4845 -405 -4703 -389
rect -4537 -389 -4521 -372
rect -4411 -372 -4341 -355
rect -4283 -355 -4033 -308
rect -4283 -372 -4213 -355
rect -4411 -389 -4395 -372
rect -4537 -405 -4395 -389
rect -4229 -389 -4213 -372
rect -4103 -372 -4033 -355
rect -3975 -355 -3725 -308
rect -3975 -372 -3905 -355
rect -4103 -389 -4087 -372
rect -4229 -405 -4087 -389
rect -3921 -389 -3905 -372
rect -3795 -372 -3725 -355
rect -3667 -355 -3417 -308
rect -3667 -372 -3597 -355
rect -3795 -389 -3779 -372
rect -3921 -405 -3779 -389
rect -3613 -389 -3597 -372
rect -3487 -372 -3417 -355
rect -3359 -355 -3109 -308
rect -3359 -372 -3289 -355
rect -3487 -389 -3471 -372
rect -3613 -405 -3471 -389
rect -3305 -389 -3289 -372
rect -3179 -372 -3109 -355
rect -3051 -355 -2801 -308
rect -3051 -372 -2981 -355
rect -3179 -389 -3163 -372
rect -3305 -405 -3163 -389
rect -2997 -389 -2981 -372
rect -2871 -372 -2801 -355
rect -2743 -355 -2493 -308
rect -2743 -372 -2673 -355
rect -2871 -389 -2855 -372
rect -2997 -405 -2855 -389
rect -2689 -389 -2673 -372
rect -2563 -372 -2493 -355
rect -2435 -355 -2185 -308
rect -2435 -372 -2365 -355
rect -2563 -389 -2547 -372
rect -2689 -405 -2547 -389
rect -2381 -389 -2365 -372
rect -2255 -372 -2185 -355
rect -2127 -355 -1877 -308
rect -2127 -372 -2057 -355
rect -2255 -389 -2239 -372
rect -2381 -405 -2239 -389
rect -2073 -389 -2057 -372
rect -1947 -372 -1877 -355
rect -1819 -355 -1569 -308
rect -1819 -372 -1749 -355
rect -1947 -389 -1931 -372
rect -2073 -405 -1931 -389
rect -1765 -389 -1749 -372
rect -1639 -372 -1569 -355
rect -1511 -355 -1261 -308
rect -1511 -372 -1441 -355
rect -1639 -389 -1623 -372
rect -1765 -405 -1623 -389
rect -1457 -389 -1441 -372
rect -1331 -372 -1261 -355
rect -1203 -355 -953 -308
rect -1203 -372 -1133 -355
rect -1331 -389 -1315 -372
rect -1457 -405 -1315 -389
rect -1149 -389 -1133 -372
rect -1023 -372 -953 -355
rect -895 -355 -645 -308
rect -895 -372 -825 -355
rect -1023 -389 -1007 -372
rect -1149 -405 -1007 -389
rect -841 -389 -825 -372
rect -715 -372 -645 -355
rect -587 -355 -337 -308
rect -587 -372 -517 -355
rect -715 -389 -699 -372
rect -841 -405 -699 -389
rect -533 -389 -517 -372
rect -407 -372 -337 -355
rect -279 -355 -29 -308
rect -279 -372 -209 -355
rect -407 -389 -391 -372
rect -533 -405 -391 -389
rect -225 -389 -209 -372
rect -99 -372 -29 -355
rect 29 -355 279 -308
rect 29 -372 99 -355
rect -99 -389 -83 -372
rect -225 -405 -83 -389
rect 83 -389 99 -372
rect 209 -372 279 -355
rect 337 -355 587 -308
rect 337 -372 407 -355
rect 209 -389 225 -372
rect 83 -405 225 -389
rect 391 -389 407 -372
rect 517 -372 587 -355
rect 645 -355 895 -308
rect 645 -372 715 -355
rect 517 -389 533 -372
rect 391 -405 533 -389
rect 699 -389 715 -372
rect 825 -372 895 -355
rect 953 -355 1203 -308
rect 953 -372 1023 -355
rect 825 -389 841 -372
rect 699 -405 841 -389
rect 1007 -389 1023 -372
rect 1133 -372 1203 -355
rect 1261 -355 1511 -308
rect 1261 -372 1331 -355
rect 1133 -389 1149 -372
rect 1007 -405 1149 -389
rect 1315 -389 1331 -372
rect 1441 -372 1511 -355
rect 1569 -355 1819 -308
rect 1569 -372 1639 -355
rect 1441 -389 1457 -372
rect 1315 -405 1457 -389
rect 1623 -389 1639 -372
rect 1749 -372 1819 -355
rect 1877 -355 2127 -308
rect 1877 -372 1947 -355
rect 1749 -389 1765 -372
rect 1623 -405 1765 -389
rect 1931 -389 1947 -372
rect 2057 -372 2127 -355
rect 2185 -355 2435 -308
rect 2185 -372 2255 -355
rect 2057 -389 2073 -372
rect 1931 -405 2073 -389
rect 2239 -389 2255 -372
rect 2365 -372 2435 -355
rect 2493 -355 2743 -308
rect 2493 -372 2563 -355
rect 2365 -389 2381 -372
rect 2239 -405 2381 -389
rect 2547 -389 2563 -372
rect 2673 -372 2743 -355
rect 2801 -355 3051 -308
rect 2801 -372 2871 -355
rect 2673 -389 2689 -372
rect 2547 -405 2689 -389
rect 2855 -389 2871 -372
rect 2981 -372 3051 -355
rect 3109 -355 3359 -308
rect 3109 -372 3179 -355
rect 2981 -389 2997 -372
rect 2855 -405 2997 -389
rect 3163 -389 3179 -372
rect 3289 -372 3359 -355
rect 3417 -355 3667 -308
rect 3417 -372 3487 -355
rect 3289 -389 3305 -372
rect 3163 -405 3305 -389
rect 3471 -389 3487 -372
rect 3597 -372 3667 -355
rect 3725 -355 3975 -308
rect 3725 -372 3795 -355
rect 3597 -389 3613 -372
rect 3471 -405 3613 -389
rect 3779 -389 3795 -372
rect 3905 -372 3975 -355
rect 4033 -355 4283 -308
rect 4033 -372 4103 -355
rect 3905 -389 3921 -372
rect 3779 -405 3921 -389
rect 4087 -389 4103 -372
rect 4213 -372 4283 -355
rect 4341 -355 4591 -308
rect 4341 -372 4411 -355
rect 4213 -389 4229 -372
rect 4087 -405 4229 -389
rect 4395 -389 4411 -372
rect 4521 -372 4591 -355
rect 4649 -355 4899 -308
rect 4649 -372 4719 -355
rect 4521 -389 4537 -372
rect 4395 -405 4537 -389
rect 4703 -389 4719 -372
rect 4829 -372 4899 -355
rect 4829 -389 4845 -372
rect 4703 -405 4845 -389
<< polycont >>
rect -4829 -389 -4719 -355
rect -4521 -389 -4411 -355
rect -4213 -389 -4103 -355
rect -3905 -389 -3795 -355
rect -3597 -389 -3487 -355
rect -3289 -389 -3179 -355
rect -2981 -389 -2871 -355
rect -2673 -389 -2563 -355
rect -2365 -389 -2255 -355
rect -2057 -389 -1947 -355
rect -1749 -389 -1639 -355
rect -1441 -389 -1331 -355
rect -1133 -389 -1023 -355
rect -825 -389 -715 -355
rect -517 -389 -407 -355
rect -209 -389 -99 -355
rect 99 -389 209 -355
rect 407 -389 517 -355
rect 715 -389 825 -355
rect 1023 -389 1133 -355
rect 1331 -389 1441 -355
rect 1639 -389 1749 -355
rect 1947 -389 2057 -355
rect 2255 -389 2365 -355
rect 2563 -389 2673 -355
rect 2871 -389 2981 -355
rect 3179 -389 3289 -355
rect 3487 -389 3597 -355
rect 3795 -389 3905 -355
rect 4103 -389 4213 -355
rect 4411 -389 4521 -355
rect 4719 -389 4829 -355
<< locali >>
rect -4945 368 -4911 384
rect -4945 -312 -4911 -296
rect -4637 368 -4603 384
rect -4637 -312 -4603 -296
rect -4329 368 -4295 384
rect -4329 -312 -4295 -296
rect -4021 368 -3987 384
rect -4021 -312 -3987 -296
rect -3713 368 -3679 384
rect -3713 -312 -3679 -296
rect -3405 368 -3371 384
rect -3405 -312 -3371 -296
rect -3097 368 -3063 384
rect -3097 -312 -3063 -296
rect -2789 368 -2755 384
rect -2789 -312 -2755 -296
rect -2481 368 -2447 384
rect -2481 -312 -2447 -296
rect -2173 368 -2139 384
rect -2173 -312 -2139 -296
rect -1865 368 -1831 384
rect -1865 -312 -1831 -296
rect -1557 368 -1523 384
rect -1557 -312 -1523 -296
rect -1249 368 -1215 384
rect -1249 -312 -1215 -296
rect -941 368 -907 384
rect -941 -312 -907 -296
rect -633 368 -599 384
rect -633 -312 -599 -296
rect -325 368 -291 384
rect -325 -312 -291 -296
rect -17 368 17 384
rect -17 -312 17 -296
rect 291 368 325 384
rect 291 -312 325 -296
rect 599 368 633 384
rect 599 -312 633 -296
rect 907 368 941 384
rect 907 -312 941 -296
rect 1215 368 1249 384
rect 1215 -312 1249 -296
rect 1523 368 1557 384
rect 1523 -312 1557 -296
rect 1831 368 1865 384
rect 1831 -312 1865 -296
rect 2139 368 2173 384
rect 2139 -312 2173 -296
rect 2447 368 2481 384
rect 2447 -312 2481 -296
rect 2755 368 2789 384
rect 2755 -312 2789 -296
rect 3063 368 3097 384
rect 3063 -312 3097 -296
rect 3371 368 3405 384
rect 3371 -312 3405 -296
rect 3679 368 3713 384
rect 3679 -312 3713 -296
rect 3987 368 4021 384
rect 3987 -312 4021 -296
rect 4295 368 4329 384
rect 4295 -312 4329 -296
rect 4603 368 4637 384
rect 4603 -312 4637 -296
rect 4911 368 4945 384
rect 4911 -312 4945 -296
rect -4845 -389 -4829 -355
rect -4719 -389 -4703 -355
rect -4537 -389 -4521 -355
rect -4411 -389 -4395 -355
rect -4229 -389 -4213 -355
rect -4103 -389 -4087 -355
rect -3921 -389 -3905 -355
rect -3795 -389 -3779 -355
rect -3613 -389 -3597 -355
rect -3487 -389 -3471 -355
rect -3305 -389 -3289 -355
rect -3179 -389 -3163 -355
rect -2997 -389 -2981 -355
rect -2871 -389 -2855 -355
rect -2689 -389 -2673 -355
rect -2563 -389 -2547 -355
rect -2381 -389 -2365 -355
rect -2255 -389 -2239 -355
rect -2073 -389 -2057 -355
rect -1947 -389 -1931 -355
rect -1765 -389 -1749 -355
rect -1639 -389 -1623 -355
rect -1457 -389 -1441 -355
rect -1331 -389 -1315 -355
rect -1149 -389 -1133 -355
rect -1023 -389 -1007 -355
rect -841 -389 -825 -355
rect -715 -389 -699 -355
rect -533 -389 -517 -355
rect -407 -389 -391 -355
rect -225 -389 -209 -355
rect -99 -389 -83 -355
rect 83 -389 99 -355
rect 209 -389 225 -355
rect 391 -389 407 -355
rect 517 -389 533 -355
rect 699 -389 715 -355
rect 825 -389 841 -355
rect 1007 -389 1023 -355
rect 1133 -389 1149 -355
rect 1315 -389 1331 -355
rect 1441 -389 1457 -355
rect 1623 -389 1639 -355
rect 1749 -389 1765 -355
rect 1931 -389 1947 -355
rect 2057 -389 2073 -355
rect 2239 -389 2255 -355
rect 2365 -389 2381 -355
rect 2547 -389 2563 -355
rect 2673 -389 2689 -355
rect 2855 -389 2871 -355
rect 2981 -389 2997 -355
rect 3163 -389 3179 -355
rect 3289 -389 3305 -355
rect 3471 -389 3487 -355
rect 3597 -389 3613 -355
rect 3779 -389 3795 -355
rect 3905 -389 3921 -355
rect 4087 -389 4103 -355
rect 4213 -389 4229 -355
rect 4395 -389 4411 -355
rect 4521 -389 4537 -355
rect 4703 -389 4719 -355
rect 4829 -389 4845 -355
<< viali >>
rect -4945 -296 -4911 368
rect -4637 -296 -4603 368
rect -4329 -296 -4295 368
rect -4021 -296 -3987 368
rect -3713 -296 -3679 368
rect -3405 -296 -3371 368
rect -3097 -296 -3063 368
rect -2789 -296 -2755 368
rect -2481 -296 -2447 368
rect -2173 -296 -2139 368
rect -1865 -296 -1831 368
rect -1557 -296 -1523 368
rect -1249 -296 -1215 368
rect -941 -296 -907 368
rect -633 -296 -599 368
rect -325 -296 -291 368
rect -17 -296 17 368
rect 291 -296 325 368
rect 599 -296 633 368
rect 907 -296 941 368
rect 1215 -296 1249 368
rect 1523 -296 1557 368
rect 1831 -296 1865 368
rect 2139 -296 2173 368
rect 2447 -296 2481 368
rect 2755 -296 2789 368
rect 3063 -296 3097 368
rect 3371 -296 3405 368
rect 3679 -296 3713 368
rect 3987 -296 4021 368
rect 4295 -296 4329 368
rect 4603 -296 4637 368
rect 4911 -296 4945 368
rect -4829 -389 -4719 -355
rect -4521 -389 -4411 -355
rect -4213 -389 -4103 -355
rect -3905 -389 -3795 -355
rect -3597 -389 -3487 -355
rect -3289 -389 -3179 -355
rect -2981 -389 -2871 -355
rect -2673 -389 -2563 -355
rect -2365 -389 -2255 -355
rect -2057 -389 -1947 -355
rect -1749 -389 -1639 -355
rect -1441 -389 -1331 -355
rect -1133 -389 -1023 -355
rect -825 -389 -715 -355
rect -517 -389 -407 -355
rect -209 -389 -99 -355
rect 99 -389 209 -355
rect 407 -389 517 -355
rect 715 -389 825 -355
rect 1023 -389 1133 -355
rect 1331 -389 1441 -355
rect 1639 -389 1749 -355
rect 1947 -389 2057 -355
rect 2255 -389 2365 -355
rect 2563 -389 2673 -355
rect 2871 -389 2981 -355
rect 3179 -389 3289 -355
rect 3487 -389 3597 -355
rect 3795 -389 3905 -355
rect 4103 -389 4213 -355
rect 4411 -389 4521 -355
rect 4719 -389 4829 -355
<< metal1 >>
rect -4951 368 -4905 380
rect -4951 -296 -4945 368
rect -4911 -296 -4905 368
rect -4951 -308 -4905 -296
rect -4643 368 -4597 380
rect -4643 -296 -4637 368
rect -4603 -296 -4597 368
rect -4643 -308 -4597 -296
rect -4335 368 -4289 380
rect -4335 -296 -4329 368
rect -4295 -296 -4289 368
rect -4335 -308 -4289 -296
rect -4027 368 -3981 380
rect -4027 -296 -4021 368
rect -3987 -296 -3981 368
rect -4027 -308 -3981 -296
rect -3719 368 -3673 380
rect -3719 -296 -3713 368
rect -3679 -296 -3673 368
rect -3719 -308 -3673 -296
rect -3411 368 -3365 380
rect -3411 -296 -3405 368
rect -3371 -296 -3365 368
rect -3411 -308 -3365 -296
rect -3103 368 -3057 380
rect -3103 -296 -3097 368
rect -3063 -296 -3057 368
rect -3103 -308 -3057 -296
rect -2795 368 -2749 380
rect -2795 -296 -2789 368
rect -2755 -296 -2749 368
rect -2795 -308 -2749 -296
rect -2487 368 -2441 380
rect -2487 -296 -2481 368
rect -2447 -296 -2441 368
rect -2487 -308 -2441 -296
rect -2179 368 -2133 380
rect -2179 -296 -2173 368
rect -2139 -296 -2133 368
rect -2179 -308 -2133 -296
rect -1871 368 -1825 380
rect -1871 -296 -1865 368
rect -1831 -296 -1825 368
rect -1871 -308 -1825 -296
rect -1563 368 -1517 380
rect -1563 -296 -1557 368
rect -1523 -296 -1517 368
rect -1563 -308 -1517 -296
rect -1255 368 -1209 380
rect -1255 -296 -1249 368
rect -1215 -296 -1209 368
rect -1255 -308 -1209 -296
rect -947 368 -901 380
rect -947 -296 -941 368
rect -907 -296 -901 368
rect -947 -308 -901 -296
rect -639 368 -593 380
rect -639 -296 -633 368
rect -599 -296 -593 368
rect -639 -308 -593 -296
rect -331 368 -285 380
rect -331 -296 -325 368
rect -291 -296 -285 368
rect -331 -308 -285 -296
rect -23 368 23 380
rect -23 -296 -17 368
rect 17 -296 23 368
rect -23 -308 23 -296
rect 285 368 331 380
rect 285 -296 291 368
rect 325 -296 331 368
rect 285 -308 331 -296
rect 593 368 639 380
rect 593 -296 599 368
rect 633 -296 639 368
rect 593 -308 639 -296
rect 901 368 947 380
rect 901 -296 907 368
rect 941 -296 947 368
rect 901 -308 947 -296
rect 1209 368 1255 380
rect 1209 -296 1215 368
rect 1249 -296 1255 368
rect 1209 -308 1255 -296
rect 1517 368 1563 380
rect 1517 -296 1523 368
rect 1557 -296 1563 368
rect 1517 -308 1563 -296
rect 1825 368 1871 380
rect 1825 -296 1831 368
rect 1865 -296 1871 368
rect 1825 -308 1871 -296
rect 2133 368 2179 380
rect 2133 -296 2139 368
rect 2173 -296 2179 368
rect 2133 -308 2179 -296
rect 2441 368 2487 380
rect 2441 -296 2447 368
rect 2481 -296 2487 368
rect 2441 -308 2487 -296
rect 2749 368 2795 380
rect 2749 -296 2755 368
rect 2789 -296 2795 368
rect 2749 -308 2795 -296
rect 3057 368 3103 380
rect 3057 -296 3063 368
rect 3097 -296 3103 368
rect 3057 -308 3103 -296
rect 3365 368 3411 380
rect 3365 -296 3371 368
rect 3405 -296 3411 368
rect 3365 -308 3411 -296
rect 3673 368 3719 380
rect 3673 -296 3679 368
rect 3713 -296 3719 368
rect 3673 -308 3719 -296
rect 3981 368 4027 380
rect 3981 -296 3987 368
rect 4021 -296 4027 368
rect 3981 -308 4027 -296
rect 4289 368 4335 380
rect 4289 -296 4295 368
rect 4329 -296 4335 368
rect 4289 -308 4335 -296
rect 4597 368 4643 380
rect 4597 -296 4603 368
rect 4637 -296 4643 368
rect 4597 -308 4643 -296
rect 4905 368 4951 380
rect 4905 -296 4911 368
rect 4945 -296 4951 368
rect 4905 -308 4951 -296
rect -4841 -355 -4707 -349
rect -4841 -389 -4829 -355
rect -4719 -389 -4707 -355
rect -4841 -395 -4707 -389
rect -4533 -355 -4399 -349
rect -4533 -389 -4521 -355
rect -4411 -389 -4399 -355
rect -4533 -395 -4399 -389
rect -4225 -355 -4091 -349
rect -4225 -389 -4213 -355
rect -4103 -389 -4091 -355
rect -4225 -395 -4091 -389
rect -3917 -355 -3783 -349
rect -3917 -389 -3905 -355
rect -3795 -389 -3783 -355
rect -3917 -395 -3783 -389
rect -3609 -355 -3475 -349
rect -3609 -389 -3597 -355
rect -3487 -389 -3475 -355
rect -3609 -395 -3475 -389
rect -3301 -355 -3167 -349
rect -3301 -389 -3289 -355
rect -3179 -389 -3167 -355
rect -3301 -395 -3167 -389
rect -2993 -355 -2859 -349
rect -2993 -389 -2981 -355
rect -2871 -389 -2859 -355
rect -2993 -395 -2859 -389
rect -2685 -355 -2551 -349
rect -2685 -389 -2673 -355
rect -2563 -389 -2551 -355
rect -2685 -395 -2551 -389
rect -2377 -355 -2243 -349
rect -2377 -389 -2365 -355
rect -2255 -389 -2243 -355
rect -2377 -395 -2243 -389
rect -2069 -355 -1935 -349
rect -2069 -389 -2057 -355
rect -1947 -389 -1935 -355
rect -2069 -395 -1935 -389
rect -1761 -355 -1627 -349
rect -1761 -389 -1749 -355
rect -1639 -389 -1627 -355
rect -1761 -395 -1627 -389
rect -1453 -355 -1319 -349
rect -1453 -389 -1441 -355
rect -1331 -389 -1319 -355
rect -1453 -395 -1319 -389
rect -1145 -355 -1011 -349
rect -1145 -389 -1133 -355
rect -1023 -389 -1011 -355
rect -1145 -395 -1011 -389
rect -837 -355 -703 -349
rect -837 -389 -825 -355
rect -715 -389 -703 -355
rect -837 -395 -703 -389
rect -529 -355 -395 -349
rect -529 -389 -517 -355
rect -407 -389 -395 -355
rect -529 -395 -395 -389
rect -221 -355 -87 -349
rect -221 -389 -209 -355
rect -99 -389 -87 -355
rect -221 -395 -87 -389
rect 87 -355 221 -349
rect 87 -389 99 -355
rect 209 -389 221 -355
rect 87 -395 221 -389
rect 395 -355 529 -349
rect 395 -389 407 -355
rect 517 -389 529 -355
rect 395 -395 529 -389
rect 703 -355 837 -349
rect 703 -389 715 -355
rect 825 -389 837 -355
rect 703 -395 837 -389
rect 1011 -355 1145 -349
rect 1011 -389 1023 -355
rect 1133 -389 1145 -355
rect 1011 -395 1145 -389
rect 1319 -355 1453 -349
rect 1319 -389 1331 -355
rect 1441 -389 1453 -355
rect 1319 -395 1453 -389
rect 1627 -355 1761 -349
rect 1627 -389 1639 -355
rect 1749 -389 1761 -355
rect 1627 -395 1761 -389
rect 1935 -355 2069 -349
rect 1935 -389 1947 -355
rect 2057 -389 2069 -355
rect 1935 -395 2069 -389
rect 2243 -355 2377 -349
rect 2243 -389 2255 -355
rect 2365 -389 2377 -355
rect 2243 -395 2377 -389
rect 2551 -355 2685 -349
rect 2551 -389 2563 -355
rect 2673 -389 2685 -355
rect 2551 -395 2685 -389
rect 2859 -355 2993 -349
rect 2859 -389 2871 -355
rect 2981 -389 2993 -355
rect 2859 -395 2993 -389
rect 3167 -355 3301 -349
rect 3167 -389 3179 -355
rect 3289 -389 3301 -355
rect 3167 -395 3301 -389
rect 3475 -355 3609 -349
rect 3475 -389 3487 -355
rect 3597 -389 3609 -355
rect 3475 -395 3609 -389
rect 3783 -355 3917 -349
rect 3783 -389 3795 -355
rect 3905 -389 3917 -355
rect 3783 -395 3917 -389
rect 4091 -355 4225 -349
rect 4091 -389 4103 -355
rect 4213 -389 4225 -355
rect 4091 -395 4225 -389
rect 4399 -355 4533 -349
rect 4399 -389 4411 -355
rect 4521 -389 4533 -355
rect 4399 -395 4533 -389
rect 4707 -355 4841 -349
rect 4707 -389 4719 -355
rect 4829 -389 4841 -355
rect 4707 -395 4841 -389
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.4375 l 1.25 m 1 nf 32 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
