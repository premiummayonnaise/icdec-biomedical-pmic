magic
tech sky130A
magscale 1 2
timestamp 1768990256
<< error_p >>
rect -3459 1038 3459 1042
rect -3459 -970 -3429 1038
rect -3393 972 -3027 976
rect -2965 972 -2599 976
rect -2537 972 -2171 976
rect -2109 972 -1743 976
rect -1681 972 -1315 976
rect -1253 972 -887 976
rect -825 972 -459 976
rect -397 972 -31 976
rect 31 972 397 976
rect 459 972 825 976
rect 887 972 1253 976
rect 1315 972 1681 976
rect 1743 972 2109 976
rect 2171 972 2537 976
rect 2599 972 2965 976
rect 3027 972 3393 976
rect -3393 -904 -3363 972
rect 3363 -904 3393 972
rect 3429 -970 3459 1038
<< nwell >>
rect -3429 -1004 3429 1038
<< mvpmos >>
rect -3335 -904 -3085 976
rect -2907 -904 -2657 976
rect -2479 -904 -2229 976
rect -2051 -904 -1801 976
rect -1623 -904 -1373 976
rect -1195 -904 -945 976
rect -767 -904 -517 976
rect -339 -904 -89 976
rect 89 -904 339 976
rect 517 -904 767 976
rect 945 -904 1195 976
rect 1373 -904 1623 976
rect 1801 -904 2051 976
rect 2229 -904 2479 976
rect 2657 -904 2907 976
rect 3085 -904 3335 976
<< mvpdiff >>
rect -3393 964 -3335 976
rect -3393 -892 -3381 964
rect -3347 -892 -3335 964
rect -3393 -904 -3335 -892
rect -3085 964 -3027 976
rect -3085 -892 -3073 964
rect -3039 -892 -3027 964
rect -3085 -904 -3027 -892
rect -2965 964 -2907 976
rect -2965 -892 -2953 964
rect -2919 -892 -2907 964
rect -2965 -904 -2907 -892
rect -2657 964 -2599 976
rect -2657 -892 -2645 964
rect -2611 -892 -2599 964
rect -2657 -904 -2599 -892
rect -2537 964 -2479 976
rect -2537 -892 -2525 964
rect -2491 -892 -2479 964
rect -2537 -904 -2479 -892
rect -2229 964 -2171 976
rect -2229 -892 -2217 964
rect -2183 -892 -2171 964
rect -2229 -904 -2171 -892
rect -2109 964 -2051 976
rect -2109 -892 -2097 964
rect -2063 -892 -2051 964
rect -2109 -904 -2051 -892
rect -1801 964 -1743 976
rect -1801 -892 -1789 964
rect -1755 -892 -1743 964
rect -1801 -904 -1743 -892
rect -1681 964 -1623 976
rect -1681 -892 -1669 964
rect -1635 -892 -1623 964
rect -1681 -904 -1623 -892
rect -1373 964 -1315 976
rect -1373 -892 -1361 964
rect -1327 -892 -1315 964
rect -1373 -904 -1315 -892
rect -1253 964 -1195 976
rect -1253 -892 -1241 964
rect -1207 -892 -1195 964
rect -1253 -904 -1195 -892
rect -945 964 -887 976
rect -945 -892 -933 964
rect -899 -892 -887 964
rect -945 -904 -887 -892
rect -825 964 -767 976
rect -825 -892 -813 964
rect -779 -892 -767 964
rect -825 -904 -767 -892
rect -517 964 -459 976
rect -517 -892 -505 964
rect -471 -892 -459 964
rect -517 -904 -459 -892
rect -397 964 -339 976
rect -397 -892 -385 964
rect -351 -892 -339 964
rect -397 -904 -339 -892
rect -89 964 -31 976
rect -89 -892 -77 964
rect -43 -892 -31 964
rect -89 -904 -31 -892
rect 31 964 89 976
rect 31 -892 43 964
rect 77 -892 89 964
rect 31 -904 89 -892
rect 339 964 397 976
rect 339 -892 351 964
rect 385 -892 397 964
rect 339 -904 397 -892
rect 459 964 517 976
rect 459 -892 471 964
rect 505 -892 517 964
rect 459 -904 517 -892
rect 767 964 825 976
rect 767 -892 779 964
rect 813 -892 825 964
rect 767 -904 825 -892
rect 887 964 945 976
rect 887 -892 899 964
rect 933 -892 945 964
rect 887 -904 945 -892
rect 1195 964 1253 976
rect 1195 -892 1207 964
rect 1241 -892 1253 964
rect 1195 -904 1253 -892
rect 1315 964 1373 976
rect 1315 -892 1327 964
rect 1361 -892 1373 964
rect 1315 -904 1373 -892
rect 1623 964 1681 976
rect 1623 -892 1635 964
rect 1669 -892 1681 964
rect 1623 -904 1681 -892
rect 1743 964 1801 976
rect 1743 -892 1755 964
rect 1789 -892 1801 964
rect 1743 -904 1801 -892
rect 2051 964 2109 976
rect 2051 -892 2063 964
rect 2097 -892 2109 964
rect 2051 -904 2109 -892
rect 2171 964 2229 976
rect 2171 -892 2183 964
rect 2217 -892 2229 964
rect 2171 -904 2229 -892
rect 2479 964 2537 976
rect 2479 -892 2491 964
rect 2525 -892 2537 964
rect 2479 -904 2537 -892
rect 2599 964 2657 976
rect 2599 -892 2611 964
rect 2645 -892 2657 964
rect 2599 -904 2657 -892
rect 2907 964 2965 976
rect 2907 -892 2919 964
rect 2953 -892 2965 964
rect 2907 -904 2965 -892
rect 3027 964 3085 976
rect 3027 -892 3039 964
rect 3073 -892 3085 964
rect 3027 -904 3085 -892
rect 3335 964 3393 976
rect 3335 -892 3347 964
rect 3381 -892 3393 964
rect 3335 -904 3393 -892
<< mvpdiffc >>
rect -3381 -892 -3347 964
rect -3073 -892 -3039 964
rect -2953 -892 -2919 964
rect -2645 -892 -2611 964
rect -2525 -892 -2491 964
rect -2217 -892 -2183 964
rect -2097 -892 -2063 964
rect -1789 -892 -1755 964
rect -1669 -892 -1635 964
rect -1361 -892 -1327 964
rect -1241 -892 -1207 964
rect -933 -892 -899 964
rect -813 -892 -779 964
rect -505 -892 -471 964
rect -385 -892 -351 964
rect -77 -892 -43 964
rect 43 -892 77 964
rect 351 -892 385 964
rect 471 -892 505 964
rect 779 -892 813 964
rect 899 -892 933 964
rect 1207 -892 1241 964
rect 1327 -892 1361 964
rect 1635 -892 1669 964
rect 1755 -892 1789 964
rect 2063 -892 2097 964
rect 2183 -892 2217 964
rect 2491 -892 2525 964
rect 2611 -892 2645 964
rect 2919 -892 2953 964
rect 3039 -892 3073 964
rect 3347 -892 3381 964
<< poly >>
rect -3335 976 -3085 1002
rect -2907 976 -2657 1002
rect -2479 976 -2229 1002
rect -2051 976 -1801 1002
rect -1623 976 -1373 1002
rect -1195 976 -945 1002
rect -767 976 -517 1002
rect -339 976 -89 1002
rect 89 976 339 1002
rect 517 976 767 1002
rect 945 976 1195 1002
rect 1373 976 1623 1002
rect 1801 976 2051 1002
rect 2229 976 2479 1002
rect 2657 976 2907 1002
rect 3085 976 3335 1002
rect -3335 -951 -3085 -904
rect -3335 -985 -3319 -951
rect -3101 -985 -3085 -951
rect -3335 -1001 -3085 -985
rect -2907 -951 -2657 -904
rect -2907 -985 -2891 -951
rect -2673 -985 -2657 -951
rect -2907 -1001 -2657 -985
rect -2479 -951 -2229 -904
rect -2479 -985 -2463 -951
rect -2245 -985 -2229 -951
rect -2479 -1001 -2229 -985
rect -2051 -951 -1801 -904
rect -2051 -985 -2035 -951
rect -1817 -985 -1801 -951
rect -2051 -1001 -1801 -985
rect -1623 -951 -1373 -904
rect -1623 -985 -1607 -951
rect -1389 -985 -1373 -951
rect -1623 -1001 -1373 -985
rect -1195 -951 -945 -904
rect -1195 -985 -1179 -951
rect -961 -985 -945 -951
rect -1195 -1001 -945 -985
rect -767 -951 -517 -904
rect -767 -985 -751 -951
rect -533 -985 -517 -951
rect -767 -1001 -517 -985
rect -339 -951 -89 -904
rect -339 -985 -323 -951
rect -105 -985 -89 -951
rect -339 -1001 -89 -985
rect 89 -951 339 -904
rect 89 -985 105 -951
rect 323 -985 339 -951
rect 89 -1001 339 -985
rect 517 -951 767 -904
rect 517 -985 533 -951
rect 751 -985 767 -951
rect 517 -1001 767 -985
rect 945 -951 1195 -904
rect 945 -985 961 -951
rect 1179 -985 1195 -951
rect 945 -1001 1195 -985
rect 1373 -951 1623 -904
rect 1373 -985 1389 -951
rect 1607 -985 1623 -951
rect 1373 -1001 1623 -985
rect 1801 -951 2051 -904
rect 1801 -985 1817 -951
rect 2035 -985 2051 -951
rect 1801 -1001 2051 -985
rect 2229 -951 2479 -904
rect 2229 -985 2245 -951
rect 2463 -985 2479 -951
rect 2229 -1001 2479 -985
rect 2657 -951 2907 -904
rect 2657 -985 2673 -951
rect 2891 -985 2907 -951
rect 2657 -1001 2907 -985
rect 3085 -951 3335 -904
rect 3085 -985 3101 -951
rect 3319 -985 3335 -951
rect 3085 -1001 3335 -985
<< polycont >>
rect -3319 -985 -3101 -951
rect -2891 -985 -2673 -951
rect -2463 -985 -2245 -951
rect -2035 -985 -1817 -951
rect -1607 -985 -1389 -951
rect -1179 -985 -961 -951
rect -751 -985 -533 -951
rect -323 -985 -105 -951
rect 105 -985 323 -951
rect 533 -985 751 -951
rect 961 -985 1179 -951
rect 1389 -985 1607 -951
rect 1817 -985 2035 -951
rect 2245 -985 2463 -951
rect 2673 -985 2891 -951
rect 3101 -985 3319 -951
<< locali >>
rect -3381 964 -3347 980
rect -3381 -908 -3347 -892
rect -3073 964 -3039 980
rect -3073 -908 -3039 -892
rect -2953 964 -2919 980
rect -2953 -908 -2919 -892
rect -2645 964 -2611 980
rect -2645 -908 -2611 -892
rect -2525 964 -2491 980
rect -2525 -908 -2491 -892
rect -2217 964 -2183 980
rect -2217 -908 -2183 -892
rect -2097 964 -2063 980
rect -2097 -908 -2063 -892
rect -1789 964 -1755 980
rect -1789 -908 -1755 -892
rect -1669 964 -1635 980
rect -1669 -908 -1635 -892
rect -1361 964 -1327 980
rect -1361 -908 -1327 -892
rect -1241 964 -1207 980
rect -1241 -908 -1207 -892
rect -933 964 -899 980
rect -933 -908 -899 -892
rect -813 964 -779 980
rect -813 -908 -779 -892
rect -505 964 -471 980
rect -505 -908 -471 -892
rect -385 964 -351 980
rect -385 -908 -351 -892
rect -77 964 -43 980
rect -77 -908 -43 -892
rect 43 964 77 980
rect 43 -908 77 -892
rect 351 964 385 980
rect 351 -908 385 -892
rect 471 964 505 980
rect 471 -908 505 -892
rect 779 964 813 980
rect 779 -908 813 -892
rect 899 964 933 980
rect 899 -908 933 -892
rect 1207 964 1241 980
rect 1207 -908 1241 -892
rect 1327 964 1361 980
rect 1327 -908 1361 -892
rect 1635 964 1669 980
rect 1635 -908 1669 -892
rect 1755 964 1789 980
rect 1755 -908 1789 -892
rect 2063 964 2097 980
rect 2063 -908 2097 -892
rect 2183 964 2217 980
rect 2183 -908 2217 -892
rect 2491 964 2525 980
rect 2491 -908 2525 -892
rect 2611 964 2645 980
rect 2611 -908 2645 -892
rect 2919 964 2953 980
rect 2919 -908 2953 -892
rect 3039 964 3073 980
rect 3039 -908 3073 -892
rect 3347 964 3381 980
rect 3347 -908 3381 -892
rect -3335 -985 -3319 -951
rect -3101 -985 -3085 -951
rect -2907 -985 -2891 -951
rect -2673 -985 -2657 -951
rect -2479 -985 -2463 -951
rect -2245 -985 -2229 -951
rect -2051 -985 -2035 -951
rect -1817 -985 -1801 -951
rect -1623 -985 -1607 -951
rect -1389 -985 -1373 -951
rect -1195 -985 -1179 -951
rect -961 -985 -945 -951
rect -767 -985 -751 -951
rect -533 -985 -517 -951
rect -339 -985 -323 -951
rect -105 -985 -89 -951
rect 89 -985 105 -951
rect 323 -985 339 -951
rect 517 -985 533 -951
rect 751 -985 767 -951
rect 945 -985 961 -951
rect 1179 -985 1195 -951
rect 1373 -985 1389 -951
rect 1607 -985 1623 -951
rect 1801 -985 1817 -951
rect 2035 -985 2051 -951
rect 2229 -985 2245 -951
rect 2463 -985 2479 -951
rect 2657 -985 2673 -951
rect 2891 -985 2907 -951
rect 3085 -985 3101 -951
rect 3319 -985 3335 -951
<< viali >>
rect -3381 -892 -3347 964
rect -3073 -892 -3039 964
rect -2953 -892 -2919 964
rect -2645 -892 -2611 964
rect -2525 -892 -2491 964
rect -2217 -892 -2183 964
rect -2097 -892 -2063 964
rect -1789 -892 -1755 964
rect -1669 -892 -1635 964
rect -1361 -892 -1327 964
rect -1241 -892 -1207 964
rect -933 -892 -899 964
rect -813 -892 -779 964
rect -505 -892 -471 964
rect -385 -892 -351 964
rect -77 -892 -43 964
rect 43 -892 77 964
rect 351 -892 385 964
rect 471 -892 505 964
rect 779 -892 813 964
rect 899 -892 933 964
rect 1207 -892 1241 964
rect 1327 -892 1361 964
rect 1635 -892 1669 964
rect 1755 -892 1789 964
rect 2063 -892 2097 964
rect 2183 -892 2217 964
rect 2491 -892 2525 964
rect 2611 -892 2645 964
rect 2919 -892 2953 964
rect 3039 -892 3073 964
rect 3347 -892 3381 964
rect -3319 -985 -3101 -951
rect -2891 -985 -2673 -951
rect -2463 -985 -2245 -951
rect -2035 -985 -1817 -951
rect -1607 -985 -1389 -951
rect -1179 -985 -961 -951
rect -751 -985 -533 -951
rect -323 -985 -105 -951
rect 105 -985 323 -951
rect 533 -985 751 -951
rect 961 -985 1179 -951
rect 1389 -985 1607 -951
rect 1817 -985 2035 -951
rect 2245 -985 2463 -951
rect 2673 -985 2891 -951
rect 3101 -985 3319 -951
<< metal1 >>
rect -3387 964 -3341 976
rect -3387 -892 -3381 964
rect -3347 -892 -3341 964
rect -3387 -904 -3341 -892
rect -3079 964 -3033 976
rect -3079 -892 -3073 964
rect -3039 -892 -3033 964
rect -3079 -904 -3033 -892
rect -2959 964 -2913 976
rect -2959 -892 -2953 964
rect -2919 -892 -2913 964
rect -2959 -904 -2913 -892
rect -2651 964 -2605 976
rect -2651 -892 -2645 964
rect -2611 -892 -2605 964
rect -2651 -904 -2605 -892
rect -2531 964 -2485 976
rect -2531 -892 -2525 964
rect -2491 -892 -2485 964
rect -2531 -904 -2485 -892
rect -2223 964 -2177 976
rect -2223 -892 -2217 964
rect -2183 -892 -2177 964
rect -2223 -904 -2177 -892
rect -2103 964 -2057 976
rect -2103 -892 -2097 964
rect -2063 -892 -2057 964
rect -2103 -904 -2057 -892
rect -1795 964 -1749 976
rect -1795 -892 -1789 964
rect -1755 -892 -1749 964
rect -1795 -904 -1749 -892
rect -1675 964 -1629 976
rect -1675 -892 -1669 964
rect -1635 -892 -1629 964
rect -1675 -904 -1629 -892
rect -1367 964 -1321 976
rect -1367 -892 -1361 964
rect -1327 -892 -1321 964
rect -1367 -904 -1321 -892
rect -1247 964 -1201 976
rect -1247 -892 -1241 964
rect -1207 -892 -1201 964
rect -1247 -904 -1201 -892
rect -939 964 -893 976
rect -939 -892 -933 964
rect -899 -892 -893 964
rect -939 -904 -893 -892
rect -819 964 -773 976
rect -819 -892 -813 964
rect -779 -892 -773 964
rect -819 -904 -773 -892
rect -511 964 -465 976
rect -511 -892 -505 964
rect -471 -892 -465 964
rect -511 -904 -465 -892
rect -391 964 -345 976
rect -391 -892 -385 964
rect -351 -892 -345 964
rect -391 -904 -345 -892
rect -83 964 -37 976
rect -83 -892 -77 964
rect -43 -892 -37 964
rect -83 -904 -37 -892
rect 37 964 83 976
rect 37 -892 43 964
rect 77 -892 83 964
rect 37 -904 83 -892
rect 345 964 391 976
rect 345 -892 351 964
rect 385 -892 391 964
rect 345 -904 391 -892
rect 465 964 511 976
rect 465 -892 471 964
rect 505 -892 511 964
rect 465 -904 511 -892
rect 773 964 819 976
rect 773 -892 779 964
rect 813 -892 819 964
rect 773 -904 819 -892
rect 893 964 939 976
rect 893 -892 899 964
rect 933 -892 939 964
rect 893 -904 939 -892
rect 1201 964 1247 976
rect 1201 -892 1207 964
rect 1241 -892 1247 964
rect 1201 -904 1247 -892
rect 1321 964 1367 976
rect 1321 -892 1327 964
rect 1361 -892 1367 964
rect 1321 -904 1367 -892
rect 1629 964 1675 976
rect 1629 -892 1635 964
rect 1669 -892 1675 964
rect 1629 -904 1675 -892
rect 1749 964 1795 976
rect 1749 -892 1755 964
rect 1789 -892 1795 964
rect 1749 -904 1795 -892
rect 2057 964 2103 976
rect 2057 -892 2063 964
rect 2097 -892 2103 964
rect 2057 -904 2103 -892
rect 2177 964 2223 976
rect 2177 -892 2183 964
rect 2217 -892 2223 964
rect 2177 -904 2223 -892
rect 2485 964 2531 976
rect 2485 -892 2491 964
rect 2525 -892 2531 964
rect 2485 -904 2531 -892
rect 2605 964 2651 976
rect 2605 -892 2611 964
rect 2645 -892 2651 964
rect 2605 -904 2651 -892
rect 2913 964 2959 976
rect 2913 -892 2919 964
rect 2953 -892 2959 964
rect 2913 -904 2959 -892
rect 3033 964 3079 976
rect 3033 -892 3039 964
rect 3073 -892 3079 964
rect 3033 -904 3079 -892
rect 3341 964 3387 976
rect 3341 -892 3347 964
rect 3381 -892 3387 964
rect 3341 -904 3387 -892
rect -3331 -951 -3089 -945
rect -3331 -985 -3319 -951
rect -3101 -985 -3089 -951
rect -3331 -991 -3089 -985
rect -2903 -951 -2661 -945
rect -2903 -985 -2891 -951
rect -2673 -985 -2661 -951
rect -2903 -991 -2661 -985
rect -2475 -951 -2233 -945
rect -2475 -985 -2463 -951
rect -2245 -985 -2233 -951
rect -2475 -991 -2233 -985
rect -2047 -951 -1805 -945
rect -2047 -985 -2035 -951
rect -1817 -985 -1805 -951
rect -2047 -991 -1805 -985
rect -1619 -951 -1377 -945
rect -1619 -985 -1607 -951
rect -1389 -985 -1377 -951
rect -1619 -991 -1377 -985
rect -1191 -951 -949 -945
rect -1191 -985 -1179 -951
rect -961 -985 -949 -951
rect -1191 -991 -949 -985
rect -763 -951 -521 -945
rect -763 -985 -751 -951
rect -533 -985 -521 -951
rect -763 -991 -521 -985
rect -335 -951 -93 -945
rect -335 -985 -323 -951
rect -105 -985 -93 -951
rect -335 -991 -93 -985
rect 93 -951 335 -945
rect 93 -985 105 -951
rect 323 -985 335 -951
rect 93 -991 335 -985
rect 521 -951 763 -945
rect 521 -985 533 -951
rect 751 -985 763 -951
rect 521 -991 763 -985
rect 949 -951 1191 -945
rect 949 -985 961 -951
rect 1179 -985 1191 -951
rect 949 -991 1191 -985
rect 1377 -951 1619 -945
rect 1377 -985 1389 -951
rect 1607 -985 1619 -951
rect 1377 -991 1619 -985
rect 1805 -951 2047 -945
rect 1805 -985 1817 -951
rect 2035 -985 2047 -951
rect 1805 -991 2047 -985
rect 2233 -951 2475 -945
rect 2233 -985 2245 -951
rect 2463 -985 2475 -951
rect 2233 -991 2475 -985
rect 2661 -951 2903 -945
rect 2661 -985 2673 -951
rect 2891 -985 2903 -951
rect 2661 -991 2903 -985
rect 3089 -951 3331 -945
rect 3089 -985 3101 -951
rect 3319 -985 3331 -951
rect 3089 -991 3331 -985
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9.4 l 1.25 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
