magic
tech sky130A
magscale 1 2
timestamp 1769400417
<< metal3 >>
rect -9104 2012 -4732 2040
rect -9104 -2012 -4816 2012
rect -4752 -2012 -4732 2012
rect -9104 -2040 -4732 -2012
rect -4492 2012 -120 2040
rect -4492 -2012 -204 2012
rect -140 -2012 -120 2012
rect -4492 -2040 -120 -2012
rect 120 2012 4492 2040
rect 120 -2012 4408 2012
rect 4472 -2012 4492 2012
rect 120 -2040 4492 -2012
rect 4732 2012 9104 2040
rect 4732 -2012 9020 2012
rect 9084 -2012 9104 2012
rect 4732 -2040 9104 -2012
<< via3 >>
rect -4816 -2012 -4752 2012
rect -204 -2012 -140 2012
rect 4408 -2012 4472 2012
rect 9020 -2012 9084 2012
<< mimcap >>
rect -9064 1960 -5064 2000
rect -9064 -1960 -9024 1960
rect -5104 -1960 -5064 1960
rect -9064 -2000 -5064 -1960
rect -4452 1960 -452 2000
rect -4452 -1960 -4412 1960
rect -492 -1960 -452 1960
rect -4452 -2000 -452 -1960
rect 160 1960 4160 2000
rect 160 -1960 200 1960
rect 4120 -1960 4160 1960
rect 160 -2000 4160 -1960
rect 4772 1960 8772 2000
rect 4772 -1960 4812 1960
rect 8732 -1960 8772 1960
rect 4772 -2000 8772 -1960
<< mimcapcontact >>
rect -9024 -1960 -5104 1960
rect -4412 -1960 -492 1960
rect 200 -1960 4120 1960
rect 4812 -1960 8732 1960
<< metal4 >>
rect -4832 2012 -4736 2028
rect -9025 1960 -5103 1961
rect -9025 -1960 -9024 1960
rect -5104 -1960 -5103 1960
rect -9025 -1961 -5103 -1960
rect -4832 -2012 -4816 2012
rect -4752 -2012 -4736 2012
rect -220 2012 -124 2028
rect -4413 1960 -491 1961
rect -4413 -1960 -4412 1960
rect -492 -1960 -491 1960
rect -4413 -1961 -491 -1960
rect -4832 -2028 -4736 -2012
rect -220 -2012 -204 2012
rect -140 -2012 -124 2012
rect 4392 2012 4488 2028
rect 199 1960 4121 1961
rect 199 -1960 200 1960
rect 4120 -1960 4121 1960
rect 199 -1961 4121 -1960
rect -220 -2028 -124 -2012
rect 4392 -2012 4408 2012
rect 4472 -2012 4488 2012
rect 9004 2012 9100 2028
rect 4811 1960 8733 1961
rect 4811 -1960 4812 1960
rect 8732 -1960 8733 1960
rect 4811 -1961 8733 -1960
rect 4392 -2028 4488 -2012
rect 9004 -2012 9020 2012
rect 9084 -2012 9100 2012
rect 9004 -2028 9100 -2012
<< properties >>
string FIXED_BBOX 4732 -2040 8812 2040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20.0 l 20.0 val 815.2 carea 2.00 cperi 0.19 class capacitor nx 4 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
