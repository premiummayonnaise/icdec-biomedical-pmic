magic
tech sky130A
magscale 1 2
timestamp 1769170054
<< nwell >>
rect -2693 -1415 2693 1415
<< mvpmos >>
rect -2435 118 -2185 1118
rect -2127 118 -1877 1118
rect -1819 118 -1569 1118
rect -1511 118 -1261 1118
rect -1203 118 -953 1118
rect -895 118 -645 1118
rect -587 118 -337 1118
rect -279 118 -29 1118
rect 29 118 279 1118
rect 337 118 587 1118
rect 645 118 895 1118
rect 953 118 1203 1118
rect 1261 118 1511 1118
rect 1569 118 1819 1118
rect 1877 118 2127 1118
rect 2185 118 2435 1118
rect -2435 -1118 -2185 -118
rect -2127 -1118 -1877 -118
rect -1819 -1118 -1569 -118
rect -1511 -1118 -1261 -118
rect -1203 -1118 -953 -118
rect -895 -1118 -645 -118
rect -587 -1118 -337 -118
rect -279 -1118 -29 -118
rect 29 -1118 279 -118
rect 337 -1118 587 -118
rect 645 -1118 895 -118
rect 953 -1118 1203 -118
rect 1261 -1118 1511 -118
rect 1569 -1118 1819 -118
rect 1877 -1118 2127 -118
rect 2185 -1118 2435 -118
<< mvpdiff >>
rect -2493 1106 -2435 1118
rect -2493 130 -2481 1106
rect -2447 130 -2435 1106
rect -2493 118 -2435 130
rect -2185 1106 -2127 1118
rect -2185 130 -2173 1106
rect -2139 130 -2127 1106
rect -2185 118 -2127 130
rect -1877 1106 -1819 1118
rect -1877 130 -1865 1106
rect -1831 130 -1819 1106
rect -1877 118 -1819 130
rect -1569 1106 -1511 1118
rect -1569 130 -1557 1106
rect -1523 130 -1511 1106
rect -1569 118 -1511 130
rect -1261 1106 -1203 1118
rect -1261 130 -1249 1106
rect -1215 130 -1203 1106
rect -1261 118 -1203 130
rect -953 1106 -895 1118
rect -953 130 -941 1106
rect -907 130 -895 1106
rect -953 118 -895 130
rect -645 1106 -587 1118
rect -645 130 -633 1106
rect -599 130 -587 1106
rect -645 118 -587 130
rect -337 1106 -279 1118
rect -337 130 -325 1106
rect -291 130 -279 1106
rect -337 118 -279 130
rect -29 1106 29 1118
rect -29 130 -17 1106
rect 17 130 29 1106
rect -29 118 29 130
rect 279 1106 337 1118
rect 279 130 291 1106
rect 325 130 337 1106
rect 279 118 337 130
rect 587 1106 645 1118
rect 587 130 599 1106
rect 633 130 645 1106
rect 587 118 645 130
rect 895 1106 953 1118
rect 895 130 907 1106
rect 941 130 953 1106
rect 895 118 953 130
rect 1203 1106 1261 1118
rect 1203 130 1215 1106
rect 1249 130 1261 1106
rect 1203 118 1261 130
rect 1511 1106 1569 1118
rect 1511 130 1523 1106
rect 1557 130 1569 1106
rect 1511 118 1569 130
rect 1819 1106 1877 1118
rect 1819 130 1831 1106
rect 1865 130 1877 1106
rect 1819 118 1877 130
rect 2127 1106 2185 1118
rect 2127 130 2139 1106
rect 2173 130 2185 1106
rect 2127 118 2185 130
rect 2435 1106 2493 1118
rect 2435 130 2447 1106
rect 2481 130 2493 1106
rect 2435 118 2493 130
rect -2493 -130 -2435 -118
rect -2493 -1106 -2481 -130
rect -2447 -1106 -2435 -130
rect -2493 -1118 -2435 -1106
rect -2185 -130 -2127 -118
rect -2185 -1106 -2173 -130
rect -2139 -1106 -2127 -130
rect -2185 -1118 -2127 -1106
rect -1877 -130 -1819 -118
rect -1877 -1106 -1865 -130
rect -1831 -1106 -1819 -130
rect -1877 -1118 -1819 -1106
rect -1569 -130 -1511 -118
rect -1569 -1106 -1557 -130
rect -1523 -1106 -1511 -130
rect -1569 -1118 -1511 -1106
rect -1261 -130 -1203 -118
rect -1261 -1106 -1249 -130
rect -1215 -1106 -1203 -130
rect -1261 -1118 -1203 -1106
rect -953 -130 -895 -118
rect -953 -1106 -941 -130
rect -907 -1106 -895 -130
rect -953 -1118 -895 -1106
rect -645 -130 -587 -118
rect -645 -1106 -633 -130
rect -599 -1106 -587 -130
rect -645 -1118 -587 -1106
rect -337 -130 -279 -118
rect -337 -1106 -325 -130
rect -291 -1106 -279 -130
rect -337 -1118 -279 -1106
rect -29 -130 29 -118
rect -29 -1106 -17 -130
rect 17 -1106 29 -130
rect -29 -1118 29 -1106
rect 279 -130 337 -118
rect 279 -1106 291 -130
rect 325 -1106 337 -130
rect 279 -1118 337 -1106
rect 587 -130 645 -118
rect 587 -1106 599 -130
rect 633 -1106 645 -130
rect 587 -1118 645 -1106
rect 895 -130 953 -118
rect 895 -1106 907 -130
rect 941 -1106 953 -130
rect 895 -1118 953 -1106
rect 1203 -130 1261 -118
rect 1203 -1106 1215 -130
rect 1249 -1106 1261 -130
rect 1203 -1118 1261 -1106
rect 1511 -130 1569 -118
rect 1511 -1106 1523 -130
rect 1557 -1106 1569 -130
rect 1511 -1118 1569 -1106
rect 1819 -130 1877 -118
rect 1819 -1106 1831 -130
rect 1865 -1106 1877 -130
rect 1819 -1118 1877 -1106
rect 2127 -130 2185 -118
rect 2127 -1106 2139 -130
rect 2173 -1106 2185 -130
rect 2127 -1118 2185 -1106
rect 2435 -130 2493 -118
rect 2435 -1106 2447 -130
rect 2481 -1106 2493 -130
rect 2435 -1118 2493 -1106
<< mvpdiffc >>
rect -2481 130 -2447 1106
rect -2173 130 -2139 1106
rect -1865 130 -1831 1106
rect -1557 130 -1523 1106
rect -1249 130 -1215 1106
rect -941 130 -907 1106
rect -633 130 -599 1106
rect -325 130 -291 1106
rect -17 130 17 1106
rect 291 130 325 1106
rect 599 130 633 1106
rect 907 130 941 1106
rect 1215 130 1249 1106
rect 1523 130 1557 1106
rect 1831 130 1865 1106
rect 2139 130 2173 1106
rect 2447 130 2481 1106
rect -2481 -1106 -2447 -130
rect -2173 -1106 -2139 -130
rect -1865 -1106 -1831 -130
rect -1557 -1106 -1523 -130
rect -1249 -1106 -1215 -130
rect -941 -1106 -907 -130
rect -633 -1106 -599 -130
rect -325 -1106 -291 -130
rect -17 -1106 17 -130
rect 291 -1106 325 -130
rect 599 -1106 633 -130
rect 907 -1106 941 -130
rect 1215 -1106 1249 -130
rect 1523 -1106 1557 -130
rect 1831 -1106 1865 -130
rect 2139 -1106 2173 -130
rect 2447 -1106 2481 -130
<< mvnsubdiff >>
rect -2627 1337 2627 1349
rect -2627 1303 -2519 1337
rect 2519 1303 2627 1337
rect -2627 1291 2627 1303
rect -2627 1241 -2569 1291
rect -2627 -1241 -2615 1241
rect -2581 -1241 -2569 1241
rect 2569 1241 2627 1291
rect -2627 -1291 -2569 -1241
rect 2569 -1241 2581 1241
rect 2615 -1241 2627 1241
rect 2569 -1291 2627 -1241
rect -2627 -1303 2627 -1291
rect -2627 -1337 -2519 -1303
rect 2519 -1337 2627 -1303
rect -2627 -1349 2627 -1337
<< mvnsubdiffcont >>
rect -2519 1303 2519 1337
rect -2615 -1241 -2581 1241
rect 2581 -1241 2615 1241
rect -2519 -1337 2519 -1303
<< poly >>
rect -2435 1199 -2185 1215
rect -2435 1165 -2419 1199
rect -2201 1165 -2185 1199
rect -2435 1118 -2185 1165
rect -2127 1199 -1877 1215
rect -2127 1165 -2111 1199
rect -1893 1165 -1877 1199
rect -2127 1118 -1877 1165
rect -1819 1199 -1569 1215
rect -1819 1165 -1803 1199
rect -1585 1165 -1569 1199
rect -1819 1118 -1569 1165
rect -1511 1199 -1261 1215
rect -1511 1165 -1495 1199
rect -1277 1165 -1261 1199
rect -1511 1118 -1261 1165
rect -1203 1199 -953 1215
rect -1203 1165 -1187 1199
rect -969 1165 -953 1199
rect -1203 1118 -953 1165
rect -895 1199 -645 1215
rect -895 1165 -879 1199
rect -661 1165 -645 1199
rect -895 1118 -645 1165
rect -587 1199 -337 1215
rect -587 1165 -571 1199
rect -353 1165 -337 1199
rect -587 1118 -337 1165
rect -279 1199 -29 1215
rect -279 1165 -263 1199
rect -45 1165 -29 1199
rect -279 1118 -29 1165
rect 29 1199 279 1215
rect 29 1165 45 1199
rect 263 1165 279 1199
rect 29 1118 279 1165
rect 337 1199 587 1215
rect 337 1165 353 1199
rect 571 1165 587 1199
rect 337 1118 587 1165
rect 645 1199 895 1215
rect 645 1165 661 1199
rect 879 1165 895 1199
rect 645 1118 895 1165
rect 953 1199 1203 1215
rect 953 1165 969 1199
rect 1187 1165 1203 1199
rect 953 1118 1203 1165
rect 1261 1199 1511 1215
rect 1261 1165 1277 1199
rect 1495 1165 1511 1199
rect 1261 1118 1511 1165
rect 1569 1199 1819 1215
rect 1569 1165 1585 1199
rect 1803 1165 1819 1199
rect 1569 1118 1819 1165
rect 1877 1199 2127 1215
rect 1877 1165 1893 1199
rect 2111 1165 2127 1199
rect 1877 1118 2127 1165
rect 2185 1199 2435 1215
rect 2185 1165 2201 1199
rect 2419 1165 2435 1199
rect 2185 1118 2435 1165
rect -2435 71 -2185 118
rect -2435 37 -2419 71
rect -2201 37 -2185 71
rect -2435 21 -2185 37
rect -2127 71 -1877 118
rect -2127 37 -2111 71
rect -1893 37 -1877 71
rect -2127 21 -1877 37
rect -1819 71 -1569 118
rect -1819 37 -1803 71
rect -1585 37 -1569 71
rect -1819 21 -1569 37
rect -1511 71 -1261 118
rect -1511 37 -1495 71
rect -1277 37 -1261 71
rect -1511 21 -1261 37
rect -1203 71 -953 118
rect -1203 37 -1187 71
rect -969 37 -953 71
rect -1203 21 -953 37
rect -895 71 -645 118
rect -895 37 -879 71
rect -661 37 -645 71
rect -895 21 -645 37
rect -587 71 -337 118
rect -587 37 -571 71
rect -353 37 -337 71
rect -587 21 -337 37
rect -279 71 -29 118
rect -279 37 -263 71
rect -45 37 -29 71
rect -279 21 -29 37
rect 29 71 279 118
rect 29 37 45 71
rect 263 37 279 71
rect 29 21 279 37
rect 337 71 587 118
rect 337 37 353 71
rect 571 37 587 71
rect 337 21 587 37
rect 645 71 895 118
rect 645 37 661 71
rect 879 37 895 71
rect 645 21 895 37
rect 953 71 1203 118
rect 953 37 969 71
rect 1187 37 1203 71
rect 953 21 1203 37
rect 1261 71 1511 118
rect 1261 37 1277 71
rect 1495 37 1511 71
rect 1261 21 1511 37
rect 1569 71 1819 118
rect 1569 37 1585 71
rect 1803 37 1819 71
rect 1569 21 1819 37
rect 1877 71 2127 118
rect 1877 37 1893 71
rect 2111 37 2127 71
rect 1877 21 2127 37
rect 2185 71 2435 118
rect 2185 37 2201 71
rect 2419 37 2435 71
rect 2185 21 2435 37
rect -2435 -37 -2185 -21
rect -2435 -71 -2419 -37
rect -2201 -71 -2185 -37
rect -2435 -118 -2185 -71
rect -2127 -37 -1877 -21
rect -2127 -71 -2111 -37
rect -1893 -71 -1877 -37
rect -2127 -118 -1877 -71
rect -1819 -37 -1569 -21
rect -1819 -71 -1803 -37
rect -1585 -71 -1569 -37
rect -1819 -118 -1569 -71
rect -1511 -37 -1261 -21
rect -1511 -71 -1495 -37
rect -1277 -71 -1261 -37
rect -1511 -118 -1261 -71
rect -1203 -37 -953 -21
rect -1203 -71 -1187 -37
rect -969 -71 -953 -37
rect -1203 -118 -953 -71
rect -895 -37 -645 -21
rect -895 -71 -879 -37
rect -661 -71 -645 -37
rect -895 -118 -645 -71
rect -587 -37 -337 -21
rect -587 -71 -571 -37
rect -353 -71 -337 -37
rect -587 -118 -337 -71
rect -279 -37 -29 -21
rect -279 -71 -263 -37
rect -45 -71 -29 -37
rect -279 -118 -29 -71
rect 29 -37 279 -21
rect 29 -71 45 -37
rect 263 -71 279 -37
rect 29 -118 279 -71
rect 337 -37 587 -21
rect 337 -71 353 -37
rect 571 -71 587 -37
rect 337 -118 587 -71
rect 645 -37 895 -21
rect 645 -71 661 -37
rect 879 -71 895 -37
rect 645 -118 895 -71
rect 953 -37 1203 -21
rect 953 -71 969 -37
rect 1187 -71 1203 -37
rect 953 -118 1203 -71
rect 1261 -37 1511 -21
rect 1261 -71 1277 -37
rect 1495 -71 1511 -37
rect 1261 -118 1511 -71
rect 1569 -37 1819 -21
rect 1569 -71 1585 -37
rect 1803 -71 1819 -37
rect 1569 -118 1819 -71
rect 1877 -37 2127 -21
rect 1877 -71 1893 -37
rect 2111 -71 2127 -37
rect 1877 -118 2127 -71
rect 2185 -37 2435 -21
rect 2185 -71 2201 -37
rect 2419 -71 2435 -37
rect 2185 -118 2435 -71
rect -2435 -1165 -2185 -1118
rect -2435 -1199 -2419 -1165
rect -2201 -1199 -2185 -1165
rect -2435 -1215 -2185 -1199
rect -2127 -1165 -1877 -1118
rect -2127 -1199 -2111 -1165
rect -1893 -1199 -1877 -1165
rect -2127 -1215 -1877 -1199
rect -1819 -1165 -1569 -1118
rect -1819 -1199 -1803 -1165
rect -1585 -1199 -1569 -1165
rect -1819 -1215 -1569 -1199
rect -1511 -1165 -1261 -1118
rect -1511 -1199 -1495 -1165
rect -1277 -1199 -1261 -1165
rect -1511 -1215 -1261 -1199
rect -1203 -1165 -953 -1118
rect -1203 -1199 -1187 -1165
rect -969 -1199 -953 -1165
rect -1203 -1215 -953 -1199
rect -895 -1165 -645 -1118
rect -895 -1199 -879 -1165
rect -661 -1199 -645 -1165
rect -895 -1215 -645 -1199
rect -587 -1165 -337 -1118
rect -587 -1199 -571 -1165
rect -353 -1199 -337 -1165
rect -587 -1215 -337 -1199
rect -279 -1165 -29 -1118
rect -279 -1199 -263 -1165
rect -45 -1199 -29 -1165
rect -279 -1215 -29 -1199
rect 29 -1165 279 -1118
rect 29 -1199 45 -1165
rect 263 -1199 279 -1165
rect 29 -1215 279 -1199
rect 337 -1165 587 -1118
rect 337 -1199 353 -1165
rect 571 -1199 587 -1165
rect 337 -1215 587 -1199
rect 645 -1165 895 -1118
rect 645 -1199 661 -1165
rect 879 -1199 895 -1165
rect 645 -1215 895 -1199
rect 953 -1165 1203 -1118
rect 953 -1199 969 -1165
rect 1187 -1199 1203 -1165
rect 953 -1215 1203 -1199
rect 1261 -1165 1511 -1118
rect 1261 -1199 1277 -1165
rect 1495 -1199 1511 -1165
rect 1261 -1215 1511 -1199
rect 1569 -1165 1819 -1118
rect 1569 -1199 1585 -1165
rect 1803 -1199 1819 -1165
rect 1569 -1215 1819 -1199
rect 1877 -1165 2127 -1118
rect 1877 -1199 1893 -1165
rect 2111 -1199 2127 -1165
rect 1877 -1215 2127 -1199
rect 2185 -1165 2435 -1118
rect 2185 -1199 2201 -1165
rect 2419 -1199 2435 -1165
rect 2185 -1215 2435 -1199
<< polycont >>
rect -2419 1165 -2201 1199
rect -2111 1165 -1893 1199
rect -1803 1165 -1585 1199
rect -1495 1165 -1277 1199
rect -1187 1165 -969 1199
rect -879 1165 -661 1199
rect -571 1165 -353 1199
rect -263 1165 -45 1199
rect 45 1165 263 1199
rect 353 1165 571 1199
rect 661 1165 879 1199
rect 969 1165 1187 1199
rect 1277 1165 1495 1199
rect 1585 1165 1803 1199
rect 1893 1165 2111 1199
rect 2201 1165 2419 1199
rect -2419 37 -2201 71
rect -2111 37 -1893 71
rect -1803 37 -1585 71
rect -1495 37 -1277 71
rect -1187 37 -969 71
rect -879 37 -661 71
rect -571 37 -353 71
rect -263 37 -45 71
rect 45 37 263 71
rect 353 37 571 71
rect 661 37 879 71
rect 969 37 1187 71
rect 1277 37 1495 71
rect 1585 37 1803 71
rect 1893 37 2111 71
rect 2201 37 2419 71
rect -2419 -71 -2201 -37
rect -2111 -71 -1893 -37
rect -1803 -71 -1585 -37
rect -1495 -71 -1277 -37
rect -1187 -71 -969 -37
rect -879 -71 -661 -37
rect -571 -71 -353 -37
rect -263 -71 -45 -37
rect 45 -71 263 -37
rect 353 -71 571 -37
rect 661 -71 879 -37
rect 969 -71 1187 -37
rect 1277 -71 1495 -37
rect 1585 -71 1803 -37
rect 1893 -71 2111 -37
rect 2201 -71 2419 -37
rect -2419 -1199 -2201 -1165
rect -2111 -1199 -1893 -1165
rect -1803 -1199 -1585 -1165
rect -1495 -1199 -1277 -1165
rect -1187 -1199 -969 -1165
rect -879 -1199 -661 -1165
rect -571 -1199 -353 -1165
rect -263 -1199 -45 -1165
rect 45 -1199 263 -1165
rect 353 -1199 571 -1165
rect 661 -1199 879 -1165
rect 969 -1199 1187 -1165
rect 1277 -1199 1495 -1165
rect 1585 -1199 1803 -1165
rect 1893 -1199 2111 -1165
rect 2201 -1199 2419 -1165
<< locali >>
rect -2615 1303 -2519 1337
rect 2519 1303 2615 1337
rect -2615 1241 -2581 1303
rect 2581 1241 2615 1303
rect -2435 1165 -2419 1199
rect -2201 1165 -2185 1199
rect -2127 1165 -2111 1199
rect -1893 1165 -1877 1199
rect -1819 1165 -1803 1199
rect -1585 1165 -1569 1199
rect -1511 1165 -1495 1199
rect -1277 1165 -1261 1199
rect -1203 1165 -1187 1199
rect -969 1165 -953 1199
rect -895 1165 -879 1199
rect -661 1165 -645 1199
rect -587 1165 -571 1199
rect -353 1165 -337 1199
rect -279 1165 -263 1199
rect -45 1165 -29 1199
rect 29 1165 45 1199
rect 263 1165 279 1199
rect 337 1165 353 1199
rect 571 1165 587 1199
rect 645 1165 661 1199
rect 879 1165 895 1199
rect 953 1165 969 1199
rect 1187 1165 1203 1199
rect 1261 1165 1277 1199
rect 1495 1165 1511 1199
rect 1569 1165 1585 1199
rect 1803 1165 1819 1199
rect 1877 1165 1893 1199
rect 2111 1165 2127 1199
rect 2185 1165 2201 1199
rect 2419 1165 2435 1199
rect -2481 1106 -2447 1122
rect -2481 114 -2447 130
rect -2173 1106 -2139 1122
rect -2173 114 -2139 130
rect -1865 1106 -1831 1122
rect -1865 114 -1831 130
rect -1557 1106 -1523 1122
rect -1557 114 -1523 130
rect -1249 1106 -1215 1122
rect -1249 114 -1215 130
rect -941 1106 -907 1122
rect -941 114 -907 130
rect -633 1106 -599 1122
rect -633 114 -599 130
rect -325 1106 -291 1122
rect -325 114 -291 130
rect -17 1106 17 1122
rect -17 114 17 130
rect 291 1106 325 1122
rect 291 114 325 130
rect 599 1106 633 1122
rect 599 114 633 130
rect 907 1106 941 1122
rect 907 114 941 130
rect 1215 1106 1249 1122
rect 1215 114 1249 130
rect 1523 1106 1557 1122
rect 1523 114 1557 130
rect 1831 1106 1865 1122
rect 1831 114 1865 130
rect 2139 1106 2173 1122
rect 2139 114 2173 130
rect 2447 1106 2481 1122
rect 2447 114 2481 130
rect -2435 37 -2419 71
rect -2201 37 -2185 71
rect -2127 37 -2111 71
rect -1893 37 -1877 71
rect -1819 37 -1803 71
rect -1585 37 -1569 71
rect -1511 37 -1495 71
rect -1277 37 -1261 71
rect -1203 37 -1187 71
rect -969 37 -953 71
rect -895 37 -879 71
rect -661 37 -645 71
rect -587 37 -571 71
rect -353 37 -337 71
rect -279 37 -263 71
rect -45 37 -29 71
rect 29 37 45 71
rect 263 37 279 71
rect 337 37 353 71
rect 571 37 587 71
rect 645 37 661 71
rect 879 37 895 71
rect 953 37 969 71
rect 1187 37 1203 71
rect 1261 37 1277 71
rect 1495 37 1511 71
rect 1569 37 1585 71
rect 1803 37 1819 71
rect 1877 37 1893 71
rect 2111 37 2127 71
rect 2185 37 2201 71
rect 2419 37 2435 71
rect -2435 -71 -2419 -37
rect -2201 -71 -2185 -37
rect -2127 -71 -2111 -37
rect -1893 -71 -1877 -37
rect -1819 -71 -1803 -37
rect -1585 -71 -1569 -37
rect -1511 -71 -1495 -37
rect -1277 -71 -1261 -37
rect -1203 -71 -1187 -37
rect -969 -71 -953 -37
rect -895 -71 -879 -37
rect -661 -71 -645 -37
rect -587 -71 -571 -37
rect -353 -71 -337 -37
rect -279 -71 -263 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 263 -71 279 -37
rect 337 -71 353 -37
rect 571 -71 587 -37
rect 645 -71 661 -37
rect 879 -71 895 -37
rect 953 -71 969 -37
rect 1187 -71 1203 -37
rect 1261 -71 1277 -37
rect 1495 -71 1511 -37
rect 1569 -71 1585 -37
rect 1803 -71 1819 -37
rect 1877 -71 1893 -37
rect 2111 -71 2127 -37
rect 2185 -71 2201 -37
rect 2419 -71 2435 -37
rect -2481 -130 -2447 -114
rect -2481 -1122 -2447 -1106
rect -2173 -130 -2139 -114
rect -2173 -1122 -2139 -1106
rect -1865 -130 -1831 -114
rect -1865 -1122 -1831 -1106
rect -1557 -130 -1523 -114
rect -1557 -1122 -1523 -1106
rect -1249 -130 -1215 -114
rect -1249 -1122 -1215 -1106
rect -941 -130 -907 -114
rect -941 -1122 -907 -1106
rect -633 -130 -599 -114
rect -633 -1122 -599 -1106
rect -325 -130 -291 -114
rect -325 -1122 -291 -1106
rect -17 -130 17 -114
rect -17 -1122 17 -1106
rect 291 -130 325 -114
rect 291 -1122 325 -1106
rect 599 -130 633 -114
rect 599 -1122 633 -1106
rect 907 -130 941 -114
rect 907 -1122 941 -1106
rect 1215 -130 1249 -114
rect 1215 -1122 1249 -1106
rect 1523 -130 1557 -114
rect 1523 -1122 1557 -1106
rect 1831 -130 1865 -114
rect 1831 -1122 1865 -1106
rect 2139 -130 2173 -114
rect 2139 -1122 2173 -1106
rect 2447 -130 2481 -114
rect 2447 -1122 2481 -1106
rect -2435 -1199 -2419 -1165
rect -2201 -1199 -2185 -1165
rect -2127 -1199 -2111 -1165
rect -1893 -1199 -1877 -1165
rect -1819 -1199 -1803 -1165
rect -1585 -1199 -1569 -1165
rect -1511 -1199 -1495 -1165
rect -1277 -1199 -1261 -1165
rect -1203 -1199 -1187 -1165
rect -969 -1199 -953 -1165
rect -895 -1199 -879 -1165
rect -661 -1199 -645 -1165
rect -587 -1199 -571 -1165
rect -353 -1199 -337 -1165
rect -279 -1199 -263 -1165
rect -45 -1199 -29 -1165
rect 29 -1199 45 -1165
rect 263 -1199 279 -1165
rect 337 -1199 353 -1165
rect 571 -1199 587 -1165
rect 645 -1199 661 -1165
rect 879 -1199 895 -1165
rect 953 -1199 969 -1165
rect 1187 -1199 1203 -1165
rect 1261 -1199 1277 -1165
rect 1495 -1199 1511 -1165
rect 1569 -1199 1585 -1165
rect 1803 -1199 1819 -1165
rect 1877 -1199 1893 -1165
rect 2111 -1199 2127 -1165
rect 2185 -1199 2201 -1165
rect 2419 -1199 2435 -1165
rect -2615 -1303 -2581 -1241
rect 2581 -1303 2615 -1241
rect -2615 -1337 -2519 -1303
rect 2519 -1337 2615 -1303
<< viali >>
rect -2419 1165 -2201 1199
rect -2111 1165 -1893 1199
rect -1803 1165 -1585 1199
rect -1495 1165 -1277 1199
rect -1187 1165 -969 1199
rect -879 1165 -661 1199
rect -571 1165 -353 1199
rect -263 1165 -45 1199
rect 45 1165 263 1199
rect 353 1165 571 1199
rect 661 1165 879 1199
rect 969 1165 1187 1199
rect 1277 1165 1495 1199
rect 1585 1165 1803 1199
rect 1893 1165 2111 1199
rect 2201 1165 2419 1199
rect -2481 130 -2447 1106
rect -2173 130 -2139 1106
rect -1865 130 -1831 1106
rect -1557 130 -1523 1106
rect -1249 130 -1215 1106
rect -941 130 -907 1106
rect -633 130 -599 1106
rect -325 130 -291 1106
rect -17 130 17 1106
rect 291 130 325 1106
rect 599 130 633 1106
rect 907 130 941 1106
rect 1215 130 1249 1106
rect 1523 130 1557 1106
rect 1831 130 1865 1106
rect 2139 130 2173 1106
rect 2447 130 2481 1106
rect -2419 37 -2201 71
rect -2111 37 -1893 71
rect -1803 37 -1585 71
rect -1495 37 -1277 71
rect -1187 37 -969 71
rect -879 37 -661 71
rect -571 37 -353 71
rect -263 37 -45 71
rect 45 37 263 71
rect 353 37 571 71
rect 661 37 879 71
rect 969 37 1187 71
rect 1277 37 1495 71
rect 1585 37 1803 71
rect 1893 37 2111 71
rect 2201 37 2419 71
rect -2419 -71 -2201 -37
rect -2111 -71 -1893 -37
rect -1803 -71 -1585 -37
rect -1495 -71 -1277 -37
rect -1187 -71 -969 -37
rect -879 -71 -661 -37
rect -571 -71 -353 -37
rect -263 -71 -45 -37
rect 45 -71 263 -37
rect 353 -71 571 -37
rect 661 -71 879 -37
rect 969 -71 1187 -37
rect 1277 -71 1495 -37
rect 1585 -71 1803 -37
rect 1893 -71 2111 -37
rect 2201 -71 2419 -37
rect -2481 -1106 -2447 -130
rect -2173 -1106 -2139 -130
rect -1865 -1106 -1831 -130
rect -1557 -1106 -1523 -130
rect -1249 -1106 -1215 -130
rect -941 -1106 -907 -130
rect -633 -1106 -599 -130
rect -325 -1106 -291 -130
rect -17 -1106 17 -130
rect 291 -1106 325 -130
rect 599 -1106 633 -130
rect 907 -1106 941 -130
rect 1215 -1106 1249 -130
rect 1523 -1106 1557 -130
rect 1831 -1106 1865 -130
rect 2139 -1106 2173 -130
rect 2447 -1106 2481 -130
rect -2419 -1199 -2201 -1165
rect -2111 -1199 -1893 -1165
rect -1803 -1199 -1585 -1165
rect -1495 -1199 -1277 -1165
rect -1187 -1199 -969 -1165
rect -879 -1199 -661 -1165
rect -571 -1199 -353 -1165
rect -263 -1199 -45 -1165
rect 45 -1199 263 -1165
rect 353 -1199 571 -1165
rect 661 -1199 879 -1165
rect 969 -1199 1187 -1165
rect 1277 -1199 1495 -1165
rect 1585 -1199 1803 -1165
rect 1893 -1199 2111 -1165
rect 2201 -1199 2419 -1165
<< metal1 >>
rect -2431 1199 -2189 1205
rect -2431 1165 -2419 1199
rect -2201 1165 -2189 1199
rect -2431 1159 -2189 1165
rect -2123 1199 -1881 1205
rect -2123 1165 -2111 1199
rect -1893 1165 -1881 1199
rect -2123 1159 -1881 1165
rect -1815 1199 -1573 1205
rect -1815 1165 -1803 1199
rect -1585 1165 -1573 1199
rect -1815 1159 -1573 1165
rect -1507 1199 -1265 1205
rect -1507 1165 -1495 1199
rect -1277 1165 -1265 1199
rect -1507 1159 -1265 1165
rect -1199 1199 -957 1205
rect -1199 1165 -1187 1199
rect -969 1165 -957 1199
rect -1199 1159 -957 1165
rect -891 1199 -649 1205
rect -891 1165 -879 1199
rect -661 1165 -649 1199
rect -891 1159 -649 1165
rect -583 1199 -341 1205
rect -583 1165 -571 1199
rect -353 1165 -341 1199
rect -583 1159 -341 1165
rect -275 1199 -33 1205
rect -275 1165 -263 1199
rect -45 1165 -33 1199
rect -275 1159 -33 1165
rect 33 1199 275 1205
rect 33 1165 45 1199
rect 263 1165 275 1199
rect 33 1159 275 1165
rect 341 1199 583 1205
rect 341 1165 353 1199
rect 571 1165 583 1199
rect 341 1159 583 1165
rect 649 1199 891 1205
rect 649 1165 661 1199
rect 879 1165 891 1199
rect 649 1159 891 1165
rect 957 1199 1199 1205
rect 957 1165 969 1199
rect 1187 1165 1199 1199
rect 957 1159 1199 1165
rect 1265 1199 1507 1205
rect 1265 1165 1277 1199
rect 1495 1165 1507 1199
rect 1265 1159 1507 1165
rect 1573 1199 1815 1205
rect 1573 1165 1585 1199
rect 1803 1165 1815 1199
rect 1573 1159 1815 1165
rect 1881 1199 2123 1205
rect 1881 1165 1893 1199
rect 2111 1165 2123 1199
rect 1881 1159 2123 1165
rect 2189 1199 2431 1205
rect 2189 1165 2201 1199
rect 2419 1165 2431 1199
rect 2189 1159 2431 1165
rect -2487 1106 -2441 1118
rect -2487 130 -2481 1106
rect -2447 130 -2441 1106
rect -2487 118 -2441 130
rect -2179 1106 -2133 1118
rect -2179 130 -2173 1106
rect -2139 130 -2133 1106
rect -2179 118 -2133 130
rect -1871 1106 -1825 1118
rect -1871 130 -1865 1106
rect -1831 130 -1825 1106
rect -1871 118 -1825 130
rect -1563 1106 -1517 1118
rect -1563 130 -1557 1106
rect -1523 130 -1517 1106
rect -1563 118 -1517 130
rect -1255 1106 -1209 1118
rect -1255 130 -1249 1106
rect -1215 130 -1209 1106
rect -1255 118 -1209 130
rect -947 1106 -901 1118
rect -947 130 -941 1106
rect -907 130 -901 1106
rect -947 118 -901 130
rect -639 1106 -593 1118
rect -639 130 -633 1106
rect -599 130 -593 1106
rect -639 118 -593 130
rect -331 1106 -285 1118
rect -331 130 -325 1106
rect -291 130 -285 1106
rect -331 118 -285 130
rect -23 1106 23 1118
rect -23 130 -17 1106
rect 17 130 23 1106
rect -23 118 23 130
rect 285 1106 331 1118
rect 285 130 291 1106
rect 325 130 331 1106
rect 285 118 331 130
rect 593 1106 639 1118
rect 593 130 599 1106
rect 633 130 639 1106
rect 593 118 639 130
rect 901 1106 947 1118
rect 901 130 907 1106
rect 941 130 947 1106
rect 901 118 947 130
rect 1209 1106 1255 1118
rect 1209 130 1215 1106
rect 1249 130 1255 1106
rect 1209 118 1255 130
rect 1517 1106 1563 1118
rect 1517 130 1523 1106
rect 1557 130 1563 1106
rect 1517 118 1563 130
rect 1825 1106 1871 1118
rect 1825 130 1831 1106
rect 1865 130 1871 1106
rect 1825 118 1871 130
rect 2133 1106 2179 1118
rect 2133 130 2139 1106
rect 2173 130 2179 1106
rect 2133 118 2179 130
rect 2441 1106 2487 1118
rect 2441 130 2447 1106
rect 2481 130 2487 1106
rect 2441 118 2487 130
rect -2431 71 -2189 77
rect -2431 37 -2419 71
rect -2201 37 -2189 71
rect -2431 31 -2189 37
rect -2123 71 -1881 77
rect -2123 37 -2111 71
rect -1893 37 -1881 71
rect -2123 31 -1881 37
rect -1815 71 -1573 77
rect -1815 37 -1803 71
rect -1585 37 -1573 71
rect -1815 31 -1573 37
rect -1507 71 -1265 77
rect -1507 37 -1495 71
rect -1277 37 -1265 71
rect -1507 31 -1265 37
rect -1199 71 -957 77
rect -1199 37 -1187 71
rect -969 37 -957 71
rect -1199 31 -957 37
rect -891 71 -649 77
rect -891 37 -879 71
rect -661 37 -649 71
rect -891 31 -649 37
rect -583 71 -341 77
rect -583 37 -571 71
rect -353 37 -341 71
rect -583 31 -341 37
rect -275 71 -33 77
rect -275 37 -263 71
rect -45 37 -33 71
rect -275 31 -33 37
rect 33 71 275 77
rect 33 37 45 71
rect 263 37 275 71
rect 33 31 275 37
rect 341 71 583 77
rect 341 37 353 71
rect 571 37 583 71
rect 341 31 583 37
rect 649 71 891 77
rect 649 37 661 71
rect 879 37 891 71
rect 649 31 891 37
rect 957 71 1199 77
rect 957 37 969 71
rect 1187 37 1199 71
rect 957 31 1199 37
rect 1265 71 1507 77
rect 1265 37 1277 71
rect 1495 37 1507 71
rect 1265 31 1507 37
rect 1573 71 1815 77
rect 1573 37 1585 71
rect 1803 37 1815 71
rect 1573 31 1815 37
rect 1881 71 2123 77
rect 1881 37 1893 71
rect 2111 37 2123 71
rect 1881 31 2123 37
rect 2189 71 2431 77
rect 2189 37 2201 71
rect 2419 37 2431 71
rect 2189 31 2431 37
rect -2431 -37 -2189 -31
rect -2431 -71 -2419 -37
rect -2201 -71 -2189 -37
rect -2431 -77 -2189 -71
rect -2123 -37 -1881 -31
rect -2123 -71 -2111 -37
rect -1893 -71 -1881 -37
rect -2123 -77 -1881 -71
rect -1815 -37 -1573 -31
rect -1815 -71 -1803 -37
rect -1585 -71 -1573 -37
rect -1815 -77 -1573 -71
rect -1507 -37 -1265 -31
rect -1507 -71 -1495 -37
rect -1277 -71 -1265 -37
rect -1507 -77 -1265 -71
rect -1199 -37 -957 -31
rect -1199 -71 -1187 -37
rect -969 -71 -957 -37
rect -1199 -77 -957 -71
rect -891 -37 -649 -31
rect -891 -71 -879 -37
rect -661 -71 -649 -37
rect -891 -77 -649 -71
rect -583 -37 -341 -31
rect -583 -71 -571 -37
rect -353 -71 -341 -37
rect -583 -77 -341 -71
rect -275 -37 -33 -31
rect -275 -71 -263 -37
rect -45 -71 -33 -37
rect -275 -77 -33 -71
rect 33 -37 275 -31
rect 33 -71 45 -37
rect 263 -71 275 -37
rect 33 -77 275 -71
rect 341 -37 583 -31
rect 341 -71 353 -37
rect 571 -71 583 -37
rect 341 -77 583 -71
rect 649 -37 891 -31
rect 649 -71 661 -37
rect 879 -71 891 -37
rect 649 -77 891 -71
rect 957 -37 1199 -31
rect 957 -71 969 -37
rect 1187 -71 1199 -37
rect 957 -77 1199 -71
rect 1265 -37 1507 -31
rect 1265 -71 1277 -37
rect 1495 -71 1507 -37
rect 1265 -77 1507 -71
rect 1573 -37 1815 -31
rect 1573 -71 1585 -37
rect 1803 -71 1815 -37
rect 1573 -77 1815 -71
rect 1881 -37 2123 -31
rect 1881 -71 1893 -37
rect 2111 -71 2123 -37
rect 1881 -77 2123 -71
rect 2189 -37 2431 -31
rect 2189 -71 2201 -37
rect 2419 -71 2431 -37
rect 2189 -77 2431 -71
rect -2487 -130 -2441 -118
rect -2487 -1106 -2481 -130
rect -2447 -1106 -2441 -130
rect -2487 -1118 -2441 -1106
rect -2179 -130 -2133 -118
rect -2179 -1106 -2173 -130
rect -2139 -1106 -2133 -130
rect -2179 -1118 -2133 -1106
rect -1871 -130 -1825 -118
rect -1871 -1106 -1865 -130
rect -1831 -1106 -1825 -130
rect -1871 -1118 -1825 -1106
rect -1563 -130 -1517 -118
rect -1563 -1106 -1557 -130
rect -1523 -1106 -1517 -130
rect -1563 -1118 -1517 -1106
rect -1255 -130 -1209 -118
rect -1255 -1106 -1249 -130
rect -1215 -1106 -1209 -130
rect -1255 -1118 -1209 -1106
rect -947 -130 -901 -118
rect -947 -1106 -941 -130
rect -907 -1106 -901 -130
rect -947 -1118 -901 -1106
rect -639 -130 -593 -118
rect -639 -1106 -633 -130
rect -599 -1106 -593 -130
rect -639 -1118 -593 -1106
rect -331 -130 -285 -118
rect -331 -1106 -325 -130
rect -291 -1106 -285 -130
rect -331 -1118 -285 -1106
rect -23 -130 23 -118
rect -23 -1106 -17 -130
rect 17 -1106 23 -130
rect -23 -1118 23 -1106
rect 285 -130 331 -118
rect 285 -1106 291 -130
rect 325 -1106 331 -130
rect 285 -1118 331 -1106
rect 593 -130 639 -118
rect 593 -1106 599 -130
rect 633 -1106 639 -130
rect 593 -1118 639 -1106
rect 901 -130 947 -118
rect 901 -1106 907 -130
rect 941 -1106 947 -130
rect 901 -1118 947 -1106
rect 1209 -130 1255 -118
rect 1209 -1106 1215 -130
rect 1249 -1106 1255 -130
rect 1209 -1118 1255 -1106
rect 1517 -130 1563 -118
rect 1517 -1106 1523 -130
rect 1557 -1106 1563 -130
rect 1517 -1118 1563 -1106
rect 1825 -130 1871 -118
rect 1825 -1106 1831 -130
rect 1865 -1106 1871 -130
rect 1825 -1118 1871 -1106
rect 2133 -130 2179 -118
rect 2133 -1106 2139 -130
rect 2173 -1106 2179 -130
rect 2133 -1118 2179 -1106
rect 2441 -130 2487 -118
rect 2441 -1106 2447 -130
rect 2481 -1106 2487 -130
rect 2441 -1118 2487 -1106
rect -2431 -1165 -2189 -1159
rect -2431 -1199 -2419 -1165
rect -2201 -1199 -2189 -1165
rect -2431 -1205 -2189 -1199
rect -2123 -1165 -1881 -1159
rect -2123 -1199 -2111 -1165
rect -1893 -1199 -1881 -1165
rect -2123 -1205 -1881 -1199
rect -1815 -1165 -1573 -1159
rect -1815 -1199 -1803 -1165
rect -1585 -1199 -1573 -1165
rect -1815 -1205 -1573 -1199
rect -1507 -1165 -1265 -1159
rect -1507 -1199 -1495 -1165
rect -1277 -1199 -1265 -1165
rect -1507 -1205 -1265 -1199
rect -1199 -1165 -957 -1159
rect -1199 -1199 -1187 -1165
rect -969 -1199 -957 -1165
rect -1199 -1205 -957 -1199
rect -891 -1165 -649 -1159
rect -891 -1199 -879 -1165
rect -661 -1199 -649 -1165
rect -891 -1205 -649 -1199
rect -583 -1165 -341 -1159
rect -583 -1199 -571 -1165
rect -353 -1199 -341 -1165
rect -583 -1205 -341 -1199
rect -275 -1165 -33 -1159
rect -275 -1199 -263 -1165
rect -45 -1199 -33 -1165
rect -275 -1205 -33 -1199
rect 33 -1165 275 -1159
rect 33 -1199 45 -1165
rect 263 -1199 275 -1165
rect 33 -1205 275 -1199
rect 341 -1165 583 -1159
rect 341 -1199 353 -1165
rect 571 -1199 583 -1165
rect 341 -1205 583 -1199
rect 649 -1165 891 -1159
rect 649 -1199 661 -1165
rect 879 -1199 891 -1165
rect 649 -1205 891 -1199
rect 957 -1165 1199 -1159
rect 957 -1199 969 -1165
rect 1187 -1199 1199 -1165
rect 957 -1205 1199 -1199
rect 1265 -1165 1507 -1159
rect 1265 -1199 1277 -1165
rect 1495 -1199 1507 -1165
rect 1265 -1205 1507 -1199
rect 1573 -1165 1815 -1159
rect 1573 -1199 1585 -1165
rect 1803 -1199 1815 -1165
rect 1573 -1205 1815 -1199
rect 1881 -1165 2123 -1159
rect 1881 -1199 1893 -1165
rect 2111 -1199 2123 -1165
rect 1881 -1205 2123 -1199
rect 2189 -1165 2431 -1159
rect 2189 -1199 2201 -1165
rect 2419 -1199 2431 -1165
rect 2189 -1205 2431 -1199
<< properties >>
string FIXED_BBOX -2598 -1320 2598 1320
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.25 m 2 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
