magic
tech sky130A
timestamp 1770177229
<< psubdiff >>
rect -750 -2875 5000 -2750
rect -750 -3125 375 -2875
rect 3875 -3125 5000 -2875
rect -750 -3250 5000 -3125
rect -750 -35750 -250 -3250
rect 3750 -15900 4250 -15750
rect 3750 -16100 3900 -15900
rect 4100 -16100 4250 -15900
rect 3750 -16250 4250 -16100
rect 4500 -35750 5000 -3250
rect -750 -35875 5000 -35750
rect -750 -36125 375 -35875
rect 3875 -36125 5000 -35875
rect -750 -36250 5000 -36125
<< psubdiffcont >>
rect 375 -3125 3875 -2875
rect 3900 -16100 4100 -15900
rect 375 -36125 3875 -35875
<< xpolycontact >>
rect 0 -4000 500 -3500
rect 0 -35500 500 -35000
<< xpolyres >>
rect 500 -4000 4250 -3500
rect 3750 -7000 4250 -4000
rect 0 -7500 4250 -7000
rect 0 -10500 500 -7500
rect 0 -11000 4250 -10500
rect 3750 -14000 4250 -11000
rect 0 -14500 4250 -14000
rect 0 -17500 500 -14500
rect 0 -18000 4250 -17500
rect 3750 -21000 4250 -18000
rect 0 -21500 4250 -21000
rect 0 -24500 500 -21500
rect 0 -25000 4250 -24500
rect 3750 -28000 4250 -25000
rect 0 -28500 4250 -28000
rect 0 -31500 500 -28500
rect 0 -32000 4250 -31500
rect 3750 -35000 4250 -32000
rect 500 -35500 4250 -35000
<< locali >>
rect -750 -2875 5000 -2750
rect -750 -3125 375 -2875
rect 3875 -3125 5000 -2875
rect -750 -3250 5000 -3125
rect -750 -35750 -250 -3250
rect 3800 -15900 4200 -15800
rect 3800 -16100 3900 -15900
rect 4100 -16100 4200 -15900
rect 3800 -16200 4200 -16100
rect 4500 -35750 5000 -3250
rect -750 -35875 5000 -35750
rect -750 -36125 375 -35875
rect 3875 -36125 5000 -35875
rect -750 -36250 5000 -36125
<< viali >>
rect 3900 -16100 4100 -15900
<< metal1 >>
rect 3800 -15900 4200 -15800
rect 3800 -16100 3900 -15900
rect 4100 -16100 4200 -15900
rect 3800 -16200 4200 -16100
<< labels >>
rlabel xpolycontact 250 -3500 250 -3500 1 A
rlabel space 0 -35750 500 -35500 1 B
rlabel space 4250 -16000 4250 -16000 3 VSS
<< end >>
