magic
tech sky130A
magscale 1 2
timestamp 1769077132
<< mvnmos >>
rect -467 -177 -367 239
rect -189 -177 -89 239
rect 89 -177 189 239
rect 367 -177 467 239
<< mvndiff >>
rect -525 227 -467 239
rect -525 -165 -513 227
rect -479 -165 -467 227
rect -525 -177 -467 -165
rect -367 227 -309 239
rect -367 -165 -355 227
rect -321 -165 -309 227
rect -367 -177 -309 -165
rect -247 227 -189 239
rect -247 -165 -235 227
rect -201 -165 -189 227
rect -247 -177 -189 -165
rect -89 227 -31 239
rect -89 -165 -77 227
rect -43 -165 -31 227
rect -89 -177 -31 -165
rect 31 227 89 239
rect 31 -165 43 227
rect 77 -165 89 227
rect 31 -177 89 -165
rect 189 227 247 239
rect 189 -165 201 227
rect 235 -165 247 227
rect 189 -177 247 -165
rect 309 227 367 239
rect 309 -165 321 227
rect 355 -165 367 227
rect 309 -177 367 -165
rect 467 227 525 239
rect 467 -165 479 227
rect 513 -165 525 227
rect 467 -177 525 -165
<< mvndiffc >>
rect -513 -165 -479 227
rect -355 -165 -321 227
rect -235 -165 -201 227
rect -77 -165 -43 227
rect 43 -165 77 227
rect 201 -165 235 227
rect 321 -165 355 227
rect 479 -165 513 227
<< poly >>
rect -467 239 -367 265
rect -189 239 -89 265
rect 89 239 189 265
rect 367 239 467 265
rect -467 -215 -367 -177
rect -467 -249 -451 -215
rect -383 -249 -367 -215
rect -467 -265 -367 -249
rect -189 -215 -89 -177
rect -189 -249 -173 -215
rect -105 -249 -89 -215
rect -189 -265 -89 -249
rect 89 -215 189 -177
rect 89 -249 105 -215
rect 173 -249 189 -215
rect 89 -265 189 -249
rect 367 -215 467 -177
rect 367 -249 383 -215
rect 451 -249 467 -215
rect 367 -265 467 -249
<< polycont >>
rect -451 -249 -383 -215
rect -173 -249 -105 -215
rect 105 -249 173 -215
rect 383 -249 451 -215
<< locali >>
rect -513 227 -479 243
rect -513 -181 -479 -165
rect -355 227 -321 243
rect -355 -181 -321 -165
rect -235 227 -201 243
rect -235 -181 -201 -165
rect -77 227 -43 243
rect -77 -181 -43 -165
rect 43 227 77 243
rect 43 -181 77 -165
rect 201 227 235 243
rect 201 -181 235 -165
rect 321 227 355 243
rect 321 -181 355 -165
rect 479 227 513 243
rect 479 -181 513 -165
rect -467 -249 -451 -215
rect -383 -249 -367 -215
rect -189 -249 -173 -215
rect -105 -249 -89 -215
rect 89 -249 105 -215
rect 173 -249 189 -215
rect 367 -249 383 -215
rect 451 -249 467 -215
<< viali >>
rect -513 -165 -479 227
rect -355 -165 -321 227
rect -235 -165 -201 227
rect -77 -165 -43 227
rect 43 -165 77 227
rect 201 -165 235 227
rect 321 -165 355 227
rect 479 -165 513 227
rect -451 -249 -383 -215
rect -173 -249 -105 -215
rect 105 -249 173 -215
rect 383 -249 451 -215
<< metal1 >>
rect -519 227 -473 239
rect -519 -165 -513 227
rect -479 -165 -473 227
rect -519 -177 -473 -165
rect -361 227 -315 239
rect -361 -165 -355 227
rect -321 -165 -315 227
rect -361 -177 -315 -165
rect -241 227 -195 239
rect -241 -165 -235 227
rect -201 -165 -195 227
rect -241 -177 -195 -165
rect -83 227 -37 239
rect -83 -165 -77 227
rect -43 -165 -37 227
rect -83 -177 -37 -165
rect 37 227 83 239
rect 37 -165 43 227
rect 77 -165 83 227
rect 37 -177 83 -165
rect 195 227 241 239
rect 195 -165 201 227
rect 235 -165 241 227
rect 195 -177 241 -165
rect 315 227 361 239
rect 315 -165 321 227
rect 355 -165 361 227
rect 315 -177 361 -165
rect 473 227 519 239
rect 473 -165 479 227
rect 513 -165 519 227
rect 473 -177 519 -165
rect -463 -215 -371 -209
rect -463 -249 -451 -215
rect -383 -249 -371 -215
rect -463 -255 -371 -249
rect -185 -215 -93 -209
rect -185 -249 -173 -215
rect -105 -249 -93 -215
rect -185 -255 -93 -249
rect 93 -215 185 -209
rect 93 -249 105 -215
rect 173 -249 185 -215
rect 93 -255 185 -249
rect 371 -215 463 -209
rect 371 -249 383 -215
rect 451 -249 463 -215
rect 371 -255 463 -249
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.08 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
