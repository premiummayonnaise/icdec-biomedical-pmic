** sch_path: /foss/designs/icdec-biomedical-pmic/xschem/5t-ota/schematics/5t-ota.sch
.subckt 5t-ota VDD OUT IBIAS VN VP VSS
*.PININFO VP:I VN:I IBIAS:I VDD:B VSS:B OUT:O
XM1 net1 VP net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.75 W=8.5 nf=4 m=1
XM2 OUT VN net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.75 W=8.5 nf=4 m=1
XM3 net2 IBIAS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1.25 W=1.58 nf=1 m=1
XM4 OUT net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.25 W=4.85 nf=2 m=1
XM5 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.25 W=4.85 nf=2 m=1
XM6 IBIAS IBIAS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1.25 W=1.58 nf=1 m=1
.ends
