magic
tech sky130A
magscale 1 2
timestamp 1769436194
<< error_p >>
rect -8931 -1129 -8901 1061
rect -8865 -1063 -8835 995
rect 8835 -1063 8865 995
rect -8865 -1067 -8649 -1063
rect -8587 -1067 -8371 -1063
rect -8309 -1067 -8093 -1063
rect -8031 -1067 -7815 -1063
rect -7753 -1067 -7537 -1063
rect -7475 -1067 -7259 -1063
rect -7197 -1067 -6981 -1063
rect -6919 -1067 -6703 -1063
rect -6641 -1067 -6425 -1063
rect -6363 -1067 -6147 -1063
rect -6085 -1067 -5869 -1063
rect -5807 -1067 -5591 -1063
rect -5529 -1067 -5313 -1063
rect -5251 -1067 -5035 -1063
rect -4973 -1067 -4757 -1063
rect -4695 -1067 -4479 -1063
rect -4417 -1067 -4201 -1063
rect -4139 -1067 -3923 -1063
rect -3861 -1067 -3645 -1063
rect -3583 -1067 -3367 -1063
rect -3305 -1067 -3089 -1063
rect -3027 -1067 -2811 -1063
rect -2749 -1067 -2533 -1063
rect -2471 -1067 -2255 -1063
rect -2193 -1067 -1977 -1063
rect -1915 -1067 -1699 -1063
rect -1637 -1067 -1421 -1063
rect -1359 -1067 -1143 -1063
rect -1081 -1067 -865 -1063
rect -803 -1067 -587 -1063
rect -525 -1067 -309 -1063
rect -247 -1067 -31 -1063
rect 31 -1067 247 -1063
rect 309 -1067 525 -1063
rect 587 -1067 803 -1063
rect 865 -1067 1081 -1063
rect 1143 -1067 1359 -1063
rect 1421 -1067 1637 -1063
rect 1699 -1067 1915 -1063
rect 1977 -1067 2193 -1063
rect 2255 -1067 2471 -1063
rect 2533 -1067 2749 -1063
rect 2811 -1067 3027 -1063
rect 3089 -1067 3305 -1063
rect 3367 -1067 3583 -1063
rect 3645 -1067 3861 -1063
rect 3923 -1067 4139 -1063
rect 4201 -1067 4417 -1063
rect 4479 -1067 4695 -1063
rect 4757 -1067 4973 -1063
rect 5035 -1067 5251 -1063
rect 5313 -1067 5529 -1063
rect 5591 -1067 5807 -1063
rect 5869 -1067 6085 -1063
rect 6147 -1067 6363 -1063
rect 6425 -1067 6641 -1063
rect 6703 -1067 6919 -1063
rect 6981 -1067 7197 -1063
rect 7259 -1067 7475 -1063
rect 7537 -1067 7753 -1063
rect 7815 -1067 8031 -1063
rect 8093 -1067 8309 -1063
rect 8371 -1067 8587 -1063
rect 8649 -1067 8865 -1063
rect 8901 -1129 8931 1061
rect -8931 -1133 8931 -1129
<< nwell >>
rect -8901 -1129 8901 1095
<< mvpmos >>
rect -8807 -1067 -8707 995
rect -8529 -1067 -8429 995
rect -8251 -1067 -8151 995
rect -7973 -1067 -7873 995
rect -7695 -1067 -7595 995
rect -7417 -1067 -7317 995
rect -7139 -1067 -7039 995
rect -6861 -1067 -6761 995
rect -6583 -1067 -6483 995
rect -6305 -1067 -6205 995
rect -6027 -1067 -5927 995
rect -5749 -1067 -5649 995
rect -5471 -1067 -5371 995
rect -5193 -1067 -5093 995
rect -4915 -1067 -4815 995
rect -4637 -1067 -4537 995
rect -4359 -1067 -4259 995
rect -4081 -1067 -3981 995
rect -3803 -1067 -3703 995
rect -3525 -1067 -3425 995
rect -3247 -1067 -3147 995
rect -2969 -1067 -2869 995
rect -2691 -1067 -2591 995
rect -2413 -1067 -2313 995
rect -2135 -1067 -2035 995
rect -1857 -1067 -1757 995
rect -1579 -1067 -1479 995
rect -1301 -1067 -1201 995
rect -1023 -1067 -923 995
rect -745 -1067 -645 995
rect -467 -1067 -367 995
rect -189 -1067 -89 995
rect 89 -1067 189 995
rect 367 -1067 467 995
rect 645 -1067 745 995
rect 923 -1067 1023 995
rect 1201 -1067 1301 995
rect 1479 -1067 1579 995
rect 1757 -1067 1857 995
rect 2035 -1067 2135 995
rect 2313 -1067 2413 995
rect 2591 -1067 2691 995
rect 2869 -1067 2969 995
rect 3147 -1067 3247 995
rect 3425 -1067 3525 995
rect 3703 -1067 3803 995
rect 3981 -1067 4081 995
rect 4259 -1067 4359 995
rect 4537 -1067 4637 995
rect 4815 -1067 4915 995
rect 5093 -1067 5193 995
rect 5371 -1067 5471 995
rect 5649 -1067 5749 995
rect 5927 -1067 6027 995
rect 6205 -1067 6305 995
rect 6483 -1067 6583 995
rect 6761 -1067 6861 995
rect 7039 -1067 7139 995
rect 7317 -1067 7417 995
rect 7595 -1067 7695 995
rect 7873 -1067 7973 995
rect 8151 -1067 8251 995
rect 8429 -1067 8529 995
rect 8707 -1067 8807 995
<< mvpdiff >>
rect -8865 983 -8807 995
rect -8865 -1055 -8853 983
rect -8819 -1055 -8807 983
rect -8865 -1067 -8807 -1055
rect -8707 983 -8649 995
rect -8707 -1055 -8695 983
rect -8661 -1055 -8649 983
rect -8707 -1067 -8649 -1055
rect -8587 983 -8529 995
rect -8587 -1055 -8575 983
rect -8541 -1055 -8529 983
rect -8587 -1067 -8529 -1055
rect -8429 983 -8371 995
rect -8429 -1055 -8417 983
rect -8383 -1055 -8371 983
rect -8429 -1067 -8371 -1055
rect -8309 983 -8251 995
rect -8309 -1055 -8297 983
rect -8263 -1055 -8251 983
rect -8309 -1067 -8251 -1055
rect -8151 983 -8093 995
rect -8151 -1055 -8139 983
rect -8105 -1055 -8093 983
rect -8151 -1067 -8093 -1055
rect -8031 983 -7973 995
rect -8031 -1055 -8019 983
rect -7985 -1055 -7973 983
rect -8031 -1067 -7973 -1055
rect -7873 983 -7815 995
rect -7873 -1055 -7861 983
rect -7827 -1055 -7815 983
rect -7873 -1067 -7815 -1055
rect -7753 983 -7695 995
rect -7753 -1055 -7741 983
rect -7707 -1055 -7695 983
rect -7753 -1067 -7695 -1055
rect -7595 983 -7537 995
rect -7595 -1055 -7583 983
rect -7549 -1055 -7537 983
rect -7595 -1067 -7537 -1055
rect -7475 983 -7417 995
rect -7475 -1055 -7463 983
rect -7429 -1055 -7417 983
rect -7475 -1067 -7417 -1055
rect -7317 983 -7259 995
rect -7317 -1055 -7305 983
rect -7271 -1055 -7259 983
rect -7317 -1067 -7259 -1055
rect -7197 983 -7139 995
rect -7197 -1055 -7185 983
rect -7151 -1055 -7139 983
rect -7197 -1067 -7139 -1055
rect -7039 983 -6981 995
rect -7039 -1055 -7027 983
rect -6993 -1055 -6981 983
rect -7039 -1067 -6981 -1055
rect -6919 983 -6861 995
rect -6919 -1055 -6907 983
rect -6873 -1055 -6861 983
rect -6919 -1067 -6861 -1055
rect -6761 983 -6703 995
rect -6761 -1055 -6749 983
rect -6715 -1055 -6703 983
rect -6761 -1067 -6703 -1055
rect -6641 983 -6583 995
rect -6641 -1055 -6629 983
rect -6595 -1055 -6583 983
rect -6641 -1067 -6583 -1055
rect -6483 983 -6425 995
rect -6483 -1055 -6471 983
rect -6437 -1055 -6425 983
rect -6483 -1067 -6425 -1055
rect -6363 983 -6305 995
rect -6363 -1055 -6351 983
rect -6317 -1055 -6305 983
rect -6363 -1067 -6305 -1055
rect -6205 983 -6147 995
rect -6205 -1055 -6193 983
rect -6159 -1055 -6147 983
rect -6205 -1067 -6147 -1055
rect -6085 983 -6027 995
rect -6085 -1055 -6073 983
rect -6039 -1055 -6027 983
rect -6085 -1067 -6027 -1055
rect -5927 983 -5869 995
rect -5927 -1055 -5915 983
rect -5881 -1055 -5869 983
rect -5927 -1067 -5869 -1055
rect -5807 983 -5749 995
rect -5807 -1055 -5795 983
rect -5761 -1055 -5749 983
rect -5807 -1067 -5749 -1055
rect -5649 983 -5591 995
rect -5649 -1055 -5637 983
rect -5603 -1055 -5591 983
rect -5649 -1067 -5591 -1055
rect -5529 983 -5471 995
rect -5529 -1055 -5517 983
rect -5483 -1055 -5471 983
rect -5529 -1067 -5471 -1055
rect -5371 983 -5313 995
rect -5371 -1055 -5359 983
rect -5325 -1055 -5313 983
rect -5371 -1067 -5313 -1055
rect -5251 983 -5193 995
rect -5251 -1055 -5239 983
rect -5205 -1055 -5193 983
rect -5251 -1067 -5193 -1055
rect -5093 983 -5035 995
rect -5093 -1055 -5081 983
rect -5047 -1055 -5035 983
rect -5093 -1067 -5035 -1055
rect -4973 983 -4915 995
rect -4973 -1055 -4961 983
rect -4927 -1055 -4915 983
rect -4973 -1067 -4915 -1055
rect -4815 983 -4757 995
rect -4815 -1055 -4803 983
rect -4769 -1055 -4757 983
rect -4815 -1067 -4757 -1055
rect -4695 983 -4637 995
rect -4695 -1055 -4683 983
rect -4649 -1055 -4637 983
rect -4695 -1067 -4637 -1055
rect -4537 983 -4479 995
rect -4537 -1055 -4525 983
rect -4491 -1055 -4479 983
rect -4537 -1067 -4479 -1055
rect -4417 983 -4359 995
rect -4417 -1055 -4405 983
rect -4371 -1055 -4359 983
rect -4417 -1067 -4359 -1055
rect -4259 983 -4201 995
rect -4259 -1055 -4247 983
rect -4213 -1055 -4201 983
rect -4259 -1067 -4201 -1055
rect -4139 983 -4081 995
rect -4139 -1055 -4127 983
rect -4093 -1055 -4081 983
rect -4139 -1067 -4081 -1055
rect -3981 983 -3923 995
rect -3981 -1055 -3969 983
rect -3935 -1055 -3923 983
rect -3981 -1067 -3923 -1055
rect -3861 983 -3803 995
rect -3861 -1055 -3849 983
rect -3815 -1055 -3803 983
rect -3861 -1067 -3803 -1055
rect -3703 983 -3645 995
rect -3703 -1055 -3691 983
rect -3657 -1055 -3645 983
rect -3703 -1067 -3645 -1055
rect -3583 983 -3525 995
rect -3583 -1055 -3571 983
rect -3537 -1055 -3525 983
rect -3583 -1067 -3525 -1055
rect -3425 983 -3367 995
rect -3425 -1055 -3413 983
rect -3379 -1055 -3367 983
rect -3425 -1067 -3367 -1055
rect -3305 983 -3247 995
rect -3305 -1055 -3293 983
rect -3259 -1055 -3247 983
rect -3305 -1067 -3247 -1055
rect -3147 983 -3089 995
rect -3147 -1055 -3135 983
rect -3101 -1055 -3089 983
rect -3147 -1067 -3089 -1055
rect -3027 983 -2969 995
rect -3027 -1055 -3015 983
rect -2981 -1055 -2969 983
rect -3027 -1067 -2969 -1055
rect -2869 983 -2811 995
rect -2869 -1055 -2857 983
rect -2823 -1055 -2811 983
rect -2869 -1067 -2811 -1055
rect -2749 983 -2691 995
rect -2749 -1055 -2737 983
rect -2703 -1055 -2691 983
rect -2749 -1067 -2691 -1055
rect -2591 983 -2533 995
rect -2591 -1055 -2579 983
rect -2545 -1055 -2533 983
rect -2591 -1067 -2533 -1055
rect -2471 983 -2413 995
rect -2471 -1055 -2459 983
rect -2425 -1055 -2413 983
rect -2471 -1067 -2413 -1055
rect -2313 983 -2255 995
rect -2313 -1055 -2301 983
rect -2267 -1055 -2255 983
rect -2313 -1067 -2255 -1055
rect -2193 983 -2135 995
rect -2193 -1055 -2181 983
rect -2147 -1055 -2135 983
rect -2193 -1067 -2135 -1055
rect -2035 983 -1977 995
rect -2035 -1055 -2023 983
rect -1989 -1055 -1977 983
rect -2035 -1067 -1977 -1055
rect -1915 983 -1857 995
rect -1915 -1055 -1903 983
rect -1869 -1055 -1857 983
rect -1915 -1067 -1857 -1055
rect -1757 983 -1699 995
rect -1757 -1055 -1745 983
rect -1711 -1055 -1699 983
rect -1757 -1067 -1699 -1055
rect -1637 983 -1579 995
rect -1637 -1055 -1625 983
rect -1591 -1055 -1579 983
rect -1637 -1067 -1579 -1055
rect -1479 983 -1421 995
rect -1479 -1055 -1467 983
rect -1433 -1055 -1421 983
rect -1479 -1067 -1421 -1055
rect -1359 983 -1301 995
rect -1359 -1055 -1347 983
rect -1313 -1055 -1301 983
rect -1359 -1067 -1301 -1055
rect -1201 983 -1143 995
rect -1201 -1055 -1189 983
rect -1155 -1055 -1143 983
rect -1201 -1067 -1143 -1055
rect -1081 983 -1023 995
rect -1081 -1055 -1069 983
rect -1035 -1055 -1023 983
rect -1081 -1067 -1023 -1055
rect -923 983 -865 995
rect -923 -1055 -911 983
rect -877 -1055 -865 983
rect -923 -1067 -865 -1055
rect -803 983 -745 995
rect -803 -1055 -791 983
rect -757 -1055 -745 983
rect -803 -1067 -745 -1055
rect -645 983 -587 995
rect -645 -1055 -633 983
rect -599 -1055 -587 983
rect -645 -1067 -587 -1055
rect -525 983 -467 995
rect -525 -1055 -513 983
rect -479 -1055 -467 983
rect -525 -1067 -467 -1055
rect -367 983 -309 995
rect -367 -1055 -355 983
rect -321 -1055 -309 983
rect -367 -1067 -309 -1055
rect -247 983 -189 995
rect -247 -1055 -235 983
rect -201 -1055 -189 983
rect -247 -1067 -189 -1055
rect -89 983 -31 995
rect -89 -1055 -77 983
rect -43 -1055 -31 983
rect -89 -1067 -31 -1055
rect 31 983 89 995
rect 31 -1055 43 983
rect 77 -1055 89 983
rect 31 -1067 89 -1055
rect 189 983 247 995
rect 189 -1055 201 983
rect 235 -1055 247 983
rect 189 -1067 247 -1055
rect 309 983 367 995
rect 309 -1055 321 983
rect 355 -1055 367 983
rect 309 -1067 367 -1055
rect 467 983 525 995
rect 467 -1055 479 983
rect 513 -1055 525 983
rect 467 -1067 525 -1055
rect 587 983 645 995
rect 587 -1055 599 983
rect 633 -1055 645 983
rect 587 -1067 645 -1055
rect 745 983 803 995
rect 745 -1055 757 983
rect 791 -1055 803 983
rect 745 -1067 803 -1055
rect 865 983 923 995
rect 865 -1055 877 983
rect 911 -1055 923 983
rect 865 -1067 923 -1055
rect 1023 983 1081 995
rect 1023 -1055 1035 983
rect 1069 -1055 1081 983
rect 1023 -1067 1081 -1055
rect 1143 983 1201 995
rect 1143 -1055 1155 983
rect 1189 -1055 1201 983
rect 1143 -1067 1201 -1055
rect 1301 983 1359 995
rect 1301 -1055 1313 983
rect 1347 -1055 1359 983
rect 1301 -1067 1359 -1055
rect 1421 983 1479 995
rect 1421 -1055 1433 983
rect 1467 -1055 1479 983
rect 1421 -1067 1479 -1055
rect 1579 983 1637 995
rect 1579 -1055 1591 983
rect 1625 -1055 1637 983
rect 1579 -1067 1637 -1055
rect 1699 983 1757 995
rect 1699 -1055 1711 983
rect 1745 -1055 1757 983
rect 1699 -1067 1757 -1055
rect 1857 983 1915 995
rect 1857 -1055 1869 983
rect 1903 -1055 1915 983
rect 1857 -1067 1915 -1055
rect 1977 983 2035 995
rect 1977 -1055 1989 983
rect 2023 -1055 2035 983
rect 1977 -1067 2035 -1055
rect 2135 983 2193 995
rect 2135 -1055 2147 983
rect 2181 -1055 2193 983
rect 2135 -1067 2193 -1055
rect 2255 983 2313 995
rect 2255 -1055 2267 983
rect 2301 -1055 2313 983
rect 2255 -1067 2313 -1055
rect 2413 983 2471 995
rect 2413 -1055 2425 983
rect 2459 -1055 2471 983
rect 2413 -1067 2471 -1055
rect 2533 983 2591 995
rect 2533 -1055 2545 983
rect 2579 -1055 2591 983
rect 2533 -1067 2591 -1055
rect 2691 983 2749 995
rect 2691 -1055 2703 983
rect 2737 -1055 2749 983
rect 2691 -1067 2749 -1055
rect 2811 983 2869 995
rect 2811 -1055 2823 983
rect 2857 -1055 2869 983
rect 2811 -1067 2869 -1055
rect 2969 983 3027 995
rect 2969 -1055 2981 983
rect 3015 -1055 3027 983
rect 2969 -1067 3027 -1055
rect 3089 983 3147 995
rect 3089 -1055 3101 983
rect 3135 -1055 3147 983
rect 3089 -1067 3147 -1055
rect 3247 983 3305 995
rect 3247 -1055 3259 983
rect 3293 -1055 3305 983
rect 3247 -1067 3305 -1055
rect 3367 983 3425 995
rect 3367 -1055 3379 983
rect 3413 -1055 3425 983
rect 3367 -1067 3425 -1055
rect 3525 983 3583 995
rect 3525 -1055 3537 983
rect 3571 -1055 3583 983
rect 3525 -1067 3583 -1055
rect 3645 983 3703 995
rect 3645 -1055 3657 983
rect 3691 -1055 3703 983
rect 3645 -1067 3703 -1055
rect 3803 983 3861 995
rect 3803 -1055 3815 983
rect 3849 -1055 3861 983
rect 3803 -1067 3861 -1055
rect 3923 983 3981 995
rect 3923 -1055 3935 983
rect 3969 -1055 3981 983
rect 3923 -1067 3981 -1055
rect 4081 983 4139 995
rect 4081 -1055 4093 983
rect 4127 -1055 4139 983
rect 4081 -1067 4139 -1055
rect 4201 983 4259 995
rect 4201 -1055 4213 983
rect 4247 -1055 4259 983
rect 4201 -1067 4259 -1055
rect 4359 983 4417 995
rect 4359 -1055 4371 983
rect 4405 -1055 4417 983
rect 4359 -1067 4417 -1055
rect 4479 983 4537 995
rect 4479 -1055 4491 983
rect 4525 -1055 4537 983
rect 4479 -1067 4537 -1055
rect 4637 983 4695 995
rect 4637 -1055 4649 983
rect 4683 -1055 4695 983
rect 4637 -1067 4695 -1055
rect 4757 983 4815 995
rect 4757 -1055 4769 983
rect 4803 -1055 4815 983
rect 4757 -1067 4815 -1055
rect 4915 983 4973 995
rect 4915 -1055 4927 983
rect 4961 -1055 4973 983
rect 4915 -1067 4973 -1055
rect 5035 983 5093 995
rect 5035 -1055 5047 983
rect 5081 -1055 5093 983
rect 5035 -1067 5093 -1055
rect 5193 983 5251 995
rect 5193 -1055 5205 983
rect 5239 -1055 5251 983
rect 5193 -1067 5251 -1055
rect 5313 983 5371 995
rect 5313 -1055 5325 983
rect 5359 -1055 5371 983
rect 5313 -1067 5371 -1055
rect 5471 983 5529 995
rect 5471 -1055 5483 983
rect 5517 -1055 5529 983
rect 5471 -1067 5529 -1055
rect 5591 983 5649 995
rect 5591 -1055 5603 983
rect 5637 -1055 5649 983
rect 5591 -1067 5649 -1055
rect 5749 983 5807 995
rect 5749 -1055 5761 983
rect 5795 -1055 5807 983
rect 5749 -1067 5807 -1055
rect 5869 983 5927 995
rect 5869 -1055 5881 983
rect 5915 -1055 5927 983
rect 5869 -1067 5927 -1055
rect 6027 983 6085 995
rect 6027 -1055 6039 983
rect 6073 -1055 6085 983
rect 6027 -1067 6085 -1055
rect 6147 983 6205 995
rect 6147 -1055 6159 983
rect 6193 -1055 6205 983
rect 6147 -1067 6205 -1055
rect 6305 983 6363 995
rect 6305 -1055 6317 983
rect 6351 -1055 6363 983
rect 6305 -1067 6363 -1055
rect 6425 983 6483 995
rect 6425 -1055 6437 983
rect 6471 -1055 6483 983
rect 6425 -1067 6483 -1055
rect 6583 983 6641 995
rect 6583 -1055 6595 983
rect 6629 -1055 6641 983
rect 6583 -1067 6641 -1055
rect 6703 983 6761 995
rect 6703 -1055 6715 983
rect 6749 -1055 6761 983
rect 6703 -1067 6761 -1055
rect 6861 983 6919 995
rect 6861 -1055 6873 983
rect 6907 -1055 6919 983
rect 6861 -1067 6919 -1055
rect 6981 983 7039 995
rect 6981 -1055 6993 983
rect 7027 -1055 7039 983
rect 6981 -1067 7039 -1055
rect 7139 983 7197 995
rect 7139 -1055 7151 983
rect 7185 -1055 7197 983
rect 7139 -1067 7197 -1055
rect 7259 983 7317 995
rect 7259 -1055 7271 983
rect 7305 -1055 7317 983
rect 7259 -1067 7317 -1055
rect 7417 983 7475 995
rect 7417 -1055 7429 983
rect 7463 -1055 7475 983
rect 7417 -1067 7475 -1055
rect 7537 983 7595 995
rect 7537 -1055 7549 983
rect 7583 -1055 7595 983
rect 7537 -1067 7595 -1055
rect 7695 983 7753 995
rect 7695 -1055 7707 983
rect 7741 -1055 7753 983
rect 7695 -1067 7753 -1055
rect 7815 983 7873 995
rect 7815 -1055 7827 983
rect 7861 -1055 7873 983
rect 7815 -1067 7873 -1055
rect 7973 983 8031 995
rect 7973 -1055 7985 983
rect 8019 -1055 8031 983
rect 7973 -1067 8031 -1055
rect 8093 983 8151 995
rect 8093 -1055 8105 983
rect 8139 -1055 8151 983
rect 8093 -1067 8151 -1055
rect 8251 983 8309 995
rect 8251 -1055 8263 983
rect 8297 -1055 8309 983
rect 8251 -1067 8309 -1055
rect 8371 983 8429 995
rect 8371 -1055 8383 983
rect 8417 -1055 8429 983
rect 8371 -1067 8429 -1055
rect 8529 983 8587 995
rect 8529 -1055 8541 983
rect 8575 -1055 8587 983
rect 8529 -1067 8587 -1055
rect 8649 983 8707 995
rect 8649 -1055 8661 983
rect 8695 -1055 8707 983
rect 8649 -1067 8707 -1055
rect 8807 983 8865 995
rect 8807 -1055 8819 983
rect 8853 -1055 8865 983
rect 8807 -1067 8865 -1055
<< mvpdiffc >>
rect -8853 -1055 -8819 983
rect -8695 -1055 -8661 983
rect -8575 -1055 -8541 983
rect -8417 -1055 -8383 983
rect -8297 -1055 -8263 983
rect -8139 -1055 -8105 983
rect -8019 -1055 -7985 983
rect -7861 -1055 -7827 983
rect -7741 -1055 -7707 983
rect -7583 -1055 -7549 983
rect -7463 -1055 -7429 983
rect -7305 -1055 -7271 983
rect -7185 -1055 -7151 983
rect -7027 -1055 -6993 983
rect -6907 -1055 -6873 983
rect -6749 -1055 -6715 983
rect -6629 -1055 -6595 983
rect -6471 -1055 -6437 983
rect -6351 -1055 -6317 983
rect -6193 -1055 -6159 983
rect -6073 -1055 -6039 983
rect -5915 -1055 -5881 983
rect -5795 -1055 -5761 983
rect -5637 -1055 -5603 983
rect -5517 -1055 -5483 983
rect -5359 -1055 -5325 983
rect -5239 -1055 -5205 983
rect -5081 -1055 -5047 983
rect -4961 -1055 -4927 983
rect -4803 -1055 -4769 983
rect -4683 -1055 -4649 983
rect -4525 -1055 -4491 983
rect -4405 -1055 -4371 983
rect -4247 -1055 -4213 983
rect -4127 -1055 -4093 983
rect -3969 -1055 -3935 983
rect -3849 -1055 -3815 983
rect -3691 -1055 -3657 983
rect -3571 -1055 -3537 983
rect -3413 -1055 -3379 983
rect -3293 -1055 -3259 983
rect -3135 -1055 -3101 983
rect -3015 -1055 -2981 983
rect -2857 -1055 -2823 983
rect -2737 -1055 -2703 983
rect -2579 -1055 -2545 983
rect -2459 -1055 -2425 983
rect -2301 -1055 -2267 983
rect -2181 -1055 -2147 983
rect -2023 -1055 -1989 983
rect -1903 -1055 -1869 983
rect -1745 -1055 -1711 983
rect -1625 -1055 -1591 983
rect -1467 -1055 -1433 983
rect -1347 -1055 -1313 983
rect -1189 -1055 -1155 983
rect -1069 -1055 -1035 983
rect -911 -1055 -877 983
rect -791 -1055 -757 983
rect -633 -1055 -599 983
rect -513 -1055 -479 983
rect -355 -1055 -321 983
rect -235 -1055 -201 983
rect -77 -1055 -43 983
rect 43 -1055 77 983
rect 201 -1055 235 983
rect 321 -1055 355 983
rect 479 -1055 513 983
rect 599 -1055 633 983
rect 757 -1055 791 983
rect 877 -1055 911 983
rect 1035 -1055 1069 983
rect 1155 -1055 1189 983
rect 1313 -1055 1347 983
rect 1433 -1055 1467 983
rect 1591 -1055 1625 983
rect 1711 -1055 1745 983
rect 1869 -1055 1903 983
rect 1989 -1055 2023 983
rect 2147 -1055 2181 983
rect 2267 -1055 2301 983
rect 2425 -1055 2459 983
rect 2545 -1055 2579 983
rect 2703 -1055 2737 983
rect 2823 -1055 2857 983
rect 2981 -1055 3015 983
rect 3101 -1055 3135 983
rect 3259 -1055 3293 983
rect 3379 -1055 3413 983
rect 3537 -1055 3571 983
rect 3657 -1055 3691 983
rect 3815 -1055 3849 983
rect 3935 -1055 3969 983
rect 4093 -1055 4127 983
rect 4213 -1055 4247 983
rect 4371 -1055 4405 983
rect 4491 -1055 4525 983
rect 4649 -1055 4683 983
rect 4769 -1055 4803 983
rect 4927 -1055 4961 983
rect 5047 -1055 5081 983
rect 5205 -1055 5239 983
rect 5325 -1055 5359 983
rect 5483 -1055 5517 983
rect 5603 -1055 5637 983
rect 5761 -1055 5795 983
rect 5881 -1055 5915 983
rect 6039 -1055 6073 983
rect 6159 -1055 6193 983
rect 6317 -1055 6351 983
rect 6437 -1055 6471 983
rect 6595 -1055 6629 983
rect 6715 -1055 6749 983
rect 6873 -1055 6907 983
rect 6993 -1055 7027 983
rect 7151 -1055 7185 983
rect 7271 -1055 7305 983
rect 7429 -1055 7463 983
rect 7549 -1055 7583 983
rect 7707 -1055 7741 983
rect 7827 -1055 7861 983
rect 7985 -1055 8019 983
rect 8105 -1055 8139 983
rect 8263 -1055 8297 983
rect 8383 -1055 8417 983
rect 8541 -1055 8575 983
rect 8661 -1055 8695 983
rect 8819 -1055 8853 983
<< poly >>
rect -8807 1076 -8707 1092
rect -8807 1042 -8791 1076
rect -8723 1042 -8707 1076
rect -8807 995 -8707 1042
rect -8529 1076 -8429 1092
rect -8529 1042 -8513 1076
rect -8445 1042 -8429 1076
rect -8529 995 -8429 1042
rect -8251 1076 -8151 1092
rect -8251 1042 -8235 1076
rect -8167 1042 -8151 1076
rect -8251 995 -8151 1042
rect -7973 1076 -7873 1092
rect -7973 1042 -7957 1076
rect -7889 1042 -7873 1076
rect -7973 995 -7873 1042
rect -7695 1076 -7595 1092
rect -7695 1042 -7679 1076
rect -7611 1042 -7595 1076
rect -7695 995 -7595 1042
rect -7417 1076 -7317 1092
rect -7417 1042 -7401 1076
rect -7333 1042 -7317 1076
rect -7417 995 -7317 1042
rect -7139 1076 -7039 1092
rect -7139 1042 -7123 1076
rect -7055 1042 -7039 1076
rect -7139 995 -7039 1042
rect -6861 1076 -6761 1092
rect -6861 1042 -6845 1076
rect -6777 1042 -6761 1076
rect -6861 995 -6761 1042
rect -6583 1076 -6483 1092
rect -6583 1042 -6567 1076
rect -6499 1042 -6483 1076
rect -6583 995 -6483 1042
rect -6305 1076 -6205 1092
rect -6305 1042 -6289 1076
rect -6221 1042 -6205 1076
rect -6305 995 -6205 1042
rect -6027 1076 -5927 1092
rect -6027 1042 -6011 1076
rect -5943 1042 -5927 1076
rect -6027 995 -5927 1042
rect -5749 1076 -5649 1092
rect -5749 1042 -5733 1076
rect -5665 1042 -5649 1076
rect -5749 995 -5649 1042
rect -5471 1076 -5371 1092
rect -5471 1042 -5455 1076
rect -5387 1042 -5371 1076
rect -5471 995 -5371 1042
rect -5193 1076 -5093 1092
rect -5193 1042 -5177 1076
rect -5109 1042 -5093 1076
rect -5193 995 -5093 1042
rect -4915 1076 -4815 1092
rect -4915 1042 -4899 1076
rect -4831 1042 -4815 1076
rect -4915 995 -4815 1042
rect -4637 1076 -4537 1092
rect -4637 1042 -4621 1076
rect -4553 1042 -4537 1076
rect -4637 995 -4537 1042
rect -4359 1076 -4259 1092
rect -4359 1042 -4343 1076
rect -4275 1042 -4259 1076
rect -4359 995 -4259 1042
rect -4081 1076 -3981 1092
rect -4081 1042 -4065 1076
rect -3997 1042 -3981 1076
rect -4081 995 -3981 1042
rect -3803 1076 -3703 1092
rect -3803 1042 -3787 1076
rect -3719 1042 -3703 1076
rect -3803 995 -3703 1042
rect -3525 1076 -3425 1092
rect -3525 1042 -3509 1076
rect -3441 1042 -3425 1076
rect -3525 995 -3425 1042
rect -3247 1076 -3147 1092
rect -3247 1042 -3231 1076
rect -3163 1042 -3147 1076
rect -3247 995 -3147 1042
rect -2969 1076 -2869 1092
rect -2969 1042 -2953 1076
rect -2885 1042 -2869 1076
rect -2969 995 -2869 1042
rect -2691 1076 -2591 1092
rect -2691 1042 -2675 1076
rect -2607 1042 -2591 1076
rect -2691 995 -2591 1042
rect -2413 1076 -2313 1092
rect -2413 1042 -2397 1076
rect -2329 1042 -2313 1076
rect -2413 995 -2313 1042
rect -2135 1076 -2035 1092
rect -2135 1042 -2119 1076
rect -2051 1042 -2035 1076
rect -2135 995 -2035 1042
rect -1857 1076 -1757 1092
rect -1857 1042 -1841 1076
rect -1773 1042 -1757 1076
rect -1857 995 -1757 1042
rect -1579 1076 -1479 1092
rect -1579 1042 -1563 1076
rect -1495 1042 -1479 1076
rect -1579 995 -1479 1042
rect -1301 1076 -1201 1092
rect -1301 1042 -1285 1076
rect -1217 1042 -1201 1076
rect -1301 995 -1201 1042
rect -1023 1076 -923 1092
rect -1023 1042 -1007 1076
rect -939 1042 -923 1076
rect -1023 995 -923 1042
rect -745 1076 -645 1092
rect -745 1042 -729 1076
rect -661 1042 -645 1076
rect -745 995 -645 1042
rect -467 1076 -367 1092
rect -467 1042 -451 1076
rect -383 1042 -367 1076
rect -467 995 -367 1042
rect -189 1076 -89 1092
rect -189 1042 -173 1076
rect -105 1042 -89 1076
rect -189 995 -89 1042
rect 89 1076 189 1092
rect 89 1042 105 1076
rect 173 1042 189 1076
rect 89 995 189 1042
rect 367 1076 467 1092
rect 367 1042 383 1076
rect 451 1042 467 1076
rect 367 995 467 1042
rect 645 1076 745 1092
rect 645 1042 661 1076
rect 729 1042 745 1076
rect 645 995 745 1042
rect 923 1076 1023 1092
rect 923 1042 939 1076
rect 1007 1042 1023 1076
rect 923 995 1023 1042
rect 1201 1076 1301 1092
rect 1201 1042 1217 1076
rect 1285 1042 1301 1076
rect 1201 995 1301 1042
rect 1479 1076 1579 1092
rect 1479 1042 1495 1076
rect 1563 1042 1579 1076
rect 1479 995 1579 1042
rect 1757 1076 1857 1092
rect 1757 1042 1773 1076
rect 1841 1042 1857 1076
rect 1757 995 1857 1042
rect 2035 1076 2135 1092
rect 2035 1042 2051 1076
rect 2119 1042 2135 1076
rect 2035 995 2135 1042
rect 2313 1076 2413 1092
rect 2313 1042 2329 1076
rect 2397 1042 2413 1076
rect 2313 995 2413 1042
rect 2591 1076 2691 1092
rect 2591 1042 2607 1076
rect 2675 1042 2691 1076
rect 2591 995 2691 1042
rect 2869 1076 2969 1092
rect 2869 1042 2885 1076
rect 2953 1042 2969 1076
rect 2869 995 2969 1042
rect 3147 1076 3247 1092
rect 3147 1042 3163 1076
rect 3231 1042 3247 1076
rect 3147 995 3247 1042
rect 3425 1076 3525 1092
rect 3425 1042 3441 1076
rect 3509 1042 3525 1076
rect 3425 995 3525 1042
rect 3703 1076 3803 1092
rect 3703 1042 3719 1076
rect 3787 1042 3803 1076
rect 3703 995 3803 1042
rect 3981 1076 4081 1092
rect 3981 1042 3997 1076
rect 4065 1042 4081 1076
rect 3981 995 4081 1042
rect 4259 1076 4359 1092
rect 4259 1042 4275 1076
rect 4343 1042 4359 1076
rect 4259 995 4359 1042
rect 4537 1076 4637 1092
rect 4537 1042 4553 1076
rect 4621 1042 4637 1076
rect 4537 995 4637 1042
rect 4815 1076 4915 1092
rect 4815 1042 4831 1076
rect 4899 1042 4915 1076
rect 4815 995 4915 1042
rect 5093 1076 5193 1092
rect 5093 1042 5109 1076
rect 5177 1042 5193 1076
rect 5093 995 5193 1042
rect 5371 1076 5471 1092
rect 5371 1042 5387 1076
rect 5455 1042 5471 1076
rect 5371 995 5471 1042
rect 5649 1076 5749 1092
rect 5649 1042 5665 1076
rect 5733 1042 5749 1076
rect 5649 995 5749 1042
rect 5927 1076 6027 1092
rect 5927 1042 5943 1076
rect 6011 1042 6027 1076
rect 5927 995 6027 1042
rect 6205 1076 6305 1092
rect 6205 1042 6221 1076
rect 6289 1042 6305 1076
rect 6205 995 6305 1042
rect 6483 1076 6583 1092
rect 6483 1042 6499 1076
rect 6567 1042 6583 1076
rect 6483 995 6583 1042
rect 6761 1076 6861 1092
rect 6761 1042 6777 1076
rect 6845 1042 6861 1076
rect 6761 995 6861 1042
rect 7039 1076 7139 1092
rect 7039 1042 7055 1076
rect 7123 1042 7139 1076
rect 7039 995 7139 1042
rect 7317 1076 7417 1092
rect 7317 1042 7333 1076
rect 7401 1042 7417 1076
rect 7317 995 7417 1042
rect 7595 1076 7695 1092
rect 7595 1042 7611 1076
rect 7679 1042 7695 1076
rect 7595 995 7695 1042
rect 7873 1076 7973 1092
rect 7873 1042 7889 1076
rect 7957 1042 7973 1076
rect 7873 995 7973 1042
rect 8151 1076 8251 1092
rect 8151 1042 8167 1076
rect 8235 1042 8251 1076
rect 8151 995 8251 1042
rect 8429 1076 8529 1092
rect 8429 1042 8445 1076
rect 8513 1042 8529 1076
rect 8429 995 8529 1042
rect 8707 1076 8807 1092
rect 8707 1042 8723 1076
rect 8791 1042 8807 1076
rect 8707 995 8807 1042
rect -8807 -1093 -8707 -1067
rect -8529 -1093 -8429 -1067
rect -8251 -1093 -8151 -1067
rect -7973 -1093 -7873 -1067
rect -7695 -1093 -7595 -1067
rect -7417 -1093 -7317 -1067
rect -7139 -1093 -7039 -1067
rect -6861 -1093 -6761 -1067
rect -6583 -1093 -6483 -1067
rect -6305 -1093 -6205 -1067
rect -6027 -1093 -5927 -1067
rect -5749 -1093 -5649 -1067
rect -5471 -1093 -5371 -1067
rect -5193 -1093 -5093 -1067
rect -4915 -1093 -4815 -1067
rect -4637 -1093 -4537 -1067
rect -4359 -1093 -4259 -1067
rect -4081 -1093 -3981 -1067
rect -3803 -1093 -3703 -1067
rect -3525 -1093 -3425 -1067
rect -3247 -1093 -3147 -1067
rect -2969 -1093 -2869 -1067
rect -2691 -1093 -2591 -1067
rect -2413 -1093 -2313 -1067
rect -2135 -1093 -2035 -1067
rect -1857 -1093 -1757 -1067
rect -1579 -1093 -1479 -1067
rect -1301 -1093 -1201 -1067
rect -1023 -1093 -923 -1067
rect -745 -1093 -645 -1067
rect -467 -1093 -367 -1067
rect -189 -1093 -89 -1067
rect 89 -1093 189 -1067
rect 367 -1093 467 -1067
rect 645 -1093 745 -1067
rect 923 -1093 1023 -1067
rect 1201 -1093 1301 -1067
rect 1479 -1093 1579 -1067
rect 1757 -1093 1857 -1067
rect 2035 -1093 2135 -1067
rect 2313 -1093 2413 -1067
rect 2591 -1093 2691 -1067
rect 2869 -1093 2969 -1067
rect 3147 -1093 3247 -1067
rect 3425 -1093 3525 -1067
rect 3703 -1093 3803 -1067
rect 3981 -1093 4081 -1067
rect 4259 -1093 4359 -1067
rect 4537 -1093 4637 -1067
rect 4815 -1093 4915 -1067
rect 5093 -1093 5193 -1067
rect 5371 -1093 5471 -1067
rect 5649 -1093 5749 -1067
rect 5927 -1093 6027 -1067
rect 6205 -1093 6305 -1067
rect 6483 -1093 6583 -1067
rect 6761 -1093 6861 -1067
rect 7039 -1093 7139 -1067
rect 7317 -1093 7417 -1067
rect 7595 -1093 7695 -1067
rect 7873 -1093 7973 -1067
rect 8151 -1093 8251 -1067
rect 8429 -1093 8529 -1067
rect 8707 -1093 8807 -1067
<< polycont >>
rect -8791 1042 -8723 1076
rect -8513 1042 -8445 1076
rect -8235 1042 -8167 1076
rect -7957 1042 -7889 1076
rect -7679 1042 -7611 1076
rect -7401 1042 -7333 1076
rect -7123 1042 -7055 1076
rect -6845 1042 -6777 1076
rect -6567 1042 -6499 1076
rect -6289 1042 -6221 1076
rect -6011 1042 -5943 1076
rect -5733 1042 -5665 1076
rect -5455 1042 -5387 1076
rect -5177 1042 -5109 1076
rect -4899 1042 -4831 1076
rect -4621 1042 -4553 1076
rect -4343 1042 -4275 1076
rect -4065 1042 -3997 1076
rect -3787 1042 -3719 1076
rect -3509 1042 -3441 1076
rect -3231 1042 -3163 1076
rect -2953 1042 -2885 1076
rect -2675 1042 -2607 1076
rect -2397 1042 -2329 1076
rect -2119 1042 -2051 1076
rect -1841 1042 -1773 1076
rect -1563 1042 -1495 1076
rect -1285 1042 -1217 1076
rect -1007 1042 -939 1076
rect -729 1042 -661 1076
rect -451 1042 -383 1076
rect -173 1042 -105 1076
rect 105 1042 173 1076
rect 383 1042 451 1076
rect 661 1042 729 1076
rect 939 1042 1007 1076
rect 1217 1042 1285 1076
rect 1495 1042 1563 1076
rect 1773 1042 1841 1076
rect 2051 1042 2119 1076
rect 2329 1042 2397 1076
rect 2607 1042 2675 1076
rect 2885 1042 2953 1076
rect 3163 1042 3231 1076
rect 3441 1042 3509 1076
rect 3719 1042 3787 1076
rect 3997 1042 4065 1076
rect 4275 1042 4343 1076
rect 4553 1042 4621 1076
rect 4831 1042 4899 1076
rect 5109 1042 5177 1076
rect 5387 1042 5455 1076
rect 5665 1042 5733 1076
rect 5943 1042 6011 1076
rect 6221 1042 6289 1076
rect 6499 1042 6567 1076
rect 6777 1042 6845 1076
rect 7055 1042 7123 1076
rect 7333 1042 7401 1076
rect 7611 1042 7679 1076
rect 7889 1042 7957 1076
rect 8167 1042 8235 1076
rect 8445 1042 8513 1076
rect 8723 1042 8791 1076
<< locali >>
rect -8807 1042 -8791 1076
rect -8723 1042 -8707 1076
rect -8529 1042 -8513 1076
rect -8445 1042 -8429 1076
rect -8251 1042 -8235 1076
rect -8167 1042 -8151 1076
rect -7973 1042 -7957 1076
rect -7889 1042 -7873 1076
rect -7695 1042 -7679 1076
rect -7611 1042 -7595 1076
rect -7417 1042 -7401 1076
rect -7333 1042 -7317 1076
rect -7139 1042 -7123 1076
rect -7055 1042 -7039 1076
rect -6861 1042 -6845 1076
rect -6777 1042 -6761 1076
rect -6583 1042 -6567 1076
rect -6499 1042 -6483 1076
rect -6305 1042 -6289 1076
rect -6221 1042 -6205 1076
rect -6027 1042 -6011 1076
rect -5943 1042 -5927 1076
rect -5749 1042 -5733 1076
rect -5665 1042 -5649 1076
rect -5471 1042 -5455 1076
rect -5387 1042 -5371 1076
rect -5193 1042 -5177 1076
rect -5109 1042 -5093 1076
rect -4915 1042 -4899 1076
rect -4831 1042 -4815 1076
rect -4637 1042 -4621 1076
rect -4553 1042 -4537 1076
rect -4359 1042 -4343 1076
rect -4275 1042 -4259 1076
rect -4081 1042 -4065 1076
rect -3997 1042 -3981 1076
rect -3803 1042 -3787 1076
rect -3719 1042 -3703 1076
rect -3525 1042 -3509 1076
rect -3441 1042 -3425 1076
rect -3247 1042 -3231 1076
rect -3163 1042 -3147 1076
rect -2969 1042 -2953 1076
rect -2885 1042 -2869 1076
rect -2691 1042 -2675 1076
rect -2607 1042 -2591 1076
rect -2413 1042 -2397 1076
rect -2329 1042 -2313 1076
rect -2135 1042 -2119 1076
rect -2051 1042 -2035 1076
rect -1857 1042 -1841 1076
rect -1773 1042 -1757 1076
rect -1579 1042 -1563 1076
rect -1495 1042 -1479 1076
rect -1301 1042 -1285 1076
rect -1217 1042 -1201 1076
rect -1023 1042 -1007 1076
rect -939 1042 -923 1076
rect -745 1042 -729 1076
rect -661 1042 -645 1076
rect -467 1042 -451 1076
rect -383 1042 -367 1076
rect -189 1042 -173 1076
rect -105 1042 -89 1076
rect 89 1042 105 1076
rect 173 1042 189 1076
rect 367 1042 383 1076
rect 451 1042 467 1076
rect 645 1042 661 1076
rect 729 1042 745 1076
rect 923 1042 939 1076
rect 1007 1042 1023 1076
rect 1201 1042 1217 1076
rect 1285 1042 1301 1076
rect 1479 1042 1495 1076
rect 1563 1042 1579 1076
rect 1757 1042 1773 1076
rect 1841 1042 1857 1076
rect 2035 1042 2051 1076
rect 2119 1042 2135 1076
rect 2313 1042 2329 1076
rect 2397 1042 2413 1076
rect 2591 1042 2607 1076
rect 2675 1042 2691 1076
rect 2869 1042 2885 1076
rect 2953 1042 2969 1076
rect 3147 1042 3163 1076
rect 3231 1042 3247 1076
rect 3425 1042 3441 1076
rect 3509 1042 3525 1076
rect 3703 1042 3719 1076
rect 3787 1042 3803 1076
rect 3981 1042 3997 1076
rect 4065 1042 4081 1076
rect 4259 1042 4275 1076
rect 4343 1042 4359 1076
rect 4537 1042 4553 1076
rect 4621 1042 4637 1076
rect 4815 1042 4831 1076
rect 4899 1042 4915 1076
rect 5093 1042 5109 1076
rect 5177 1042 5193 1076
rect 5371 1042 5387 1076
rect 5455 1042 5471 1076
rect 5649 1042 5665 1076
rect 5733 1042 5749 1076
rect 5927 1042 5943 1076
rect 6011 1042 6027 1076
rect 6205 1042 6221 1076
rect 6289 1042 6305 1076
rect 6483 1042 6499 1076
rect 6567 1042 6583 1076
rect 6761 1042 6777 1076
rect 6845 1042 6861 1076
rect 7039 1042 7055 1076
rect 7123 1042 7139 1076
rect 7317 1042 7333 1076
rect 7401 1042 7417 1076
rect 7595 1042 7611 1076
rect 7679 1042 7695 1076
rect 7873 1042 7889 1076
rect 7957 1042 7973 1076
rect 8151 1042 8167 1076
rect 8235 1042 8251 1076
rect 8429 1042 8445 1076
rect 8513 1042 8529 1076
rect 8707 1042 8723 1076
rect 8791 1042 8807 1076
rect -8853 983 -8819 999
rect -8853 -1071 -8819 -1055
rect -8695 983 -8661 999
rect -8695 -1071 -8661 -1055
rect -8575 983 -8541 999
rect -8575 -1071 -8541 -1055
rect -8417 983 -8383 999
rect -8417 -1071 -8383 -1055
rect -8297 983 -8263 999
rect -8297 -1071 -8263 -1055
rect -8139 983 -8105 999
rect -8139 -1071 -8105 -1055
rect -8019 983 -7985 999
rect -8019 -1071 -7985 -1055
rect -7861 983 -7827 999
rect -7861 -1071 -7827 -1055
rect -7741 983 -7707 999
rect -7741 -1071 -7707 -1055
rect -7583 983 -7549 999
rect -7583 -1071 -7549 -1055
rect -7463 983 -7429 999
rect -7463 -1071 -7429 -1055
rect -7305 983 -7271 999
rect -7305 -1071 -7271 -1055
rect -7185 983 -7151 999
rect -7185 -1071 -7151 -1055
rect -7027 983 -6993 999
rect -7027 -1071 -6993 -1055
rect -6907 983 -6873 999
rect -6907 -1071 -6873 -1055
rect -6749 983 -6715 999
rect -6749 -1071 -6715 -1055
rect -6629 983 -6595 999
rect -6629 -1071 -6595 -1055
rect -6471 983 -6437 999
rect -6471 -1071 -6437 -1055
rect -6351 983 -6317 999
rect -6351 -1071 -6317 -1055
rect -6193 983 -6159 999
rect -6193 -1071 -6159 -1055
rect -6073 983 -6039 999
rect -6073 -1071 -6039 -1055
rect -5915 983 -5881 999
rect -5915 -1071 -5881 -1055
rect -5795 983 -5761 999
rect -5795 -1071 -5761 -1055
rect -5637 983 -5603 999
rect -5637 -1071 -5603 -1055
rect -5517 983 -5483 999
rect -5517 -1071 -5483 -1055
rect -5359 983 -5325 999
rect -5359 -1071 -5325 -1055
rect -5239 983 -5205 999
rect -5239 -1071 -5205 -1055
rect -5081 983 -5047 999
rect -5081 -1071 -5047 -1055
rect -4961 983 -4927 999
rect -4961 -1071 -4927 -1055
rect -4803 983 -4769 999
rect -4803 -1071 -4769 -1055
rect -4683 983 -4649 999
rect -4683 -1071 -4649 -1055
rect -4525 983 -4491 999
rect -4525 -1071 -4491 -1055
rect -4405 983 -4371 999
rect -4405 -1071 -4371 -1055
rect -4247 983 -4213 999
rect -4247 -1071 -4213 -1055
rect -4127 983 -4093 999
rect -4127 -1071 -4093 -1055
rect -3969 983 -3935 999
rect -3969 -1071 -3935 -1055
rect -3849 983 -3815 999
rect -3849 -1071 -3815 -1055
rect -3691 983 -3657 999
rect -3691 -1071 -3657 -1055
rect -3571 983 -3537 999
rect -3571 -1071 -3537 -1055
rect -3413 983 -3379 999
rect -3413 -1071 -3379 -1055
rect -3293 983 -3259 999
rect -3293 -1071 -3259 -1055
rect -3135 983 -3101 999
rect -3135 -1071 -3101 -1055
rect -3015 983 -2981 999
rect -3015 -1071 -2981 -1055
rect -2857 983 -2823 999
rect -2857 -1071 -2823 -1055
rect -2737 983 -2703 999
rect -2737 -1071 -2703 -1055
rect -2579 983 -2545 999
rect -2579 -1071 -2545 -1055
rect -2459 983 -2425 999
rect -2459 -1071 -2425 -1055
rect -2301 983 -2267 999
rect -2301 -1071 -2267 -1055
rect -2181 983 -2147 999
rect -2181 -1071 -2147 -1055
rect -2023 983 -1989 999
rect -2023 -1071 -1989 -1055
rect -1903 983 -1869 999
rect -1903 -1071 -1869 -1055
rect -1745 983 -1711 999
rect -1745 -1071 -1711 -1055
rect -1625 983 -1591 999
rect -1625 -1071 -1591 -1055
rect -1467 983 -1433 999
rect -1467 -1071 -1433 -1055
rect -1347 983 -1313 999
rect -1347 -1071 -1313 -1055
rect -1189 983 -1155 999
rect -1189 -1071 -1155 -1055
rect -1069 983 -1035 999
rect -1069 -1071 -1035 -1055
rect -911 983 -877 999
rect -911 -1071 -877 -1055
rect -791 983 -757 999
rect -791 -1071 -757 -1055
rect -633 983 -599 999
rect -633 -1071 -599 -1055
rect -513 983 -479 999
rect -513 -1071 -479 -1055
rect -355 983 -321 999
rect -355 -1071 -321 -1055
rect -235 983 -201 999
rect -235 -1071 -201 -1055
rect -77 983 -43 999
rect -77 -1071 -43 -1055
rect 43 983 77 999
rect 43 -1071 77 -1055
rect 201 983 235 999
rect 201 -1071 235 -1055
rect 321 983 355 999
rect 321 -1071 355 -1055
rect 479 983 513 999
rect 479 -1071 513 -1055
rect 599 983 633 999
rect 599 -1071 633 -1055
rect 757 983 791 999
rect 757 -1071 791 -1055
rect 877 983 911 999
rect 877 -1071 911 -1055
rect 1035 983 1069 999
rect 1035 -1071 1069 -1055
rect 1155 983 1189 999
rect 1155 -1071 1189 -1055
rect 1313 983 1347 999
rect 1313 -1071 1347 -1055
rect 1433 983 1467 999
rect 1433 -1071 1467 -1055
rect 1591 983 1625 999
rect 1591 -1071 1625 -1055
rect 1711 983 1745 999
rect 1711 -1071 1745 -1055
rect 1869 983 1903 999
rect 1869 -1071 1903 -1055
rect 1989 983 2023 999
rect 1989 -1071 2023 -1055
rect 2147 983 2181 999
rect 2147 -1071 2181 -1055
rect 2267 983 2301 999
rect 2267 -1071 2301 -1055
rect 2425 983 2459 999
rect 2425 -1071 2459 -1055
rect 2545 983 2579 999
rect 2545 -1071 2579 -1055
rect 2703 983 2737 999
rect 2703 -1071 2737 -1055
rect 2823 983 2857 999
rect 2823 -1071 2857 -1055
rect 2981 983 3015 999
rect 2981 -1071 3015 -1055
rect 3101 983 3135 999
rect 3101 -1071 3135 -1055
rect 3259 983 3293 999
rect 3259 -1071 3293 -1055
rect 3379 983 3413 999
rect 3379 -1071 3413 -1055
rect 3537 983 3571 999
rect 3537 -1071 3571 -1055
rect 3657 983 3691 999
rect 3657 -1071 3691 -1055
rect 3815 983 3849 999
rect 3815 -1071 3849 -1055
rect 3935 983 3969 999
rect 3935 -1071 3969 -1055
rect 4093 983 4127 999
rect 4093 -1071 4127 -1055
rect 4213 983 4247 999
rect 4213 -1071 4247 -1055
rect 4371 983 4405 999
rect 4371 -1071 4405 -1055
rect 4491 983 4525 999
rect 4491 -1071 4525 -1055
rect 4649 983 4683 999
rect 4649 -1071 4683 -1055
rect 4769 983 4803 999
rect 4769 -1071 4803 -1055
rect 4927 983 4961 999
rect 4927 -1071 4961 -1055
rect 5047 983 5081 999
rect 5047 -1071 5081 -1055
rect 5205 983 5239 999
rect 5205 -1071 5239 -1055
rect 5325 983 5359 999
rect 5325 -1071 5359 -1055
rect 5483 983 5517 999
rect 5483 -1071 5517 -1055
rect 5603 983 5637 999
rect 5603 -1071 5637 -1055
rect 5761 983 5795 999
rect 5761 -1071 5795 -1055
rect 5881 983 5915 999
rect 5881 -1071 5915 -1055
rect 6039 983 6073 999
rect 6039 -1071 6073 -1055
rect 6159 983 6193 999
rect 6159 -1071 6193 -1055
rect 6317 983 6351 999
rect 6317 -1071 6351 -1055
rect 6437 983 6471 999
rect 6437 -1071 6471 -1055
rect 6595 983 6629 999
rect 6595 -1071 6629 -1055
rect 6715 983 6749 999
rect 6715 -1071 6749 -1055
rect 6873 983 6907 999
rect 6873 -1071 6907 -1055
rect 6993 983 7027 999
rect 6993 -1071 7027 -1055
rect 7151 983 7185 999
rect 7151 -1071 7185 -1055
rect 7271 983 7305 999
rect 7271 -1071 7305 -1055
rect 7429 983 7463 999
rect 7429 -1071 7463 -1055
rect 7549 983 7583 999
rect 7549 -1071 7583 -1055
rect 7707 983 7741 999
rect 7707 -1071 7741 -1055
rect 7827 983 7861 999
rect 7827 -1071 7861 -1055
rect 7985 983 8019 999
rect 7985 -1071 8019 -1055
rect 8105 983 8139 999
rect 8105 -1071 8139 -1055
rect 8263 983 8297 999
rect 8263 -1071 8297 -1055
rect 8383 983 8417 999
rect 8383 -1071 8417 -1055
rect 8541 983 8575 999
rect 8541 -1071 8575 -1055
rect 8661 983 8695 999
rect 8661 -1071 8695 -1055
rect 8819 983 8853 999
rect 8819 -1071 8853 -1055
<< viali >>
rect -8791 1042 -8723 1076
rect -8513 1042 -8445 1076
rect -8235 1042 -8167 1076
rect -7957 1042 -7889 1076
rect -7679 1042 -7611 1076
rect -7401 1042 -7333 1076
rect -7123 1042 -7055 1076
rect -6845 1042 -6777 1076
rect -6567 1042 -6499 1076
rect -6289 1042 -6221 1076
rect -6011 1042 -5943 1076
rect -5733 1042 -5665 1076
rect -5455 1042 -5387 1076
rect -5177 1042 -5109 1076
rect -4899 1042 -4831 1076
rect -4621 1042 -4553 1076
rect -4343 1042 -4275 1076
rect -4065 1042 -3997 1076
rect -3787 1042 -3719 1076
rect -3509 1042 -3441 1076
rect -3231 1042 -3163 1076
rect -2953 1042 -2885 1076
rect -2675 1042 -2607 1076
rect -2397 1042 -2329 1076
rect -2119 1042 -2051 1076
rect -1841 1042 -1773 1076
rect -1563 1042 -1495 1076
rect -1285 1042 -1217 1076
rect -1007 1042 -939 1076
rect -729 1042 -661 1076
rect -451 1042 -383 1076
rect -173 1042 -105 1076
rect 105 1042 173 1076
rect 383 1042 451 1076
rect 661 1042 729 1076
rect 939 1042 1007 1076
rect 1217 1042 1285 1076
rect 1495 1042 1563 1076
rect 1773 1042 1841 1076
rect 2051 1042 2119 1076
rect 2329 1042 2397 1076
rect 2607 1042 2675 1076
rect 2885 1042 2953 1076
rect 3163 1042 3231 1076
rect 3441 1042 3509 1076
rect 3719 1042 3787 1076
rect 3997 1042 4065 1076
rect 4275 1042 4343 1076
rect 4553 1042 4621 1076
rect 4831 1042 4899 1076
rect 5109 1042 5177 1076
rect 5387 1042 5455 1076
rect 5665 1042 5733 1076
rect 5943 1042 6011 1076
rect 6221 1042 6289 1076
rect 6499 1042 6567 1076
rect 6777 1042 6845 1076
rect 7055 1042 7123 1076
rect 7333 1042 7401 1076
rect 7611 1042 7679 1076
rect 7889 1042 7957 1076
rect 8167 1042 8235 1076
rect 8445 1042 8513 1076
rect 8723 1042 8791 1076
rect -8853 -1055 -8819 983
rect -8695 -1055 -8661 983
rect -8575 -1055 -8541 983
rect -8417 -1055 -8383 983
rect -8297 -1055 -8263 983
rect -8139 -1055 -8105 983
rect -8019 -1055 -7985 983
rect -7861 -1055 -7827 983
rect -7741 -1055 -7707 983
rect -7583 -1055 -7549 983
rect -7463 -1055 -7429 983
rect -7305 -1055 -7271 983
rect -7185 -1055 -7151 983
rect -7027 -1055 -6993 983
rect -6907 -1055 -6873 983
rect -6749 -1055 -6715 983
rect -6629 -1055 -6595 983
rect -6471 -1055 -6437 983
rect -6351 -1055 -6317 983
rect -6193 -1055 -6159 983
rect -6073 -1055 -6039 983
rect -5915 -1055 -5881 983
rect -5795 -1055 -5761 983
rect -5637 -1055 -5603 983
rect -5517 -1055 -5483 983
rect -5359 -1055 -5325 983
rect -5239 -1055 -5205 983
rect -5081 -1055 -5047 983
rect -4961 -1055 -4927 983
rect -4803 -1055 -4769 983
rect -4683 -1055 -4649 983
rect -4525 -1055 -4491 983
rect -4405 -1055 -4371 983
rect -4247 -1055 -4213 983
rect -4127 -1055 -4093 983
rect -3969 -1055 -3935 983
rect -3849 -1055 -3815 983
rect -3691 -1055 -3657 983
rect -3571 -1055 -3537 983
rect -3413 -1055 -3379 983
rect -3293 -1055 -3259 983
rect -3135 -1055 -3101 983
rect -3015 -1055 -2981 983
rect -2857 -1055 -2823 983
rect -2737 -1055 -2703 983
rect -2579 -1055 -2545 983
rect -2459 -1055 -2425 983
rect -2301 -1055 -2267 983
rect -2181 -1055 -2147 983
rect -2023 -1055 -1989 983
rect -1903 -1055 -1869 983
rect -1745 -1055 -1711 983
rect -1625 -1055 -1591 983
rect -1467 -1055 -1433 983
rect -1347 -1055 -1313 983
rect -1189 -1055 -1155 983
rect -1069 -1055 -1035 983
rect -911 -1055 -877 983
rect -791 -1055 -757 983
rect -633 -1055 -599 983
rect -513 -1055 -479 983
rect -355 -1055 -321 983
rect -235 -1055 -201 983
rect -77 -1055 -43 983
rect 43 -1055 77 983
rect 201 -1055 235 983
rect 321 -1055 355 983
rect 479 -1055 513 983
rect 599 -1055 633 983
rect 757 -1055 791 983
rect 877 -1055 911 983
rect 1035 -1055 1069 983
rect 1155 -1055 1189 983
rect 1313 -1055 1347 983
rect 1433 -1055 1467 983
rect 1591 -1055 1625 983
rect 1711 -1055 1745 983
rect 1869 -1055 1903 983
rect 1989 -1055 2023 983
rect 2147 -1055 2181 983
rect 2267 -1055 2301 983
rect 2425 -1055 2459 983
rect 2545 -1055 2579 983
rect 2703 -1055 2737 983
rect 2823 -1055 2857 983
rect 2981 -1055 3015 983
rect 3101 -1055 3135 983
rect 3259 -1055 3293 983
rect 3379 -1055 3413 983
rect 3537 -1055 3571 983
rect 3657 -1055 3691 983
rect 3815 -1055 3849 983
rect 3935 -1055 3969 983
rect 4093 -1055 4127 983
rect 4213 -1055 4247 983
rect 4371 -1055 4405 983
rect 4491 -1055 4525 983
rect 4649 -1055 4683 983
rect 4769 -1055 4803 983
rect 4927 -1055 4961 983
rect 5047 -1055 5081 983
rect 5205 -1055 5239 983
rect 5325 -1055 5359 983
rect 5483 -1055 5517 983
rect 5603 -1055 5637 983
rect 5761 -1055 5795 983
rect 5881 -1055 5915 983
rect 6039 -1055 6073 983
rect 6159 -1055 6193 983
rect 6317 -1055 6351 983
rect 6437 -1055 6471 983
rect 6595 -1055 6629 983
rect 6715 -1055 6749 983
rect 6873 -1055 6907 983
rect 6993 -1055 7027 983
rect 7151 -1055 7185 983
rect 7271 -1055 7305 983
rect 7429 -1055 7463 983
rect 7549 -1055 7583 983
rect 7707 -1055 7741 983
rect 7827 -1055 7861 983
rect 7985 -1055 8019 983
rect 8105 -1055 8139 983
rect 8263 -1055 8297 983
rect 8383 -1055 8417 983
rect 8541 -1055 8575 983
rect 8661 -1055 8695 983
rect 8819 -1055 8853 983
<< metal1 >>
rect -8803 1076 -8711 1082
rect -8803 1042 -8791 1076
rect -8723 1042 -8711 1076
rect -8803 1036 -8711 1042
rect -8525 1076 -8433 1082
rect -8525 1042 -8513 1076
rect -8445 1042 -8433 1076
rect -8525 1036 -8433 1042
rect -8247 1076 -8155 1082
rect -8247 1042 -8235 1076
rect -8167 1042 -8155 1076
rect -8247 1036 -8155 1042
rect -7969 1076 -7877 1082
rect -7969 1042 -7957 1076
rect -7889 1042 -7877 1076
rect -7969 1036 -7877 1042
rect -7691 1076 -7599 1082
rect -7691 1042 -7679 1076
rect -7611 1042 -7599 1076
rect -7691 1036 -7599 1042
rect -7413 1076 -7321 1082
rect -7413 1042 -7401 1076
rect -7333 1042 -7321 1076
rect -7413 1036 -7321 1042
rect -7135 1076 -7043 1082
rect -7135 1042 -7123 1076
rect -7055 1042 -7043 1076
rect -7135 1036 -7043 1042
rect -6857 1076 -6765 1082
rect -6857 1042 -6845 1076
rect -6777 1042 -6765 1076
rect -6857 1036 -6765 1042
rect -6579 1076 -6487 1082
rect -6579 1042 -6567 1076
rect -6499 1042 -6487 1076
rect -6579 1036 -6487 1042
rect -6301 1076 -6209 1082
rect -6301 1042 -6289 1076
rect -6221 1042 -6209 1076
rect -6301 1036 -6209 1042
rect -6023 1076 -5931 1082
rect -6023 1042 -6011 1076
rect -5943 1042 -5931 1076
rect -6023 1036 -5931 1042
rect -5745 1076 -5653 1082
rect -5745 1042 -5733 1076
rect -5665 1042 -5653 1076
rect -5745 1036 -5653 1042
rect -5467 1076 -5375 1082
rect -5467 1042 -5455 1076
rect -5387 1042 -5375 1076
rect -5467 1036 -5375 1042
rect -5189 1076 -5097 1082
rect -5189 1042 -5177 1076
rect -5109 1042 -5097 1076
rect -5189 1036 -5097 1042
rect -4911 1076 -4819 1082
rect -4911 1042 -4899 1076
rect -4831 1042 -4819 1076
rect -4911 1036 -4819 1042
rect -4633 1076 -4541 1082
rect -4633 1042 -4621 1076
rect -4553 1042 -4541 1076
rect -4633 1036 -4541 1042
rect -4355 1076 -4263 1082
rect -4355 1042 -4343 1076
rect -4275 1042 -4263 1076
rect -4355 1036 -4263 1042
rect -4077 1076 -3985 1082
rect -4077 1042 -4065 1076
rect -3997 1042 -3985 1076
rect -4077 1036 -3985 1042
rect -3799 1076 -3707 1082
rect -3799 1042 -3787 1076
rect -3719 1042 -3707 1076
rect -3799 1036 -3707 1042
rect -3521 1076 -3429 1082
rect -3521 1042 -3509 1076
rect -3441 1042 -3429 1076
rect -3521 1036 -3429 1042
rect -3243 1076 -3151 1082
rect -3243 1042 -3231 1076
rect -3163 1042 -3151 1076
rect -3243 1036 -3151 1042
rect -2965 1076 -2873 1082
rect -2965 1042 -2953 1076
rect -2885 1042 -2873 1076
rect -2965 1036 -2873 1042
rect -2687 1076 -2595 1082
rect -2687 1042 -2675 1076
rect -2607 1042 -2595 1076
rect -2687 1036 -2595 1042
rect -2409 1076 -2317 1082
rect -2409 1042 -2397 1076
rect -2329 1042 -2317 1076
rect -2409 1036 -2317 1042
rect -2131 1076 -2039 1082
rect -2131 1042 -2119 1076
rect -2051 1042 -2039 1076
rect -2131 1036 -2039 1042
rect -1853 1076 -1761 1082
rect -1853 1042 -1841 1076
rect -1773 1042 -1761 1076
rect -1853 1036 -1761 1042
rect -1575 1076 -1483 1082
rect -1575 1042 -1563 1076
rect -1495 1042 -1483 1076
rect -1575 1036 -1483 1042
rect -1297 1076 -1205 1082
rect -1297 1042 -1285 1076
rect -1217 1042 -1205 1076
rect -1297 1036 -1205 1042
rect -1019 1076 -927 1082
rect -1019 1042 -1007 1076
rect -939 1042 -927 1076
rect -1019 1036 -927 1042
rect -741 1076 -649 1082
rect -741 1042 -729 1076
rect -661 1042 -649 1076
rect -741 1036 -649 1042
rect -463 1076 -371 1082
rect -463 1042 -451 1076
rect -383 1042 -371 1076
rect -463 1036 -371 1042
rect -185 1076 -93 1082
rect -185 1042 -173 1076
rect -105 1042 -93 1076
rect -185 1036 -93 1042
rect 93 1076 185 1082
rect 93 1042 105 1076
rect 173 1042 185 1076
rect 93 1036 185 1042
rect 371 1076 463 1082
rect 371 1042 383 1076
rect 451 1042 463 1076
rect 371 1036 463 1042
rect 649 1076 741 1082
rect 649 1042 661 1076
rect 729 1042 741 1076
rect 649 1036 741 1042
rect 927 1076 1019 1082
rect 927 1042 939 1076
rect 1007 1042 1019 1076
rect 927 1036 1019 1042
rect 1205 1076 1297 1082
rect 1205 1042 1217 1076
rect 1285 1042 1297 1076
rect 1205 1036 1297 1042
rect 1483 1076 1575 1082
rect 1483 1042 1495 1076
rect 1563 1042 1575 1076
rect 1483 1036 1575 1042
rect 1761 1076 1853 1082
rect 1761 1042 1773 1076
rect 1841 1042 1853 1076
rect 1761 1036 1853 1042
rect 2039 1076 2131 1082
rect 2039 1042 2051 1076
rect 2119 1042 2131 1076
rect 2039 1036 2131 1042
rect 2317 1076 2409 1082
rect 2317 1042 2329 1076
rect 2397 1042 2409 1076
rect 2317 1036 2409 1042
rect 2595 1076 2687 1082
rect 2595 1042 2607 1076
rect 2675 1042 2687 1076
rect 2595 1036 2687 1042
rect 2873 1076 2965 1082
rect 2873 1042 2885 1076
rect 2953 1042 2965 1076
rect 2873 1036 2965 1042
rect 3151 1076 3243 1082
rect 3151 1042 3163 1076
rect 3231 1042 3243 1076
rect 3151 1036 3243 1042
rect 3429 1076 3521 1082
rect 3429 1042 3441 1076
rect 3509 1042 3521 1076
rect 3429 1036 3521 1042
rect 3707 1076 3799 1082
rect 3707 1042 3719 1076
rect 3787 1042 3799 1076
rect 3707 1036 3799 1042
rect 3985 1076 4077 1082
rect 3985 1042 3997 1076
rect 4065 1042 4077 1076
rect 3985 1036 4077 1042
rect 4263 1076 4355 1082
rect 4263 1042 4275 1076
rect 4343 1042 4355 1076
rect 4263 1036 4355 1042
rect 4541 1076 4633 1082
rect 4541 1042 4553 1076
rect 4621 1042 4633 1076
rect 4541 1036 4633 1042
rect 4819 1076 4911 1082
rect 4819 1042 4831 1076
rect 4899 1042 4911 1076
rect 4819 1036 4911 1042
rect 5097 1076 5189 1082
rect 5097 1042 5109 1076
rect 5177 1042 5189 1076
rect 5097 1036 5189 1042
rect 5375 1076 5467 1082
rect 5375 1042 5387 1076
rect 5455 1042 5467 1076
rect 5375 1036 5467 1042
rect 5653 1076 5745 1082
rect 5653 1042 5665 1076
rect 5733 1042 5745 1076
rect 5653 1036 5745 1042
rect 5931 1076 6023 1082
rect 5931 1042 5943 1076
rect 6011 1042 6023 1076
rect 5931 1036 6023 1042
rect 6209 1076 6301 1082
rect 6209 1042 6221 1076
rect 6289 1042 6301 1076
rect 6209 1036 6301 1042
rect 6487 1076 6579 1082
rect 6487 1042 6499 1076
rect 6567 1042 6579 1076
rect 6487 1036 6579 1042
rect 6765 1076 6857 1082
rect 6765 1042 6777 1076
rect 6845 1042 6857 1076
rect 6765 1036 6857 1042
rect 7043 1076 7135 1082
rect 7043 1042 7055 1076
rect 7123 1042 7135 1076
rect 7043 1036 7135 1042
rect 7321 1076 7413 1082
rect 7321 1042 7333 1076
rect 7401 1042 7413 1076
rect 7321 1036 7413 1042
rect 7599 1076 7691 1082
rect 7599 1042 7611 1076
rect 7679 1042 7691 1076
rect 7599 1036 7691 1042
rect 7877 1076 7969 1082
rect 7877 1042 7889 1076
rect 7957 1042 7969 1076
rect 7877 1036 7969 1042
rect 8155 1076 8247 1082
rect 8155 1042 8167 1076
rect 8235 1042 8247 1076
rect 8155 1036 8247 1042
rect 8433 1076 8525 1082
rect 8433 1042 8445 1076
rect 8513 1042 8525 1076
rect 8433 1036 8525 1042
rect 8711 1076 8803 1082
rect 8711 1042 8723 1076
rect 8791 1042 8803 1076
rect 8711 1036 8803 1042
rect -8859 983 -8813 995
rect -8859 -1055 -8853 983
rect -8819 -1055 -8813 983
rect -8859 -1067 -8813 -1055
rect -8701 983 -8655 995
rect -8701 -1055 -8695 983
rect -8661 -1055 -8655 983
rect -8701 -1067 -8655 -1055
rect -8581 983 -8535 995
rect -8581 -1055 -8575 983
rect -8541 -1055 -8535 983
rect -8581 -1067 -8535 -1055
rect -8423 983 -8377 995
rect -8423 -1055 -8417 983
rect -8383 -1055 -8377 983
rect -8423 -1067 -8377 -1055
rect -8303 983 -8257 995
rect -8303 -1055 -8297 983
rect -8263 -1055 -8257 983
rect -8303 -1067 -8257 -1055
rect -8145 983 -8099 995
rect -8145 -1055 -8139 983
rect -8105 -1055 -8099 983
rect -8145 -1067 -8099 -1055
rect -8025 983 -7979 995
rect -8025 -1055 -8019 983
rect -7985 -1055 -7979 983
rect -8025 -1067 -7979 -1055
rect -7867 983 -7821 995
rect -7867 -1055 -7861 983
rect -7827 -1055 -7821 983
rect -7867 -1067 -7821 -1055
rect -7747 983 -7701 995
rect -7747 -1055 -7741 983
rect -7707 -1055 -7701 983
rect -7747 -1067 -7701 -1055
rect -7589 983 -7543 995
rect -7589 -1055 -7583 983
rect -7549 -1055 -7543 983
rect -7589 -1067 -7543 -1055
rect -7469 983 -7423 995
rect -7469 -1055 -7463 983
rect -7429 -1055 -7423 983
rect -7469 -1067 -7423 -1055
rect -7311 983 -7265 995
rect -7311 -1055 -7305 983
rect -7271 -1055 -7265 983
rect -7311 -1067 -7265 -1055
rect -7191 983 -7145 995
rect -7191 -1055 -7185 983
rect -7151 -1055 -7145 983
rect -7191 -1067 -7145 -1055
rect -7033 983 -6987 995
rect -7033 -1055 -7027 983
rect -6993 -1055 -6987 983
rect -7033 -1067 -6987 -1055
rect -6913 983 -6867 995
rect -6913 -1055 -6907 983
rect -6873 -1055 -6867 983
rect -6913 -1067 -6867 -1055
rect -6755 983 -6709 995
rect -6755 -1055 -6749 983
rect -6715 -1055 -6709 983
rect -6755 -1067 -6709 -1055
rect -6635 983 -6589 995
rect -6635 -1055 -6629 983
rect -6595 -1055 -6589 983
rect -6635 -1067 -6589 -1055
rect -6477 983 -6431 995
rect -6477 -1055 -6471 983
rect -6437 -1055 -6431 983
rect -6477 -1067 -6431 -1055
rect -6357 983 -6311 995
rect -6357 -1055 -6351 983
rect -6317 -1055 -6311 983
rect -6357 -1067 -6311 -1055
rect -6199 983 -6153 995
rect -6199 -1055 -6193 983
rect -6159 -1055 -6153 983
rect -6199 -1067 -6153 -1055
rect -6079 983 -6033 995
rect -6079 -1055 -6073 983
rect -6039 -1055 -6033 983
rect -6079 -1067 -6033 -1055
rect -5921 983 -5875 995
rect -5921 -1055 -5915 983
rect -5881 -1055 -5875 983
rect -5921 -1067 -5875 -1055
rect -5801 983 -5755 995
rect -5801 -1055 -5795 983
rect -5761 -1055 -5755 983
rect -5801 -1067 -5755 -1055
rect -5643 983 -5597 995
rect -5643 -1055 -5637 983
rect -5603 -1055 -5597 983
rect -5643 -1067 -5597 -1055
rect -5523 983 -5477 995
rect -5523 -1055 -5517 983
rect -5483 -1055 -5477 983
rect -5523 -1067 -5477 -1055
rect -5365 983 -5319 995
rect -5365 -1055 -5359 983
rect -5325 -1055 -5319 983
rect -5365 -1067 -5319 -1055
rect -5245 983 -5199 995
rect -5245 -1055 -5239 983
rect -5205 -1055 -5199 983
rect -5245 -1067 -5199 -1055
rect -5087 983 -5041 995
rect -5087 -1055 -5081 983
rect -5047 -1055 -5041 983
rect -5087 -1067 -5041 -1055
rect -4967 983 -4921 995
rect -4967 -1055 -4961 983
rect -4927 -1055 -4921 983
rect -4967 -1067 -4921 -1055
rect -4809 983 -4763 995
rect -4809 -1055 -4803 983
rect -4769 -1055 -4763 983
rect -4809 -1067 -4763 -1055
rect -4689 983 -4643 995
rect -4689 -1055 -4683 983
rect -4649 -1055 -4643 983
rect -4689 -1067 -4643 -1055
rect -4531 983 -4485 995
rect -4531 -1055 -4525 983
rect -4491 -1055 -4485 983
rect -4531 -1067 -4485 -1055
rect -4411 983 -4365 995
rect -4411 -1055 -4405 983
rect -4371 -1055 -4365 983
rect -4411 -1067 -4365 -1055
rect -4253 983 -4207 995
rect -4253 -1055 -4247 983
rect -4213 -1055 -4207 983
rect -4253 -1067 -4207 -1055
rect -4133 983 -4087 995
rect -4133 -1055 -4127 983
rect -4093 -1055 -4087 983
rect -4133 -1067 -4087 -1055
rect -3975 983 -3929 995
rect -3975 -1055 -3969 983
rect -3935 -1055 -3929 983
rect -3975 -1067 -3929 -1055
rect -3855 983 -3809 995
rect -3855 -1055 -3849 983
rect -3815 -1055 -3809 983
rect -3855 -1067 -3809 -1055
rect -3697 983 -3651 995
rect -3697 -1055 -3691 983
rect -3657 -1055 -3651 983
rect -3697 -1067 -3651 -1055
rect -3577 983 -3531 995
rect -3577 -1055 -3571 983
rect -3537 -1055 -3531 983
rect -3577 -1067 -3531 -1055
rect -3419 983 -3373 995
rect -3419 -1055 -3413 983
rect -3379 -1055 -3373 983
rect -3419 -1067 -3373 -1055
rect -3299 983 -3253 995
rect -3299 -1055 -3293 983
rect -3259 -1055 -3253 983
rect -3299 -1067 -3253 -1055
rect -3141 983 -3095 995
rect -3141 -1055 -3135 983
rect -3101 -1055 -3095 983
rect -3141 -1067 -3095 -1055
rect -3021 983 -2975 995
rect -3021 -1055 -3015 983
rect -2981 -1055 -2975 983
rect -3021 -1067 -2975 -1055
rect -2863 983 -2817 995
rect -2863 -1055 -2857 983
rect -2823 -1055 -2817 983
rect -2863 -1067 -2817 -1055
rect -2743 983 -2697 995
rect -2743 -1055 -2737 983
rect -2703 -1055 -2697 983
rect -2743 -1067 -2697 -1055
rect -2585 983 -2539 995
rect -2585 -1055 -2579 983
rect -2545 -1055 -2539 983
rect -2585 -1067 -2539 -1055
rect -2465 983 -2419 995
rect -2465 -1055 -2459 983
rect -2425 -1055 -2419 983
rect -2465 -1067 -2419 -1055
rect -2307 983 -2261 995
rect -2307 -1055 -2301 983
rect -2267 -1055 -2261 983
rect -2307 -1067 -2261 -1055
rect -2187 983 -2141 995
rect -2187 -1055 -2181 983
rect -2147 -1055 -2141 983
rect -2187 -1067 -2141 -1055
rect -2029 983 -1983 995
rect -2029 -1055 -2023 983
rect -1989 -1055 -1983 983
rect -2029 -1067 -1983 -1055
rect -1909 983 -1863 995
rect -1909 -1055 -1903 983
rect -1869 -1055 -1863 983
rect -1909 -1067 -1863 -1055
rect -1751 983 -1705 995
rect -1751 -1055 -1745 983
rect -1711 -1055 -1705 983
rect -1751 -1067 -1705 -1055
rect -1631 983 -1585 995
rect -1631 -1055 -1625 983
rect -1591 -1055 -1585 983
rect -1631 -1067 -1585 -1055
rect -1473 983 -1427 995
rect -1473 -1055 -1467 983
rect -1433 -1055 -1427 983
rect -1473 -1067 -1427 -1055
rect -1353 983 -1307 995
rect -1353 -1055 -1347 983
rect -1313 -1055 -1307 983
rect -1353 -1067 -1307 -1055
rect -1195 983 -1149 995
rect -1195 -1055 -1189 983
rect -1155 -1055 -1149 983
rect -1195 -1067 -1149 -1055
rect -1075 983 -1029 995
rect -1075 -1055 -1069 983
rect -1035 -1055 -1029 983
rect -1075 -1067 -1029 -1055
rect -917 983 -871 995
rect -917 -1055 -911 983
rect -877 -1055 -871 983
rect -917 -1067 -871 -1055
rect -797 983 -751 995
rect -797 -1055 -791 983
rect -757 -1055 -751 983
rect -797 -1067 -751 -1055
rect -639 983 -593 995
rect -639 -1055 -633 983
rect -599 -1055 -593 983
rect -639 -1067 -593 -1055
rect -519 983 -473 995
rect -519 -1055 -513 983
rect -479 -1055 -473 983
rect -519 -1067 -473 -1055
rect -361 983 -315 995
rect -361 -1055 -355 983
rect -321 -1055 -315 983
rect -361 -1067 -315 -1055
rect -241 983 -195 995
rect -241 -1055 -235 983
rect -201 -1055 -195 983
rect -241 -1067 -195 -1055
rect -83 983 -37 995
rect -83 -1055 -77 983
rect -43 -1055 -37 983
rect -83 -1067 -37 -1055
rect 37 983 83 995
rect 37 -1055 43 983
rect 77 -1055 83 983
rect 37 -1067 83 -1055
rect 195 983 241 995
rect 195 -1055 201 983
rect 235 -1055 241 983
rect 195 -1067 241 -1055
rect 315 983 361 995
rect 315 -1055 321 983
rect 355 -1055 361 983
rect 315 -1067 361 -1055
rect 473 983 519 995
rect 473 -1055 479 983
rect 513 -1055 519 983
rect 473 -1067 519 -1055
rect 593 983 639 995
rect 593 -1055 599 983
rect 633 -1055 639 983
rect 593 -1067 639 -1055
rect 751 983 797 995
rect 751 -1055 757 983
rect 791 -1055 797 983
rect 751 -1067 797 -1055
rect 871 983 917 995
rect 871 -1055 877 983
rect 911 -1055 917 983
rect 871 -1067 917 -1055
rect 1029 983 1075 995
rect 1029 -1055 1035 983
rect 1069 -1055 1075 983
rect 1029 -1067 1075 -1055
rect 1149 983 1195 995
rect 1149 -1055 1155 983
rect 1189 -1055 1195 983
rect 1149 -1067 1195 -1055
rect 1307 983 1353 995
rect 1307 -1055 1313 983
rect 1347 -1055 1353 983
rect 1307 -1067 1353 -1055
rect 1427 983 1473 995
rect 1427 -1055 1433 983
rect 1467 -1055 1473 983
rect 1427 -1067 1473 -1055
rect 1585 983 1631 995
rect 1585 -1055 1591 983
rect 1625 -1055 1631 983
rect 1585 -1067 1631 -1055
rect 1705 983 1751 995
rect 1705 -1055 1711 983
rect 1745 -1055 1751 983
rect 1705 -1067 1751 -1055
rect 1863 983 1909 995
rect 1863 -1055 1869 983
rect 1903 -1055 1909 983
rect 1863 -1067 1909 -1055
rect 1983 983 2029 995
rect 1983 -1055 1989 983
rect 2023 -1055 2029 983
rect 1983 -1067 2029 -1055
rect 2141 983 2187 995
rect 2141 -1055 2147 983
rect 2181 -1055 2187 983
rect 2141 -1067 2187 -1055
rect 2261 983 2307 995
rect 2261 -1055 2267 983
rect 2301 -1055 2307 983
rect 2261 -1067 2307 -1055
rect 2419 983 2465 995
rect 2419 -1055 2425 983
rect 2459 -1055 2465 983
rect 2419 -1067 2465 -1055
rect 2539 983 2585 995
rect 2539 -1055 2545 983
rect 2579 -1055 2585 983
rect 2539 -1067 2585 -1055
rect 2697 983 2743 995
rect 2697 -1055 2703 983
rect 2737 -1055 2743 983
rect 2697 -1067 2743 -1055
rect 2817 983 2863 995
rect 2817 -1055 2823 983
rect 2857 -1055 2863 983
rect 2817 -1067 2863 -1055
rect 2975 983 3021 995
rect 2975 -1055 2981 983
rect 3015 -1055 3021 983
rect 2975 -1067 3021 -1055
rect 3095 983 3141 995
rect 3095 -1055 3101 983
rect 3135 -1055 3141 983
rect 3095 -1067 3141 -1055
rect 3253 983 3299 995
rect 3253 -1055 3259 983
rect 3293 -1055 3299 983
rect 3253 -1067 3299 -1055
rect 3373 983 3419 995
rect 3373 -1055 3379 983
rect 3413 -1055 3419 983
rect 3373 -1067 3419 -1055
rect 3531 983 3577 995
rect 3531 -1055 3537 983
rect 3571 -1055 3577 983
rect 3531 -1067 3577 -1055
rect 3651 983 3697 995
rect 3651 -1055 3657 983
rect 3691 -1055 3697 983
rect 3651 -1067 3697 -1055
rect 3809 983 3855 995
rect 3809 -1055 3815 983
rect 3849 -1055 3855 983
rect 3809 -1067 3855 -1055
rect 3929 983 3975 995
rect 3929 -1055 3935 983
rect 3969 -1055 3975 983
rect 3929 -1067 3975 -1055
rect 4087 983 4133 995
rect 4087 -1055 4093 983
rect 4127 -1055 4133 983
rect 4087 -1067 4133 -1055
rect 4207 983 4253 995
rect 4207 -1055 4213 983
rect 4247 -1055 4253 983
rect 4207 -1067 4253 -1055
rect 4365 983 4411 995
rect 4365 -1055 4371 983
rect 4405 -1055 4411 983
rect 4365 -1067 4411 -1055
rect 4485 983 4531 995
rect 4485 -1055 4491 983
rect 4525 -1055 4531 983
rect 4485 -1067 4531 -1055
rect 4643 983 4689 995
rect 4643 -1055 4649 983
rect 4683 -1055 4689 983
rect 4643 -1067 4689 -1055
rect 4763 983 4809 995
rect 4763 -1055 4769 983
rect 4803 -1055 4809 983
rect 4763 -1067 4809 -1055
rect 4921 983 4967 995
rect 4921 -1055 4927 983
rect 4961 -1055 4967 983
rect 4921 -1067 4967 -1055
rect 5041 983 5087 995
rect 5041 -1055 5047 983
rect 5081 -1055 5087 983
rect 5041 -1067 5087 -1055
rect 5199 983 5245 995
rect 5199 -1055 5205 983
rect 5239 -1055 5245 983
rect 5199 -1067 5245 -1055
rect 5319 983 5365 995
rect 5319 -1055 5325 983
rect 5359 -1055 5365 983
rect 5319 -1067 5365 -1055
rect 5477 983 5523 995
rect 5477 -1055 5483 983
rect 5517 -1055 5523 983
rect 5477 -1067 5523 -1055
rect 5597 983 5643 995
rect 5597 -1055 5603 983
rect 5637 -1055 5643 983
rect 5597 -1067 5643 -1055
rect 5755 983 5801 995
rect 5755 -1055 5761 983
rect 5795 -1055 5801 983
rect 5755 -1067 5801 -1055
rect 5875 983 5921 995
rect 5875 -1055 5881 983
rect 5915 -1055 5921 983
rect 5875 -1067 5921 -1055
rect 6033 983 6079 995
rect 6033 -1055 6039 983
rect 6073 -1055 6079 983
rect 6033 -1067 6079 -1055
rect 6153 983 6199 995
rect 6153 -1055 6159 983
rect 6193 -1055 6199 983
rect 6153 -1067 6199 -1055
rect 6311 983 6357 995
rect 6311 -1055 6317 983
rect 6351 -1055 6357 983
rect 6311 -1067 6357 -1055
rect 6431 983 6477 995
rect 6431 -1055 6437 983
rect 6471 -1055 6477 983
rect 6431 -1067 6477 -1055
rect 6589 983 6635 995
rect 6589 -1055 6595 983
rect 6629 -1055 6635 983
rect 6589 -1067 6635 -1055
rect 6709 983 6755 995
rect 6709 -1055 6715 983
rect 6749 -1055 6755 983
rect 6709 -1067 6755 -1055
rect 6867 983 6913 995
rect 6867 -1055 6873 983
rect 6907 -1055 6913 983
rect 6867 -1067 6913 -1055
rect 6987 983 7033 995
rect 6987 -1055 6993 983
rect 7027 -1055 7033 983
rect 6987 -1067 7033 -1055
rect 7145 983 7191 995
rect 7145 -1055 7151 983
rect 7185 -1055 7191 983
rect 7145 -1067 7191 -1055
rect 7265 983 7311 995
rect 7265 -1055 7271 983
rect 7305 -1055 7311 983
rect 7265 -1067 7311 -1055
rect 7423 983 7469 995
rect 7423 -1055 7429 983
rect 7463 -1055 7469 983
rect 7423 -1067 7469 -1055
rect 7543 983 7589 995
rect 7543 -1055 7549 983
rect 7583 -1055 7589 983
rect 7543 -1067 7589 -1055
rect 7701 983 7747 995
rect 7701 -1055 7707 983
rect 7741 -1055 7747 983
rect 7701 -1067 7747 -1055
rect 7821 983 7867 995
rect 7821 -1055 7827 983
rect 7861 -1055 7867 983
rect 7821 -1067 7867 -1055
rect 7979 983 8025 995
rect 7979 -1055 7985 983
rect 8019 -1055 8025 983
rect 7979 -1067 8025 -1055
rect 8099 983 8145 995
rect 8099 -1055 8105 983
rect 8139 -1055 8145 983
rect 8099 -1067 8145 -1055
rect 8257 983 8303 995
rect 8257 -1055 8263 983
rect 8297 -1055 8303 983
rect 8257 -1067 8303 -1055
rect 8377 983 8423 995
rect 8377 -1055 8383 983
rect 8417 -1055 8423 983
rect 8377 -1067 8423 -1055
rect 8535 983 8581 995
rect 8535 -1055 8541 983
rect 8575 -1055 8581 983
rect 8535 -1067 8581 -1055
rect 8655 983 8701 995
rect 8655 -1055 8661 983
rect 8695 -1055 8701 983
rect 8655 -1067 8701 -1055
rect 8813 983 8859 995
rect 8813 -1055 8819 983
rect 8853 -1055 8859 983
rect 8813 -1067 8859 -1055
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.3125 l 0.5 m 1 nf 64 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
