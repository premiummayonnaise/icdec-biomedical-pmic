magic
tech sky130A
magscale 1 2
timestamp 1769411983
<< mvnmos >>
rect -2435 -781 -2185 719
rect -2127 -781 -1877 719
rect -1819 -781 -1569 719
rect -1511 -781 -1261 719
rect -1203 -781 -953 719
rect -895 -781 -645 719
rect -587 -781 -337 719
rect -279 -781 -29 719
rect 29 -781 279 719
rect 337 -781 587 719
rect 645 -781 895 719
rect 953 -781 1203 719
rect 1261 -781 1511 719
rect 1569 -781 1819 719
rect 1877 -781 2127 719
rect 2185 -781 2435 719
<< mvndiff >>
rect -2493 707 -2435 719
rect -2493 -769 -2481 707
rect -2447 -769 -2435 707
rect -2493 -781 -2435 -769
rect -2185 707 -2127 719
rect -2185 -769 -2173 707
rect -2139 -769 -2127 707
rect -2185 -781 -2127 -769
rect -1877 707 -1819 719
rect -1877 -769 -1865 707
rect -1831 -769 -1819 707
rect -1877 -781 -1819 -769
rect -1569 707 -1511 719
rect -1569 -769 -1557 707
rect -1523 -769 -1511 707
rect -1569 -781 -1511 -769
rect -1261 707 -1203 719
rect -1261 -769 -1249 707
rect -1215 -769 -1203 707
rect -1261 -781 -1203 -769
rect -953 707 -895 719
rect -953 -769 -941 707
rect -907 -769 -895 707
rect -953 -781 -895 -769
rect -645 707 -587 719
rect -645 -769 -633 707
rect -599 -769 -587 707
rect -645 -781 -587 -769
rect -337 707 -279 719
rect -337 -769 -325 707
rect -291 -769 -279 707
rect -337 -781 -279 -769
rect -29 707 29 719
rect -29 -769 -17 707
rect 17 -769 29 707
rect -29 -781 29 -769
rect 279 707 337 719
rect 279 -769 291 707
rect 325 -769 337 707
rect 279 -781 337 -769
rect 587 707 645 719
rect 587 -769 599 707
rect 633 -769 645 707
rect 587 -781 645 -769
rect 895 707 953 719
rect 895 -769 907 707
rect 941 -769 953 707
rect 895 -781 953 -769
rect 1203 707 1261 719
rect 1203 -769 1215 707
rect 1249 -769 1261 707
rect 1203 -781 1261 -769
rect 1511 707 1569 719
rect 1511 -769 1523 707
rect 1557 -769 1569 707
rect 1511 -781 1569 -769
rect 1819 707 1877 719
rect 1819 -769 1831 707
rect 1865 -769 1877 707
rect 1819 -781 1877 -769
rect 2127 707 2185 719
rect 2127 -769 2139 707
rect 2173 -769 2185 707
rect 2127 -781 2185 -769
rect 2435 707 2493 719
rect 2435 -769 2447 707
rect 2481 -769 2493 707
rect 2435 -781 2493 -769
<< mvndiffc >>
rect -2481 -769 -2447 707
rect -2173 -769 -2139 707
rect -1865 -769 -1831 707
rect -1557 -769 -1523 707
rect -1249 -769 -1215 707
rect -941 -769 -907 707
rect -633 -769 -599 707
rect -325 -769 -291 707
rect -17 -769 17 707
rect 291 -769 325 707
rect 599 -769 633 707
rect 907 -769 941 707
rect 1215 -769 1249 707
rect 1523 -769 1557 707
rect 1831 -769 1865 707
rect 2139 -769 2173 707
rect 2447 -769 2481 707
<< poly >>
rect -2435 791 -2185 807
rect -2435 757 -2419 791
rect -2201 757 -2185 791
rect -2435 719 -2185 757
rect -2127 791 -1877 807
rect -2127 757 -2111 791
rect -1893 757 -1877 791
rect -2127 719 -1877 757
rect -1819 791 -1569 807
rect -1819 757 -1803 791
rect -1585 757 -1569 791
rect -1819 719 -1569 757
rect -1511 791 -1261 807
rect -1511 757 -1495 791
rect -1277 757 -1261 791
rect -1511 719 -1261 757
rect -1203 791 -953 807
rect -1203 757 -1187 791
rect -969 757 -953 791
rect -1203 719 -953 757
rect -895 791 -645 807
rect -895 757 -879 791
rect -661 757 -645 791
rect -895 719 -645 757
rect -587 791 -337 807
rect -587 757 -571 791
rect -353 757 -337 791
rect -587 719 -337 757
rect -279 791 -29 807
rect -279 757 -263 791
rect -45 757 -29 791
rect -279 719 -29 757
rect 29 791 279 807
rect 29 757 45 791
rect 263 757 279 791
rect 29 719 279 757
rect 337 791 587 807
rect 337 757 353 791
rect 571 757 587 791
rect 337 719 587 757
rect 645 791 895 807
rect 645 757 661 791
rect 879 757 895 791
rect 645 719 895 757
rect 953 791 1203 807
rect 953 757 969 791
rect 1187 757 1203 791
rect 953 719 1203 757
rect 1261 791 1511 807
rect 1261 757 1277 791
rect 1495 757 1511 791
rect 1261 719 1511 757
rect 1569 791 1819 807
rect 1569 757 1585 791
rect 1803 757 1819 791
rect 1569 719 1819 757
rect 1877 791 2127 807
rect 1877 757 1893 791
rect 2111 757 2127 791
rect 1877 719 2127 757
rect 2185 791 2435 807
rect 2185 757 2201 791
rect 2419 757 2435 791
rect 2185 719 2435 757
rect -2435 -807 -2185 -781
rect -2127 -807 -1877 -781
rect -1819 -807 -1569 -781
rect -1511 -807 -1261 -781
rect -1203 -807 -953 -781
rect -895 -807 -645 -781
rect -587 -807 -337 -781
rect -279 -807 -29 -781
rect 29 -807 279 -781
rect 337 -807 587 -781
rect 645 -807 895 -781
rect 953 -807 1203 -781
rect 1261 -807 1511 -781
rect 1569 -807 1819 -781
rect 1877 -807 2127 -781
rect 2185 -807 2435 -781
<< polycont >>
rect -2419 757 -2201 791
rect -2111 757 -1893 791
rect -1803 757 -1585 791
rect -1495 757 -1277 791
rect -1187 757 -969 791
rect -879 757 -661 791
rect -571 757 -353 791
rect -263 757 -45 791
rect 45 757 263 791
rect 353 757 571 791
rect 661 757 879 791
rect 969 757 1187 791
rect 1277 757 1495 791
rect 1585 757 1803 791
rect 1893 757 2111 791
rect 2201 757 2419 791
<< locali >>
rect -2435 757 -2419 791
rect -2201 757 -2185 791
rect -2127 757 -2111 791
rect -1893 757 -1877 791
rect -1819 757 -1803 791
rect -1585 757 -1569 791
rect -1511 757 -1495 791
rect -1277 757 -1261 791
rect -1203 757 -1187 791
rect -969 757 -953 791
rect -895 757 -879 791
rect -661 757 -645 791
rect -587 757 -571 791
rect -353 757 -337 791
rect -279 757 -263 791
rect -45 757 -29 791
rect 29 757 45 791
rect 263 757 279 791
rect 337 757 353 791
rect 571 757 587 791
rect 645 757 661 791
rect 879 757 895 791
rect 953 757 969 791
rect 1187 757 1203 791
rect 1261 757 1277 791
rect 1495 757 1511 791
rect 1569 757 1585 791
rect 1803 757 1819 791
rect 1877 757 1893 791
rect 2111 757 2127 791
rect 2185 757 2201 791
rect 2419 757 2435 791
rect -2481 707 -2447 723
rect -2481 -785 -2447 -769
rect -2173 707 -2139 723
rect -2173 -785 -2139 -769
rect -1865 707 -1831 723
rect -1865 -785 -1831 -769
rect -1557 707 -1523 723
rect -1557 -785 -1523 -769
rect -1249 707 -1215 723
rect -1249 -785 -1215 -769
rect -941 707 -907 723
rect -941 -785 -907 -769
rect -633 707 -599 723
rect -633 -785 -599 -769
rect -325 707 -291 723
rect -325 -785 -291 -769
rect -17 707 17 723
rect -17 -785 17 -769
rect 291 707 325 723
rect 291 -785 325 -769
rect 599 707 633 723
rect 599 -785 633 -769
rect 907 707 941 723
rect 907 -785 941 -769
rect 1215 707 1249 723
rect 1215 -785 1249 -769
rect 1523 707 1557 723
rect 1523 -785 1557 -769
rect 1831 707 1865 723
rect 1831 -785 1865 -769
rect 2139 707 2173 723
rect 2139 -785 2173 -769
rect 2447 707 2481 723
rect 2447 -785 2481 -769
<< viali >>
rect -2419 757 -2201 791
rect -2111 757 -1893 791
rect -1803 757 -1585 791
rect -1495 757 -1277 791
rect -1187 757 -969 791
rect -879 757 -661 791
rect -571 757 -353 791
rect -263 757 -45 791
rect 45 757 263 791
rect 353 757 571 791
rect 661 757 879 791
rect 969 757 1187 791
rect 1277 757 1495 791
rect 1585 757 1803 791
rect 1893 757 2111 791
rect 2201 757 2419 791
rect -2481 -769 -2447 707
rect -2173 -769 -2139 707
rect -1865 -769 -1831 707
rect -1557 -769 -1523 707
rect -1249 -769 -1215 707
rect -941 -769 -907 707
rect -633 -769 -599 707
rect -325 -769 -291 707
rect -17 -769 17 707
rect 291 -769 325 707
rect 599 -769 633 707
rect 907 -769 941 707
rect 1215 -769 1249 707
rect 1523 -769 1557 707
rect 1831 -769 1865 707
rect 2139 -769 2173 707
rect 2447 -769 2481 707
<< metal1 >>
rect -2431 791 -2189 797
rect -2431 757 -2419 791
rect -2201 757 -2189 791
rect -2431 751 -2189 757
rect -2123 791 -1881 797
rect -2123 757 -2111 791
rect -1893 757 -1881 791
rect -2123 751 -1881 757
rect -1815 791 -1573 797
rect -1815 757 -1803 791
rect -1585 757 -1573 791
rect -1815 751 -1573 757
rect -1507 791 -1265 797
rect -1507 757 -1495 791
rect -1277 757 -1265 791
rect -1507 751 -1265 757
rect -1199 791 -957 797
rect -1199 757 -1187 791
rect -969 757 -957 791
rect -1199 751 -957 757
rect -891 791 -649 797
rect -891 757 -879 791
rect -661 757 -649 791
rect -891 751 -649 757
rect -583 791 -341 797
rect -583 757 -571 791
rect -353 757 -341 791
rect -583 751 -341 757
rect -275 791 -33 797
rect -275 757 -263 791
rect -45 757 -33 791
rect -275 751 -33 757
rect 33 791 275 797
rect 33 757 45 791
rect 263 757 275 791
rect 33 751 275 757
rect 341 791 583 797
rect 341 757 353 791
rect 571 757 583 791
rect 341 751 583 757
rect 649 791 891 797
rect 649 757 661 791
rect 879 757 891 791
rect 649 751 891 757
rect 957 791 1199 797
rect 957 757 969 791
rect 1187 757 1199 791
rect 957 751 1199 757
rect 1265 791 1507 797
rect 1265 757 1277 791
rect 1495 757 1507 791
rect 1265 751 1507 757
rect 1573 791 1815 797
rect 1573 757 1585 791
rect 1803 757 1815 791
rect 1573 751 1815 757
rect 1881 791 2123 797
rect 1881 757 1893 791
rect 2111 757 2123 791
rect 1881 751 2123 757
rect 2189 791 2431 797
rect 2189 757 2201 791
rect 2419 757 2431 791
rect 2189 751 2431 757
rect -2487 707 -2441 719
rect -2487 -769 -2481 707
rect -2447 -769 -2441 707
rect -2487 -781 -2441 -769
rect -2179 707 -2133 719
rect -2179 -769 -2173 707
rect -2139 -769 -2133 707
rect -2179 -781 -2133 -769
rect -1871 707 -1825 719
rect -1871 -769 -1865 707
rect -1831 -769 -1825 707
rect -1871 -781 -1825 -769
rect -1563 707 -1517 719
rect -1563 -769 -1557 707
rect -1523 -769 -1517 707
rect -1563 -781 -1517 -769
rect -1255 707 -1209 719
rect -1255 -769 -1249 707
rect -1215 -769 -1209 707
rect -1255 -781 -1209 -769
rect -947 707 -901 719
rect -947 -769 -941 707
rect -907 -769 -901 707
rect -947 -781 -901 -769
rect -639 707 -593 719
rect -639 -769 -633 707
rect -599 -769 -593 707
rect -639 -781 -593 -769
rect -331 707 -285 719
rect -331 -769 -325 707
rect -291 -769 -285 707
rect -331 -781 -285 -769
rect -23 707 23 719
rect -23 -769 -17 707
rect 17 -769 23 707
rect -23 -781 23 -769
rect 285 707 331 719
rect 285 -769 291 707
rect 325 -769 331 707
rect 285 -781 331 -769
rect 593 707 639 719
rect 593 -769 599 707
rect 633 -769 639 707
rect 593 -781 639 -769
rect 901 707 947 719
rect 901 -769 907 707
rect 941 -769 947 707
rect 901 -781 947 -769
rect 1209 707 1255 719
rect 1209 -769 1215 707
rect 1249 -769 1255 707
rect 1209 -781 1255 -769
rect 1517 707 1563 719
rect 1517 -769 1523 707
rect 1557 -769 1563 707
rect 1517 -781 1563 -769
rect 1825 707 1871 719
rect 1825 -769 1831 707
rect 1865 -769 1871 707
rect 1825 -781 1871 -769
rect 2133 707 2179 719
rect 2133 -769 2139 707
rect 2173 -769 2179 707
rect 2133 -781 2179 -769
rect 2441 707 2487 719
rect 2441 -769 2447 707
rect 2481 -769 2487 707
rect 2441 -781 2487 -769
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
