magic
tech sky130A
magscale 1 2
timestamp 1770003941
<< pwell >>
rect -7400 9090 3200 35418
<< psubdiff >>
rect -7392 35354 3208 35390
rect -7396 34998 3208 35354
rect -7396 34992 3204 34998
rect -7398 34962 3204 34992
rect -7398 34870 3196 34962
rect -7402 34820 3196 34870
rect -7402 34602 3198 34820
rect -7402 33366 -6602 34602
rect -7398 32428 -6604 33366
rect 2398 33316 3198 34602
rect 2400 32770 3196 33316
rect -7400 30924 -6600 32428
rect 2398 31840 3202 32770
rect 2396 31302 3202 31840
rect -7398 9896 -6604 30924
rect 2396 30372 3200 31302
rect 2400 9896 3196 30372
rect -7398 9696 3196 9896
rect -7398 9632 -6202 9696
rect -7400 9298 -6202 9632
rect 1998 9632 3196 9696
rect 1998 9492 3200 9632
rect 1998 9298 3204 9492
rect -7400 9240 3204 9298
rect -7396 9100 3204 9240
<< psubdiffcont >>
rect -6202 9298 1998 9696
<< locali >>
rect -7392 35354 3208 35390
rect -7396 34998 3208 35354
rect -7396 34992 3204 34998
rect -7398 34962 3204 34992
rect -7398 34870 3196 34962
rect -7402 34820 3196 34870
rect -7402 34602 3198 34820
rect -7402 33366 -6602 34602
rect -7398 32428 -6604 33366
rect 2398 33316 3198 34602
rect 2400 32770 3196 33316
rect -7400 30924 -6600 32428
rect 2398 31840 3202 32770
rect 2396 31302 3202 31840
rect -7398 9898 -6604 30924
rect 2396 30372 3200 31302
rect -2934 17684 -2362 17696
rect -2934 17676 -2506 17684
rect -2386 17676 -2362 17684
rect -2934 17266 -2362 17676
rect 2400 9898 3196 30372
rect -7402 9754 3198 9898
rect -7402 9252 -6252 9754
rect 2048 9632 3198 9754
rect 2048 9492 3200 9632
rect 2048 9252 3204 9492
rect -7402 9100 3204 9252
rect -7402 8298 3198 9100
<< viali >>
rect -6252 9696 2048 9754
rect -6252 9298 -6202 9696
rect -6202 9298 1998 9696
rect 1998 9298 2048 9696
rect -6252 9252 2048 9298
<< metal1 >>
rect -6248 36200 -5684 36254
rect -6248 35906 -6168 36200
rect -5754 35906 -5684 36200
rect -6248 35854 -5684 35906
rect 1466 36102 2036 36188
rect 1466 35750 1546 36102
rect 1940 35750 2036 36102
rect 1466 35658 2036 35750
rect -6242 34148 -5674 34232
rect -6242 33900 -6150 34148
rect -5750 33900 -5674 34148
rect -6242 33802 -5674 33900
rect -5148 34148 -4580 34236
rect -5148 33900 -5050 34148
rect -4650 33900 -4580 34148
rect -5148 33806 -4580 33900
rect -4042 34148 -3474 34234
rect -4042 33900 -3954 34148
rect -3554 33900 -3474 34148
rect -4042 33804 -3474 33900
rect -2940 34154 -2372 34238
rect -2940 33906 -2848 34154
rect -2448 33906 -2372 34154
rect -2940 33808 -2372 33906
rect -1838 34148 -1270 34234
rect -1838 33900 -1752 34148
rect -1352 33900 -1270 34148
rect -1838 33804 -1270 33900
rect -738 34148 -170 34232
rect -738 33900 -650 34148
rect -250 33900 -170 34148
rect -738 33802 -170 33900
rect 362 34150 930 34230
rect 362 33902 452 34150
rect 852 33902 930 34150
rect 362 33800 930 33902
rect 1464 34152 2032 34230
rect 1464 33904 1548 34152
rect 1948 33904 2032 34152
rect 1464 33800 2032 33904
rect -6240 31596 -5672 31700
rect -6240 31348 -6152 31596
rect -5752 31348 -5672 31596
rect -6240 31270 -5672 31348
rect -5144 31596 -4576 31706
rect -5144 31348 -5050 31596
rect -4650 31348 -4576 31596
rect -5144 31276 -4576 31348
rect -4044 31600 -3476 31706
rect -4044 31352 -3952 31600
rect -3552 31352 -3476 31600
rect -4044 31276 -3476 31352
rect -2942 31598 -2374 31706
rect -2942 31350 -2854 31598
rect -2454 31350 -2374 31598
rect -2942 31276 -2374 31350
rect -1836 31598 -1268 31694
rect -1836 31350 -1752 31598
rect -1352 31350 -1268 31598
rect -1836 31264 -1268 31350
rect -740 31596 -172 31698
rect -740 31348 -650 31596
rect -250 31348 -172 31596
rect -740 31268 -172 31348
rect 360 31598 928 31698
rect 360 31350 448 31598
rect 848 31350 928 31598
rect 360 31268 928 31350
rect 1464 31596 2032 31700
rect 1464 31348 1548 31596
rect 1948 31348 2032 31596
rect 1464 31270 2032 31348
rect -6236 30650 -5664 30728
rect -6236 30398 -6152 30650
rect -5748 30398 -5664 30650
rect -6236 30298 -5664 30398
rect -5118 30312 -3490 30706
rect -2942 30648 -2374 30740
rect -2942 30400 -2848 30648
rect -2448 30400 -2374 30648
rect -2942 30310 -2374 30400
rect -1844 30650 -1276 30746
rect -1844 30402 -1752 30650
rect -1352 30402 -1276 30650
rect -1844 30316 -1276 30402
rect -718 30318 910 30712
rect 1466 30652 2038 30732
rect 1466 30400 1548 30652
rect 1948 30400 2038 30652
rect 1466 30296 2038 30400
rect -6220 26814 -5682 28180
rect -5114 26814 -4576 28180
rect -4016 26814 -3478 28180
rect -2946 28100 -2378 28208
rect -2946 27852 -2850 28100
rect -2450 27852 -2378 28100
rect -2946 27778 -2378 27852
rect -1844 28100 -1276 28216
rect -1844 27852 -1754 28100
rect -1354 27852 -1276 28100
rect -1844 27786 -1276 27852
rect -2912 26814 -1284 27208
rect -720 26814 -182 28180
rect 380 26814 918 28180
rect 1484 26812 2022 28178
rect -6220 23314 -5682 24680
rect -5116 23314 -4578 24680
rect -4016 23310 -3478 24676
rect -2914 23326 -2388 24676
rect -1840 23646 -1272 23740
rect -1840 23398 -1752 23646
rect -1352 23398 -1272 23646
rect -1840 23310 -1272 23398
rect -720 23316 -182 24682
rect 380 23312 918 24678
rect 1484 23312 2022 24678
rect -6216 19814 -5678 21180
rect -5116 19812 -4578 21178
rect -4012 19810 -3474 21176
rect -2914 19818 -2388 21168
rect -1836 21126 -1268 21208
rect -1836 20878 -1752 21126
rect -1352 20878 -1268 21126
rect -1836 20778 -1268 20878
rect -722 19812 -184 21178
rect 384 19814 922 21180
rect 1484 19814 2022 21180
rect -2934 17684 -2362 17696
rect -6216 16314 -5678 17680
rect -5114 16314 -4576 17680
rect -4018 16312 -3480 17678
rect -2934 17676 -2506 17684
rect -2386 17676 -2362 17684
rect -2934 17600 -2362 17676
rect -2934 17350 -2850 17600
rect -2448 17350 -2362 17600
rect -2934 17266 -2362 17350
rect -2938 16652 -2370 16724
rect -2938 16404 -2850 16652
rect -2450 16404 -2370 16652
rect -2938 16294 -2370 16404
rect -1840 16650 -1272 16740
rect -1840 16402 -1752 16650
rect -1352 16402 -1272 16650
rect -1840 16310 -1272 16402
rect -720 16314 -182 17680
rect 380 16316 918 17682
rect 1488 16312 2026 17678
rect -6216 13784 -4588 14178
rect -2942 14100 -2374 14188
rect -2942 13852 -2854 14100
rect -2454 13852 -2374 14100
rect -2942 13758 -2374 13852
rect -1840 14102 -1272 14200
rect -1840 13854 -1752 14102
rect -1352 13854 -1272 14102
rect -1840 13770 -1272 13854
rect 386 13788 2014 14182
rect -6242 13146 -5674 13240
rect -4048 13232 -3480 13238
rect -1838 13236 -1270 13238
rect -6242 12898 -6154 13146
rect -5754 12898 -5674 13146
rect -6242 12810 -5674 12898
rect -6240 12804 -5674 12810
rect -5138 13154 -4572 13232
rect -5138 12906 -5056 13154
rect -4656 12906 -4572 13154
rect -5138 12802 -4572 12906
rect -4048 13148 -3476 13232
rect -4048 12900 -3952 13148
rect -3552 12900 -3476 13148
rect -4048 12808 -3476 12900
rect -4044 12804 -3476 12808
rect -2930 13148 -2360 13232
rect -2930 12900 -2850 13148
rect -2450 12900 -2360 13148
rect -2930 12804 -2360 12900
rect -1838 13144 -1268 13236
rect -1838 12896 -1752 13144
rect -1352 12896 -1268 13144
rect -1838 12808 -1268 12896
rect -1834 12804 -1268 12808
rect -740 13150 -170 13232
rect -740 12902 -650 13150
rect -250 12902 -170 13150
rect -740 12804 -170 12902
rect -4044 12800 -3478 12804
rect -2928 12802 -2360 12804
rect -738 12802 -170 12804
rect 358 13144 932 13232
rect 358 12896 450 13144
rect 850 12896 932 13144
rect 358 12804 932 12896
rect 1460 13150 2030 13232
rect 1460 12902 1552 13150
rect 1952 12902 2030 13150
rect 1460 12804 2030 12902
rect 358 12802 926 12804
rect 1462 12802 2030 12804
rect -6242 10698 -5674 10704
rect -6244 10616 -5674 10698
rect -6244 10368 -6152 10616
rect -5752 10368 -5674 10616
rect -6244 10274 -5674 10368
rect -5142 10702 -4574 10704
rect -5142 10624 -4572 10702
rect -5142 10376 -5050 10624
rect -4650 10376 -4572 10624
rect -5142 10274 -4572 10376
rect -4046 10618 -3478 10704
rect -4046 10370 -3950 10618
rect -3550 10370 -3478 10618
rect -4046 10274 -3478 10370
rect -2930 10620 -2362 10704
rect -2930 10372 -2848 10620
rect -2448 10372 -2362 10620
rect -2930 10274 -2362 10372
rect -1842 10702 -1274 10708
rect -1842 10630 -1268 10702
rect -1842 10382 -1750 10630
rect -1350 10382 -1268 10630
rect -1842 10278 -1268 10382
rect -1834 10274 -1268 10278
rect -742 10622 -174 10700
rect -742 10374 -650 10622
rect -250 10374 -174 10622
rect -6244 10270 -5678 10274
rect -2928 10270 -2362 10274
rect -742 10270 -174 10374
rect 358 10698 926 10700
rect 358 10624 930 10698
rect 358 10376 448 10624
rect 848 10376 930 10624
rect 358 10270 930 10376
rect 1462 10618 2030 10704
rect 1462 10370 1550 10618
rect 1950 10370 2030 10618
rect 1462 10274 2030 10370
rect 1462 10266 2028 10274
rect -7398 9898 3196 9900
rect -7402 9754 3198 9898
rect -7402 9252 -6252 9754
rect 2048 9752 3198 9754
rect -7402 9250 -6250 9252
rect 2050 9250 3198 9752
rect -7402 8298 3198 9250
<< via1 >>
rect -6168 35906 -5754 36200
rect 1546 35750 1940 36102
rect -6150 33900 -5750 34148
rect -5050 33900 -4650 34148
rect -3954 33900 -3554 34148
rect -2848 33906 -2448 34154
rect -1752 33900 -1352 34148
rect -650 33900 -250 34148
rect 452 33902 852 34150
rect 1548 33904 1948 34152
rect -6152 31348 -5752 31596
rect -5050 31348 -4650 31596
rect -3952 31352 -3552 31600
rect -2854 31350 -2454 31598
rect -1752 31350 -1352 31598
rect -650 31348 -250 31596
rect 448 31350 848 31598
rect 1548 31348 1948 31596
rect -6152 30398 -5748 30650
rect -2848 30400 -2448 30648
rect -1752 30402 -1352 30650
rect 1548 30400 1948 30652
rect -2850 27852 -2450 28100
rect -1754 27852 -1354 28100
rect -1750 24358 -1352 24600
rect -1752 23398 -1352 23646
rect -1752 20878 -1352 21126
rect -1748 19900 -1350 20142
rect -2850 17350 -2448 17600
rect -1750 17356 -1352 17606
rect -2850 16404 -2450 16652
rect -1752 16402 -1352 16650
rect -3952 13852 -3550 14102
rect -2854 13852 -2454 14100
rect -1752 13854 -1352 14102
rect -648 13850 -250 14100
rect -6154 12898 -5754 13146
rect -5056 12906 -4656 13154
rect -3952 12900 -3552 13148
rect -2850 12900 -2450 13148
rect -1752 12896 -1352 13144
rect -650 12902 -250 13150
rect 450 12896 850 13144
rect 1552 12902 1952 13150
rect -6152 10368 -5752 10616
rect -5050 10376 -4650 10624
rect -3950 10370 -3550 10618
rect -2848 10372 -2448 10620
rect -1750 10382 -1350 10630
rect -650 10374 -250 10622
rect 448 10376 848 10624
rect 1550 10370 1950 10618
rect -6252 9252 2048 9754
rect 2048 9252 2050 9752
rect -6250 9250 2050 9252
<< metal2 >>
rect -6248 36200 -5684 36254
rect -6248 35906 -6168 36200
rect -5754 35906 -5684 36200
rect -6248 35854 -5684 35906
rect 1466 36102 2036 36188
rect 1466 35750 1546 36102
rect 1940 35750 2036 36102
rect 1466 35658 2036 35750
rect -6242 34148 -5674 34232
rect -6242 33900 -6150 34148
rect -5750 33900 -5674 34148
rect -6242 33802 -5674 33900
rect -5148 34148 -4580 34236
rect -5148 33900 -5050 34148
rect -4650 33900 -4580 34148
rect -5148 33806 -4580 33900
rect -4042 34148 -3474 34234
rect -4042 33900 -3954 34148
rect -3554 33900 -3474 34148
rect -4042 33804 -3474 33900
rect -2940 34154 -2372 34238
rect -2940 33906 -2848 34154
rect -2448 33906 -2372 34154
rect -2940 33808 -2372 33906
rect -1838 34148 -1270 34234
rect -1838 33900 -1752 34148
rect -1352 33900 -1270 34148
rect -1838 33804 -1270 33900
rect -738 34148 -170 34232
rect -738 33900 -650 34148
rect -250 33900 -170 34148
rect -738 33802 -170 33900
rect 362 34150 930 34230
rect 362 33902 452 34150
rect 852 33902 930 34150
rect 362 33800 930 33902
rect 1464 34152 2032 34230
rect 1464 33904 1548 34152
rect 1948 33904 2032 34152
rect 1464 33800 2032 33904
rect -6240 31596 -5672 31700
rect -6240 31348 -6152 31596
rect -5752 31348 -5672 31596
rect -6240 31270 -5672 31348
rect -5144 31596 -4576 31706
rect -5144 31348 -5050 31596
rect -4650 31348 -4576 31596
rect -5144 31276 -4576 31348
rect -4044 31600 -3476 31706
rect -4044 31352 -3952 31600
rect -3552 31352 -3476 31600
rect -4044 31276 -3476 31352
rect -2942 31598 -2374 31706
rect -2942 31350 -2854 31598
rect -2454 31350 -2374 31598
rect -2942 31276 -2374 31350
rect -1836 31598 -1268 31694
rect -1836 31350 -1752 31598
rect -1352 31350 -1268 31598
rect -1836 31264 -1268 31350
rect -740 31596 -172 31698
rect -740 31348 -650 31596
rect -250 31348 -172 31596
rect -740 31268 -172 31348
rect 360 31598 928 31698
rect 360 31350 448 31598
rect 848 31350 928 31598
rect 360 31268 928 31350
rect 1464 31596 2032 31700
rect 1464 31348 1548 31596
rect 1948 31348 2032 31596
rect 1464 31270 2032 31348
rect -6236 30650 -5664 30728
rect -6236 30398 -6152 30650
rect -5748 30398 -5664 30650
rect -6236 30298 -5664 30398
rect -2942 30648 -2374 30740
rect -2942 30400 -2848 30648
rect -2448 30400 -2374 30648
rect -2942 30310 -2374 30400
rect -1844 30650 -1276 30746
rect -1844 30402 -1752 30650
rect -1352 30402 -1276 30650
rect -1844 30316 -1276 30402
rect 1466 30652 2038 30732
rect 1466 30400 1548 30652
rect 1948 30400 2038 30652
rect 1466 30296 2038 30400
rect -2946 28100 -2378 28208
rect -2946 27852 -2850 28100
rect -2450 27852 -2378 28100
rect -2946 27778 -2378 27852
rect -1844 28100 -1276 28216
rect -1844 27852 -1754 28100
rect -1354 27852 -1276 28100
rect -1844 27786 -1276 27852
rect -1836 24600 -166 24704
rect -1836 24358 -1750 24600
rect -1352 24358 -166 24600
rect -1836 24272 -166 24358
rect -1840 23646 -1272 23740
rect -1840 23398 -1752 23646
rect -1352 23398 -1272 23646
rect -1840 23310 -1272 23398
rect -1836 21126 -1268 21208
rect -1836 20878 -1752 21126
rect -1352 20878 -1268 21126
rect -1836 20778 -1268 20878
rect -734 20230 -166 24272
rect -1834 20142 -164 20230
rect -1834 19900 -1748 20142
rect -1350 19900 -164 20142
rect -1834 19798 -164 19900
rect -4036 17600 -2366 17700
rect -4036 17350 -2850 17600
rect -2448 17350 -2366 17600
rect -4036 17272 -2366 17350
rect -1834 17606 -164 17700
rect -1834 17356 -1750 17606
rect -1352 17356 -164 17606
rect -1834 17274 -164 17356
rect -4034 14102 -3466 17272
rect -2938 16652 -2370 16724
rect -2938 16404 -2850 16652
rect -2450 16404 -2370 16652
rect -2938 16294 -2370 16404
rect -1840 16650 -1272 16740
rect -1840 16402 -1752 16650
rect -1352 16402 -1272 16650
rect -1840 16310 -1272 16402
rect -4034 13852 -3952 14102
rect -3550 13852 -3466 14102
rect -4034 13770 -3466 13852
rect -2942 14100 -2374 14188
rect -2942 13852 -2854 14100
rect -2454 13852 -2374 14100
rect -2942 13758 -2374 13852
rect -1840 14102 -1272 14200
rect -1840 13854 -1752 14102
rect -1352 13854 -1272 14102
rect -1840 13770 -1272 13854
rect -734 14100 -166 17274
rect -734 13850 -648 14100
rect -250 13850 -166 14100
rect -734 13766 -166 13850
rect -6242 13146 -5674 13240
rect -6242 12898 -6154 13146
rect -5754 12898 -5674 13146
rect -6242 12810 -5674 12898
rect -6240 12804 -5674 12810
rect -5142 13232 -4574 13236
rect -4048 13232 -3480 13238
rect -1838 13236 -1270 13238
rect -5142 13154 -4572 13232
rect -5142 12906 -5056 13154
rect -4656 12906 -4572 13154
rect -5142 12806 -4572 12906
rect -4048 13148 -3476 13232
rect -4048 12900 -3952 13148
rect -3552 12900 -3476 13148
rect -4048 12808 -3476 12900
rect -5138 12802 -4572 12806
rect -4044 12804 -3476 12808
rect -2930 13148 -2360 13232
rect -2930 12900 -2850 13148
rect -2450 12900 -2360 13148
rect -2930 12804 -2360 12900
rect -1838 13144 -1268 13236
rect -1838 12896 -1752 13144
rect -1352 12896 -1268 13144
rect -1838 12808 -1268 12896
rect -1834 12804 -1268 12808
rect -740 13150 -170 13232
rect -740 12902 -650 13150
rect -250 12902 -170 13150
rect -740 12804 -170 12902
rect -4044 12800 -3478 12804
rect -2928 12802 -2360 12804
rect -738 12802 -170 12804
rect 358 13144 932 13232
rect 358 12896 450 13144
rect 850 12896 932 13144
rect 358 12804 932 12896
rect 1460 13150 2030 13232
rect 1460 12902 1552 13150
rect 1952 12902 2030 13150
rect 1460 12804 2030 12902
rect 358 12802 926 12804
rect 1462 12802 2030 12804
rect -6242 10698 -5674 10704
rect -6244 10616 -5674 10698
rect -6244 10368 -6152 10616
rect -5752 10368 -5674 10616
rect -6244 10274 -5674 10368
rect -5142 10702 -4574 10704
rect -5142 10624 -4572 10702
rect -5142 10376 -5050 10624
rect -4650 10376 -4572 10624
rect -5142 10274 -4572 10376
rect -4046 10618 -3478 10704
rect -4046 10370 -3950 10618
rect -3550 10370 -3478 10618
rect -4046 10274 -3478 10370
rect -2930 10620 -2362 10704
rect -2930 10372 -2848 10620
rect -2448 10372 -2362 10620
rect -2930 10274 -2362 10372
rect -1842 10702 -1274 10708
rect -1842 10630 -1268 10702
rect -1842 10382 -1750 10630
rect -1350 10382 -1268 10630
rect -1842 10278 -1268 10382
rect -1834 10274 -1268 10278
rect -742 10622 -174 10700
rect -742 10374 -650 10622
rect -250 10374 -174 10622
rect -6244 10270 -5678 10274
rect -2928 10270 -2362 10274
rect -742 10270 -174 10374
rect 358 10698 926 10700
rect 358 10624 930 10698
rect 358 10376 448 10624
rect 848 10376 930 10624
rect 358 10270 930 10376
rect 1462 10618 2030 10704
rect 1462 10370 1550 10618
rect 1950 10370 2030 10618
rect 1462 10274 2030 10370
rect 1462 10266 2028 10274
rect -7398 9754 3196 9900
rect -7398 9252 -6252 9754
rect 2048 9752 3196 9754
rect -7398 9250 -6250 9252
rect 2050 9250 3196 9752
rect -7398 8298 3196 9250
<< via2 >>
rect -6168 35906 -5754 36200
rect 1546 35750 1940 36102
rect -6150 33900 -5750 34148
rect -5050 33900 -4650 34148
rect -3954 33900 -3554 34148
rect -2848 33906 -2448 34154
rect -1752 33900 -1352 34148
rect -650 33900 -250 34148
rect 452 33902 852 34150
rect 1548 33904 1948 34152
rect -6152 31348 -5752 31596
rect -5050 31348 -4650 31596
rect -3952 31352 -3552 31600
rect -2854 31350 -2454 31598
rect -1752 31350 -1352 31598
rect -650 31348 -250 31596
rect 448 31350 848 31598
rect 1548 31348 1948 31596
rect -6152 30398 -5748 30650
rect -2848 30400 -2448 30648
rect -1752 30402 -1352 30650
rect 1548 30400 1948 30652
rect -2850 27852 -2450 28100
rect -1754 27852 -1354 28100
rect -1752 23398 -1352 23646
rect -1752 20878 -1352 21126
rect -2850 16404 -2450 16652
rect -1752 16402 -1352 16650
rect -2854 13852 -2454 14100
rect -1752 13854 -1352 14102
rect -6154 12898 -5754 13146
rect -5056 12906 -4656 13154
rect -3952 12900 -3552 13148
rect -2850 12900 -2450 13148
rect -1752 12896 -1352 13144
rect -650 12902 -250 13150
rect 450 12896 850 13144
rect 1552 12902 1952 13150
rect -6152 10368 -5752 10616
rect -5050 10376 -4650 10624
rect -3950 10370 -3550 10618
rect -2848 10372 -2448 10620
rect -1750 10382 -1350 10630
rect -650 10374 -250 10622
rect 448 10376 848 10624
rect 1550 10370 1950 10618
rect -6252 9752 2048 9754
rect -6252 9252 2050 9752
rect -6250 9250 2050 9252
<< metal3 >>
rect -6248 36200 -5684 36254
rect -6248 35906 -6168 36200
rect -5754 35906 -5684 36200
rect -6248 35854 -5684 35906
rect 1466 36102 2036 36188
rect 1466 35750 1546 36102
rect 1940 35750 2036 36102
rect 1466 35658 2036 35750
rect -2940 34236 -2372 34238
rect -6242 34148 -5674 34232
rect -6242 33900 -6150 34148
rect -5750 33900 -5674 34148
rect -6242 33802 -5674 33900
rect -5148 34148 -4580 34236
rect -5148 33900 -5050 34148
rect -4650 33900 -4580 34148
rect -5148 33806 -4580 33900
rect -4042 34148 -3474 34234
rect -2940 34232 -2358 34236
rect -4042 33900 -3954 34148
rect -3554 33900 -3474 34148
rect -4042 33804 -3474 33900
rect -2940 34154 -2372 34232
rect -2940 33906 -2848 34154
rect -2448 33906 -2372 34154
rect -2940 33808 -2372 33906
rect -1838 34148 -1270 34234
rect -1838 33900 -1752 34148
rect -1352 33900 -1270 34148
rect -1838 33804 -1270 33900
rect -738 34148 -170 34232
rect -738 33900 -650 34148
rect -250 33900 -170 34148
rect -738 33802 -170 33900
rect 362 34150 930 34230
rect 362 33902 452 34150
rect 852 33902 930 34150
rect 362 33800 930 33902
rect 1464 34152 2032 34230
rect 1464 33904 1548 34152
rect 1948 33904 2032 34152
rect 1464 33800 2032 33904
rect -2940 33394 -2358 33798
rect -1836 33394 -1254 33798
rect -2940 31890 -2354 33394
rect -1840 31890 -1254 33394
rect -2940 31706 -2358 31890
rect -5144 31704 -4576 31706
rect -4044 31704 -3476 31706
rect -2942 31704 -2358 31706
rect -1836 31704 -1254 31890
rect -6246 31700 2028 31704
rect -6246 31600 2032 31700
rect -6246 31596 -3952 31600
rect -6246 31348 -6152 31596
rect -5752 31348 -5050 31596
rect -4650 31352 -3952 31596
rect -3552 31598 2032 31600
rect -3552 31352 -2854 31598
rect -4650 31350 -2854 31352
rect -2454 31350 -1752 31598
rect -1352 31596 448 31598
rect -1352 31350 -650 31596
rect -4650 31348 -650 31350
rect -250 31350 448 31596
rect 848 31596 2032 31598
rect 848 31350 1548 31596
rect -250 31348 1548 31350
rect 1948 31348 2032 31596
rect -6246 31270 2032 31348
rect -2940 30970 -2358 31270
rect -1836 30970 -1254 31270
rect -740 31268 -172 31270
rect 360 31268 928 31270
rect -2940 30740 -2354 30970
rect -1840 30746 -1254 30970
rect -6236 30650 -5664 30728
rect -6236 30398 -6152 30650
rect -5748 30398 -5664 30650
rect -6236 30298 -5664 30398
rect -2942 30648 -2354 30740
rect -2942 30400 -2848 30648
rect -2448 30400 -2354 30648
rect -2942 30310 -2354 30400
rect -1844 30650 -1254 30746
rect -1844 30402 -1752 30650
rect -1352 30402 -1254 30650
rect -1844 30316 -1254 30402
rect -2940 28208 -2354 30310
rect -1840 28216 -1254 30316
rect 1466 30652 2038 30732
rect 1466 30400 1548 30652
rect 1948 30400 2038 30652
rect 1466 30296 2038 30400
rect -2946 28100 -2354 28208
rect -2946 27852 -2850 28100
rect -2450 27852 -2354 28100
rect -2946 27778 -2354 27852
rect -1844 28100 -1254 28216
rect -1844 27852 -1754 28100
rect -1354 27852 -1254 28100
rect -1844 27786 -1254 27852
rect -2940 16652 -2354 27778
rect -2940 16404 -2850 16652
rect -2450 16404 -2354 16652
rect -2940 14188 -2354 16404
rect -2942 14100 -2354 14188
rect -2942 13852 -2854 14100
rect -2454 13852 -2354 14100
rect -2942 13758 -2354 13852
rect -6242 13236 -5674 13240
rect -4048 13236 -3480 13238
rect -2940 13236 -2354 13758
rect -1840 23646 -1254 27786
rect -1840 23398 -1752 23646
rect -1352 23398 -1254 23646
rect -1840 21126 -1254 23398
rect -1840 20878 -1752 21126
rect -1352 20878 -1254 21126
rect -1840 16650 -1254 20878
rect -1840 16402 -1752 16650
rect -1352 16402 -1254 16650
rect -1840 14102 -1254 16402
rect -1840 13854 -1752 14102
rect -1352 13854 -1254 14102
rect -1840 13236 -1254 13854
rect -6242 13154 2034 13236
rect -6242 13146 -5056 13154
rect -6242 12898 -6154 13146
rect -5754 12906 -5056 13146
rect -4656 13150 2034 13154
rect -4656 13148 -650 13150
rect -4656 12906 -3952 13148
rect -5754 12900 -3952 12906
rect -3552 12900 -2850 13148
rect -2450 13144 -650 13148
rect -2450 12900 -1752 13144
rect -5754 12898 -1752 12900
rect -6242 12896 -1752 12898
rect -1352 12902 -650 13144
rect -250 13144 1552 13150
rect -250 12902 450 13144
rect -1352 12896 450 12902
rect 850 12902 1552 13144
rect 1952 12902 2034 13150
rect 850 12896 2034 12902
rect -6242 12810 2034 12896
rect -6240 12802 2034 12810
rect -4044 12800 -3478 12802
rect -2940 10710 -2354 12802
rect -1840 10710 -1254 12802
rect -6244 10704 2030 10710
rect -6244 10630 2036 10704
rect -6244 10624 -1750 10630
rect -6244 10616 -5050 10624
rect -6244 10368 -6152 10616
rect -5752 10376 -5050 10616
rect -4650 10620 -1750 10624
rect -4650 10618 -2848 10620
rect -4650 10376 -3950 10618
rect -5752 10370 -3950 10376
rect -3550 10372 -2848 10618
rect -2448 10382 -1750 10620
rect -1350 10624 2036 10630
rect -1350 10622 448 10624
rect -1350 10382 -650 10622
rect -2448 10374 -650 10382
rect -250 10376 448 10622
rect 848 10618 2036 10624
rect 848 10376 1550 10618
rect -250 10374 1550 10376
rect -2448 10372 1550 10374
rect -3550 10370 1550 10372
rect 1950 10492 2036 10618
rect 1950 10370 2038 10492
rect -5752 10368 2038 10370
rect -6244 10270 2038 10368
rect -6242 10054 2038 10270
rect -6240 9900 2036 10054
rect -7398 9754 3196 9900
rect -7398 9252 -6252 9754
rect 2048 9752 3196 9754
rect -7398 9250 -6250 9252
rect 2050 9250 3196 9752
rect -7398 8298 3196 9250
<< rmetal3 >>
rect -5674 33806 -5148 34232
rect -4580 33806 -4042 34232
rect -5674 33804 -4042 33806
rect -3474 33808 -2940 34232
rect -2372 33808 -1838 34232
rect -3474 33804 -1838 33808
rect -1270 33804 -738 34232
rect -170 34230 2034 34232
rect -5674 33802 -738 33804
rect -170 33802 362 34230
rect -6240 33800 362 33802
rect 930 33800 1464 34230
rect 2032 33800 2034 34230
rect -6240 33798 2034 33800
<< via3 >>
rect -6168 35906 -5754 36200
rect 1546 35750 1940 36102
rect -6152 30398 -5748 30650
rect 1548 30400 1948 30652
<< metal4 >>
rect -6248 36200 -5684 36254
rect -6248 35906 -6168 36200
rect -5754 35906 -5684 36200
rect 1466 36148 2036 36188
rect -6248 35778 -5684 35906
rect 1464 36102 2036 36148
rect -6248 35614 -5674 35778
rect 1464 35750 1546 36102
rect 1940 35750 2036 36102
rect 1464 35618 2036 35750
rect -6244 34226 -5674 35614
rect -6246 32822 -5674 34226
rect -6246 31852 -5676 32822
rect 1466 31858 2036 35618
rect -6246 30650 -5662 31852
rect -6246 30398 -6152 30650
rect -5748 30398 -5662 30650
rect -6246 30298 -5662 30398
rect 1460 30652 2044 31858
rect 1460 30400 1548 30652
rect 1948 30400 2044 30652
rect 1460 30304 2044 30400
rect 1466 30296 2038 30304
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_0
timestamp 1769960253
transform 1 0 -5957 0 1 32749
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_1
timestamp 1769960253
transform 1 0 -4861 0 1 32753
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_2
timestamp 1769960253
transform 1 0 -3757 0 1 32753
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_3
timestamp 1769960253
transform 1 0 -2653 0 1 32755
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_4
timestamp 1769960253
transform 1 0 -1551 0 1 32751
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_5
timestamp 1769960253
transform 1 0 -451 0 1 32749
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_6
timestamp 1769960253
transform 1 0 647 0 1 32751
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_7
timestamp 1769960253
transform 1 0 1751 0 1 32749
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_8
timestamp 1769960253
transform 1 0 -2655 0 1 29257
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_9
timestamp 1769960253
transform 1 0 -1559 0 1 29265
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_10
timestamp 1769960253
transform 1 0 -1551 0 1 22253
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_11
timestamp 1769960253
transform 1 0 -2653 0 1 15235
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_12
timestamp 1769960253
transform 1 0 -1553 0 1 15251
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_13
timestamp 1769960253
transform 1 0 -5955 0 1 11753
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_14
timestamp 1769960253
transform 1 0 -4855 0 1 11753
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_15
timestamp 1769960253
transform 1 0 -3761 0 1 11753
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_16
timestamp 1769960253
transform 1 0 -2643 0 1 11751
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_17
timestamp 1769960253
transform 1 0 -1551 0 1 11753
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_18
timestamp 1769960253
transform 1 0 -455 0 1 11749
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_19
timestamp 1769960253
transform 1 0 647 0 1 11749
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  sky130_fd_pr__res_xhigh_po_2p85_789E74_20
timestamp 1769960253
transform 1 0 1747 0 1 11751
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR1
timestamp 1769960253
transform 1 0 -5949 0 1 29247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR2
timestamp 1769960253
transform 1 0 -5949 0 1 25747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR3
timestamp 1769960253
transform 1 0 -5949 0 1 22247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR4
timestamp 1769960253
transform 1 0 -5949 0 1 18747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR5
timestamp 1769960253
transform 1 0 -5949 0 1 15247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR6
timestamp 1769960253
transform 1 0 -4849 0 1 15247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR7
timestamp 1769960253
transform 1 0 -4849 0 1 18747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR8
timestamp 1769960253
transform 1 0 -4849 0 1 22247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR9
timestamp 1769960253
transform 1 0 -4849 0 1 25747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR10
timestamp 1769960253
transform 1 0 -4849 0 1 29247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR11
timestamp 1769960253
transform 1 0 -3749 0 1 15247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR12
timestamp 1769960253
transform 1 0 -3749 0 1 18747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR13
timestamp 1769960253
transform 1 0 -3749 0 1 22247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR14
timestamp 1769960253
transform 1 0 -3749 0 1 25747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR15
timestamp 1769960253
transform 1 0 -3749 0 1 29247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR16
timestamp 1769960253
transform 1 0 -2649 0 1 18747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR17
timestamp 1769960253
transform 1 0 -2649 0 1 22247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR18
timestamp 1769960253
transform 1 0 -2649 0 1 25747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR19
timestamp 1769960253
transform 1 0 -1549 0 1 25747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR20
timestamp 1769960253
transform 1 0 -1549 0 1 18747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR21
timestamp 1769960253
transform 1 0 -449 0 1 15247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR22
timestamp 1769960253
transform 1 0 -449 0 1 18747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR23
timestamp 1769960253
transform 1 0 -449 0 1 22247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR24
timestamp 1769960253
transform 1 0 -449 0 1 25747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR25
timestamp 1769960253
transform 1 0 -449 0 1 29247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR26
timestamp 1769960253
transform 1 0 651 0 1 29247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR27
timestamp 1769960253
transform 1 0 651 0 1 25747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR28
timestamp 1769960253
transform 1 0 651 0 1 22247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR29
timestamp 1769960253
transform 1 0 651 0 1 18747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR30
timestamp 1769960253
transform 1 0 651 0 1 15247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR31
timestamp 1769960253
transform 1 0 1751 0 1 15247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR32
timestamp 1769960253
transform 1 0 1751 0 1 18747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR33
timestamp 1769960253
transform 1 0 1751 0 1 22247
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR34
timestamp 1769960253
transform 1 0 1751 0 1 25747
box -451 -1647 451 1647
use sky130_fd_pr__res_xhigh_po_2p85_789E74  XR35
timestamp 1769960253
transform 1 0 1751 0 1 29247
box -451 -1647 451 1647
<< labels >>
flabel metal1 -2232 8568 -2032 8768 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel via1 -6048 35946 -5848 36146 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel via1 1644 35852 1844 36052 0 FreeSans 256 0 0 0 B
port 2 nsew
<< end >>
