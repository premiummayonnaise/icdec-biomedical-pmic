magic
tech sky130A
magscale 1 2
timestamp 1769999431
<< error_p >>
rect -2867 1038 2867 1042
rect -2867 -970 -2837 1038
rect -2801 972 2801 976
rect -2801 -904 -2771 972
rect 2771 -904 2801 972
rect 2837 -970 2867 1038
<< nwell >>
rect -2837 -1004 2837 1038
<< mvpmos >>
rect -2743 -904 -2493 976
rect -2435 -904 -2185 976
rect -2127 -904 -1877 976
rect -1819 -904 -1569 976
rect -1511 -904 -1261 976
rect -1203 -904 -953 976
rect -895 -904 -645 976
rect -587 -904 -337 976
rect -279 -904 -29 976
rect 29 -904 279 976
rect 337 -904 587 976
rect 645 -904 895 976
rect 953 -904 1203 976
rect 1261 -904 1511 976
rect 1569 -904 1819 976
rect 1877 -904 2127 976
rect 2185 -904 2435 976
rect 2493 -904 2743 976
<< mvpdiff >>
rect -2801 964 -2743 976
rect -2801 -892 -2789 964
rect -2755 -892 -2743 964
rect -2801 -904 -2743 -892
rect -2493 964 -2435 976
rect -2493 -892 -2481 964
rect -2447 -892 -2435 964
rect -2493 -904 -2435 -892
rect -2185 964 -2127 976
rect -2185 -892 -2173 964
rect -2139 -892 -2127 964
rect -2185 -904 -2127 -892
rect -1877 964 -1819 976
rect -1877 -892 -1865 964
rect -1831 -892 -1819 964
rect -1877 -904 -1819 -892
rect -1569 964 -1511 976
rect -1569 -892 -1557 964
rect -1523 -892 -1511 964
rect -1569 -904 -1511 -892
rect -1261 964 -1203 976
rect -1261 -892 -1249 964
rect -1215 -892 -1203 964
rect -1261 -904 -1203 -892
rect -953 964 -895 976
rect -953 -892 -941 964
rect -907 -892 -895 964
rect -953 -904 -895 -892
rect -645 964 -587 976
rect -645 -892 -633 964
rect -599 -892 -587 964
rect -645 -904 -587 -892
rect -337 964 -279 976
rect -337 -892 -325 964
rect -291 -892 -279 964
rect -337 -904 -279 -892
rect -29 964 29 976
rect -29 -892 -17 964
rect 17 -892 29 964
rect -29 -904 29 -892
rect 279 964 337 976
rect 279 -892 291 964
rect 325 -892 337 964
rect 279 -904 337 -892
rect 587 964 645 976
rect 587 -892 599 964
rect 633 -892 645 964
rect 587 -904 645 -892
rect 895 964 953 976
rect 895 -892 907 964
rect 941 -892 953 964
rect 895 -904 953 -892
rect 1203 964 1261 976
rect 1203 -892 1215 964
rect 1249 -892 1261 964
rect 1203 -904 1261 -892
rect 1511 964 1569 976
rect 1511 -892 1523 964
rect 1557 -892 1569 964
rect 1511 -904 1569 -892
rect 1819 964 1877 976
rect 1819 -892 1831 964
rect 1865 -892 1877 964
rect 1819 -904 1877 -892
rect 2127 964 2185 976
rect 2127 -892 2139 964
rect 2173 -892 2185 964
rect 2127 -904 2185 -892
rect 2435 964 2493 976
rect 2435 -892 2447 964
rect 2481 -892 2493 964
rect 2435 -904 2493 -892
rect 2743 964 2801 976
rect 2743 -892 2755 964
rect 2789 -892 2801 964
rect 2743 -904 2801 -892
<< mvpdiffc >>
rect -2789 -892 -2755 964
rect -2481 -892 -2447 964
rect -2173 -892 -2139 964
rect -1865 -892 -1831 964
rect -1557 -892 -1523 964
rect -1249 -892 -1215 964
rect -941 -892 -907 964
rect -633 -892 -599 964
rect -325 -892 -291 964
rect -17 -892 17 964
rect 291 -892 325 964
rect 599 -892 633 964
rect 907 -892 941 964
rect 1215 -892 1249 964
rect 1523 -892 1557 964
rect 1831 -892 1865 964
rect 2139 -892 2173 964
rect 2447 -892 2481 964
rect 2755 -892 2789 964
<< poly >>
rect -2743 976 -2493 1002
rect -2435 976 -2185 1002
rect -2127 976 -1877 1002
rect -1819 976 -1569 1002
rect -1511 976 -1261 1002
rect -1203 976 -953 1002
rect -895 976 -645 1002
rect -587 976 -337 1002
rect -279 976 -29 1002
rect 29 976 279 1002
rect 337 976 587 1002
rect 645 976 895 1002
rect 953 976 1203 1002
rect 1261 976 1511 1002
rect 1569 976 1819 1002
rect 1877 976 2127 1002
rect 2185 976 2435 1002
rect 2493 976 2743 1002
rect -2743 -951 -2493 -904
rect -2743 -968 -2689 -951
rect -2705 -985 -2689 -968
rect -2547 -968 -2493 -951
rect -2435 -951 -2185 -904
rect -2435 -968 -2381 -951
rect -2547 -985 -2531 -968
rect -2705 -1001 -2531 -985
rect -2397 -985 -2381 -968
rect -2239 -968 -2185 -951
rect -2127 -951 -1877 -904
rect -2127 -968 -2073 -951
rect -2239 -985 -2223 -968
rect -2397 -1001 -2223 -985
rect -2089 -985 -2073 -968
rect -1931 -968 -1877 -951
rect -1819 -951 -1569 -904
rect -1819 -968 -1765 -951
rect -1931 -985 -1915 -968
rect -2089 -1001 -1915 -985
rect -1781 -985 -1765 -968
rect -1623 -968 -1569 -951
rect -1511 -951 -1261 -904
rect -1511 -968 -1457 -951
rect -1623 -985 -1607 -968
rect -1781 -1001 -1607 -985
rect -1473 -985 -1457 -968
rect -1315 -968 -1261 -951
rect -1203 -951 -953 -904
rect -1203 -968 -1149 -951
rect -1315 -985 -1299 -968
rect -1473 -1001 -1299 -985
rect -1165 -985 -1149 -968
rect -1007 -968 -953 -951
rect -895 -951 -645 -904
rect -895 -968 -841 -951
rect -1007 -985 -991 -968
rect -1165 -1001 -991 -985
rect -857 -985 -841 -968
rect -699 -968 -645 -951
rect -587 -951 -337 -904
rect -587 -968 -533 -951
rect -699 -985 -683 -968
rect -857 -1001 -683 -985
rect -549 -985 -533 -968
rect -391 -968 -337 -951
rect -279 -951 -29 -904
rect -279 -968 -225 -951
rect -391 -985 -375 -968
rect -549 -1001 -375 -985
rect -241 -985 -225 -968
rect -83 -968 -29 -951
rect 29 -951 279 -904
rect 29 -968 83 -951
rect -83 -985 -67 -968
rect -241 -1001 -67 -985
rect 67 -985 83 -968
rect 225 -968 279 -951
rect 337 -951 587 -904
rect 337 -968 391 -951
rect 225 -985 241 -968
rect 67 -1001 241 -985
rect 375 -985 391 -968
rect 533 -968 587 -951
rect 645 -951 895 -904
rect 645 -968 699 -951
rect 533 -985 549 -968
rect 375 -1001 549 -985
rect 683 -985 699 -968
rect 841 -968 895 -951
rect 953 -951 1203 -904
rect 953 -968 1007 -951
rect 841 -985 857 -968
rect 683 -1001 857 -985
rect 991 -985 1007 -968
rect 1149 -968 1203 -951
rect 1261 -951 1511 -904
rect 1261 -968 1315 -951
rect 1149 -985 1165 -968
rect 991 -1001 1165 -985
rect 1299 -985 1315 -968
rect 1457 -968 1511 -951
rect 1569 -951 1819 -904
rect 1569 -968 1623 -951
rect 1457 -985 1473 -968
rect 1299 -1001 1473 -985
rect 1607 -985 1623 -968
rect 1765 -968 1819 -951
rect 1877 -951 2127 -904
rect 1877 -968 1931 -951
rect 1765 -985 1781 -968
rect 1607 -1001 1781 -985
rect 1915 -985 1931 -968
rect 2073 -968 2127 -951
rect 2185 -951 2435 -904
rect 2185 -968 2239 -951
rect 2073 -985 2089 -968
rect 1915 -1001 2089 -985
rect 2223 -985 2239 -968
rect 2381 -968 2435 -951
rect 2493 -951 2743 -904
rect 2493 -968 2547 -951
rect 2381 -985 2397 -968
rect 2223 -1001 2397 -985
rect 2531 -985 2547 -968
rect 2689 -968 2743 -951
rect 2689 -985 2705 -968
rect 2531 -1001 2705 -985
<< polycont >>
rect -2689 -985 -2547 -951
rect -2381 -985 -2239 -951
rect -2073 -985 -1931 -951
rect -1765 -985 -1623 -951
rect -1457 -985 -1315 -951
rect -1149 -985 -1007 -951
rect -841 -985 -699 -951
rect -533 -985 -391 -951
rect -225 -985 -83 -951
rect 83 -985 225 -951
rect 391 -985 533 -951
rect 699 -985 841 -951
rect 1007 -985 1149 -951
rect 1315 -985 1457 -951
rect 1623 -985 1765 -951
rect 1931 -985 2073 -951
rect 2239 -985 2381 -951
rect 2547 -985 2689 -951
<< locali >>
rect -2789 964 -2755 980
rect -2789 -908 -2755 -892
rect -2481 964 -2447 980
rect -2481 -908 -2447 -892
rect -2173 964 -2139 980
rect -2173 -908 -2139 -892
rect -1865 964 -1831 980
rect -1865 -908 -1831 -892
rect -1557 964 -1523 980
rect -1557 -908 -1523 -892
rect -1249 964 -1215 980
rect -1249 -908 -1215 -892
rect -941 964 -907 980
rect -941 -908 -907 -892
rect -633 964 -599 980
rect -633 -908 -599 -892
rect -325 964 -291 980
rect -325 -908 -291 -892
rect -17 964 17 980
rect -17 -908 17 -892
rect 291 964 325 980
rect 291 -908 325 -892
rect 599 964 633 980
rect 599 -908 633 -892
rect 907 964 941 980
rect 907 -908 941 -892
rect 1215 964 1249 980
rect 1215 -908 1249 -892
rect 1523 964 1557 980
rect 1523 -908 1557 -892
rect 1831 964 1865 980
rect 1831 -908 1865 -892
rect 2139 964 2173 980
rect 2139 -908 2173 -892
rect 2447 964 2481 980
rect 2447 -908 2481 -892
rect 2755 964 2789 980
rect 2755 -908 2789 -892
rect -2705 -985 -2689 -951
rect -2547 -985 -2531 -951
rect -2397 -985 -2381 -951
rect -2239 -985 -2223 -951
rect -2089 -985 -2073 -951
rect -1931 -985 -1915 -951
rect -1781 -985 -1765 -951
rect -1623 -985 -1607 -951
rect -1473 -985 -1457 -951
rect -1315 -985 -1299 -951
rect -1165 -985 -1149 -951
rect -1007 -985 -991 -951
rect -857 -985 -841 -951
rect -699 -985 -683 -951
rect -549 -985 -533 -951
rect -391 -985 -375 -951
rect -241 -985 -225 -951
rect -83 -985 -67 -951
rect 67 -985 83 -951
rect 225 -985 241 -951
rect 375 -985 391 -951
rect 533 -985 549 -951
rect 683 -985 699 -951
rect 841 -985 857 -951
rect 991 -985 1007 -951
rect 1149 -985 1165 -951
rect 1299 -985 1315 -951
rect 1457 -985 1473 -951
rect 1607 -985 1623 -951
rect 1765 -985 1781 -951
rect 1915 -985 1931 -951
rect 2073 -985 2089 -951
rect 2223 -985 2239 -951
rect 2381 -985 2397 -951
rect 2531 -985 2547 -951
rect 2689 -985 2705 -951
<< viali >>
rect -2789 -892 -2755 964
rect -2481 -892 -2447 964
rect -2173 -892 -2139 964
rect -1865 -892 -1831 964
rect -1557 -892 -1523 964
rect -1249 -892 -1215 964
rect -941 -892 -907 964
rect -633 -892 -599 964
rect -325 -892 -291 964
rect -17 -892 17 964
rect 291 -892 325 964
rect 599 -892 633 964
rect 907 -892 941 964
rect 1215 -892 1249 964
rect 1523 -892 1557 964
rect 1831 -892 1865 964
rect 2139 -892 2173 964
rect 2447 -892 2481 964
rect 2755 -892 2789 964
rect -2689 -985 -2547 -951
rect -2381 -985 -2239 -951
rect -2073 -985 -1931 -951
rect -1765 -985 -1623 -951
rect -1457 -985 -1315 -951
rect -1149 -985 -1007 -951
rect -841 -985 -699 -951
rect -533 -985 -391 -951
rect -225 -985 -83 -951
rect 83 -985 225 -951
rect 391 -985 533 -951
rect 699 -985 841 -951
rect 1007 -985 1149 -951
rect 1315 -985 1457 -951
rect 1623 -985 1765 -951
rect 1931 -985 2073 -951
rect 2239 -985 2381 -951
rect 2547 -985 2689 -951
<< metal1 >>
rect -2795 964 -2749 976
rect -2795 -892 -2789 964
rect -2755 -892 -2749 964
rect -2795 -904 -2749 -892
rect -2487 964 -2441 976
rect -2487 -892 -2481 964
rect -2447 -892 -2441 964
rect -2487 -904 -2441 -892
rect -2179 964 -2133 976
rect -2179 -892 -2173 964
rect -2139 -892 -2133 964
rect -2179 -904 -2133 -892
rect -1871 964 -1825 976
rect -1871 -892 -1865 964
rect -1831 -892 -1825 964
rect -1871 -904 -1825 -892
rect -1563 964 -1517 976
rect -1563 -892 -1557 964
rect -1523 -892 -1517 964
rect -1563 -904 -1517 -892
rect -1255 964 -1209 976
rect -1255 -892 -1249 964
rect -1215 -892 -1209 964
rect -1255 -904 -1209 -892
rect -947 964 -901 976
rect -947 -892 -941 964
rect -907 -892 -901 964
rect -947 -904 -901 -892
rect -639 964 -593 976
rect -639 -892 -633 964
rect -599 -892 -593 964
rect -639 -904 -593 -892
rect -331 964 -285 976
rect -331 -892 -325 964
rect -291 -892 -285 964
rect -331 -904 -285 -892
rect -23 964 23 976
rect -23 -892 -17 964
rect 17 -892 23 964
rect -23 -904 23 -892
rect 285 964 331 976
rect 285 -892 291 964
rect 325 -892 331 964
rect 285 -904 331 -892
rect 593 964 639 976
rect 593 -892 599 964
rect 633 -892 639 964
rect 593 -904 639 -892
rect 901 964 947 976
rect 901 -892 907 964
rect 941 -892 947 964
rect 901 -904 947 -892
rect 1209 964 1255 976
rect 1209 -892 1215 964
rect 1249 -892 1255 964
rect 1209 -904 1255 -892
rect 1517 964 1563 976
rect 1517 -892 1523 964
rect 1557 -892 1563 964
rect 1517 -904 1563 -892
rect 1825 964 1871 976
rect 1825 -892 1831 964
rect 1865 -892 1871 964
rect 1825 -904 1871 -892
rect 2133 964 2179 976
rect 2133 -892 2139 964
rect 2173 -892 2179 964
rect 2133 -904 2179 -892
rect 2441 964 2487 976
rect 2441 -892 2447 964
rect 2481 -892 2487 964
rect 2441 -904 2487 -892
rect 2749 964 2795 976
rect 2749 -892 2755 964
rect 2789 -892 2795 964
rect 2749 -904 2795 -892
rect -2701 -951 -2535 -945
rect -2701 -985 -2689 -951
rect -2547 -985 -2535 -951
rect -2701 -991 -2535 -985
rect -2393 -951 -2227 -945
rect -2393 -985 -2381 -951
rect -2239 -985 -2227 -951
rect -2393 -991 -2227 -985
rect -2085 -951 -1919 -945
rect -2085 -985 -2073 -951
rect -1931 -985 -1919 -951
rect -2085 -991 -1919 -985
rect -1777 -951 -1611 -945
rect -1777 -985 -1765 -951
rect -1623 -985 -1611 -951
rect -1777 -991 -1611 -985
rect -1469 -951 -1303 -945
rect -1469 -985 -1457 -951
rect -1315 -985 -1303 -951
rect -1469 -991 -1303 -985
rect -1161 -951 -995 -945
rect -1161 -985 -1149 -951
rect -1007 -985 -995 -951
rect -1161 -991 -995 -985
rect -853 -951 -687 -945
rect -853 -985 -841 -951
rect -699 -985 -687 -951
rect -853 -991 -687 -985
rect -545 -951 -379 -945
rect -545 -985 -533 -951
rect -391 -985 -379 -951
rect -545 -991 -379 -985
rect -237 -951 -71 -945
rect -237 -985 -225 -951
rect -83 -985 -71 -951
rect -237 -991 -71 -985
rect 71 -951 237 -945
rect 71 -985 83 -951
rect 225 -985 237 -951
rect 71 -991 237 -985
rect 379 -951 545 -945
rect 379 -985 391 -951
rect 533 -985 545 -951
rect 379 -991 545 -985
rect 687 -951 853 -945
rect 687 -985 699 -951
rect 841 -985 853 -951
rect 687 -991 853 -985
rect 995 -951 1161 -945
rect 995 -985 1007 -951
rect 1149 -985 1161 -951
rect 995 -991 1161 -985
rect 1303 -951 1469 -945
rect 1303 -985 1315 -951
rect 1457 -985 1469 -951
rect 1303 -991 1469 -985
rect 1611 -951 1777 -945
rect 1611 -985 1623 -951
rect 1765 -985 1777 -951
rect 1611 -991 1777 -985
rect 1919 -951 2085 -945
rect 1919 -985 1931 -951
rect 2073 -985 2085 -951
rect 1919 -991 2085 -985
rect 2227 -951 2393 -945
rect 2227 -985 2239 -951
rect 2381 -985 2393 -951
rect 2227 -991 2393 -985
rect 2535 -951 2701 -945
rect 2535 -985 2547 -951
rect 2689 -985 2701 -951
rect 2535 -991 2701 -985
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9.4 l 1.25 m 1 nf 18 diffcov 100 polycov 65 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 65 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
