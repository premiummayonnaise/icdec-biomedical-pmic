magic
tech sky130A
magscale 1 2
timestamp 1769400417
<< nwell >>
rect -1297 -334 1297 368
<< pmos >>
rect -1203 -234 -953 306
rect -895 -234 -645 306
rect -587 -234 -337 306
rect -279 -234 -29 306
rect 29 -234 279 306
rect 337 -234 587 306
rect 645 -234 895 306
rect 953 -234 1203 306
<< pdiff >>
rect -1261 294 -1203 306
rect -1261 -222 -1249 294
rect -1215 -222 -1203 294
rect -1261 -234 -1203 -222
rect -953 294 -895 306
rect -953 -222 -941 294
rect -907 -222 -895 294
rect -953 -234 -895 -222
rect -645 294 -587 306
rect -645 -222 -633 294
rect -599 -222 -587 294
rect -645 -234 -587 -222
rect -337 294 -279 306
rect -337 -222 -325 294
rect -291 -222 -279 294
rect -337 -234 -279 -222
rect -29 294 29 306
rect -29 -222 -17 294
rect 17 -222 29 294
rect -29 -234 29 -222
rect 279 294 337 306
rect 279 -222 291 294
rect 325 -222 337 294
rect 279 -234 337 -222
rect 587 294 645 306
rect 587 -222 599 294
rect 633 -222 645 294
rect 587 -234 645 -222
rect 895 294 953 306
rect 895 -222 907 294
rect 941 -222 953 294
rect 895 -234 953 -222
rect 1203 294 1261 306
rect 1203 -222 1215 294
rect 1249 -222 1261 294
rect 1203 -234 1261 -222
<< pdiffc >>
rect -1249 -222 -1215 294
rect -941 -222 -907 294
rect -633 -222 -599 294
rect -325 -222 -291 294
rect -17 -222 17 294
rect 291 -222 325 294
rect 599 -222 633 294
rect 907 -222 941 294
rect 1215 -222 1249 294
<< poly >>
rect -1203 306 -953 332
rect -895 306 -645 332
rect -587 306 -337 332
rect -279 306 -29 332
rect 29 306 279 332
rect 337 306 587 332
rect 645 306 895 332
rect 953 306 1203 332
rect -1203 -281 -953 -234
rect -1203 -315 -1187 -281
rect -969 -315 -953 -281
rect -1203 -331 -953 -315
rect -895 -281 -645 -234
rect -895 -315 -879 -281
rect -661 -315 -645 -281
rect -895 -331 -645 -315
rect -587 -281 -337 -234
rect -587 -315 -571 -281
rect -353 -315 -337 -281
rect -587 -331 -337 -315
rect -279 -281 -29 -234
rect -279 -315 -263 -281
rect -45 -315 -29 -281
rect -279 -331 -29 -315
rect 29 -281 279 -234
rect 29 -315 45 -281
rect 263 -315 279 -281
rect 29 -331 279 -315
rect 337 -281 587 -234
rect 337 -315 353 -281
rect 571 -315 587 -281
rect 337 -331 587 -315
rect 645 -281 895 -234
rect 645 -315 661 -281
rect 879 -315 895 -281
rect 645 -331 895 -315
rect 953 -281 1203 -234
rect 953 -315 969 -281
rect 1187 -315 1203 -281
rect 953 -331 1203 -315
<< polycont >>
rect -1187 -315 -969 -281
rect -879 -315 -661 -281
rect -571 -315 -353 -281
rect -263 -315 -45 -281
rect 45 -315 263 -281
rect 353 -315 571 -281
rect 661 -315 879 -281
rect 969 -315 1187 -281
<< locali >>
rect -1249 294 -1215 310
rect -1249 -238 -1215 -222
rect -941 294 -907 310
rect -941 -238 -907 -222
rect -633 294 -599 310
rect -633 -238 -599 -222
rect -325 294 -291 310
rect -325 -238 -291 -222
rect -17 294 17 310
rect -17 -238 17 -222
rect 291 294 325 310
rect 291 -238 325 -222
rect 599 294 633 310
rect 599 -238 633 -222
rect 907 294 941 310
rect 907 -238 941 -222
rect 1215 294 1249 310
rect 1215 -238 1249 -222
rect -1203 -315 -1187 -281
rect -969 -315 -953 -281
rect -895 -315 -879 -281
rect -661 -315 -645 -281
rect -587 -315 -571 -281
rect -353 -315 -337 -281
rect -279 -315 -263 -281
rect -45 -315 -29 -281
rect 29 -315 45 -281
rect 263 -315 279 -281
rect 337 -315 353 -281
rect 571 -315 587 -281
rect 645 -315 661 -281
rect 879 -315 895 -281
rect 953 -315 969 -281
rect 1187 -315 1203 -281
<< viali >>
rect -1249 -222 -1215 294
rect -941 -222 -907 294
rect -633 -222 -599 294
rect -325 -222 -291 294
rect -17 -222 17 294
rect 291 -222 325 294
rect 599 -222 633 294
rect 907 -222 941 294
rect 1215 -222 1249 294
rect -1187 -315 -969 -281
rect -879 -315 -661 -281
rect -571 -315 -353 -281
rect -263 -315 -45 -281
rect 45 -315 263 -281
rect 353 -315 571 -281
rect 661 -315 879 -281
rect 969 -315 1187 -281
<< metal1 >>
rect -1255 294 -1209 306
rect -1255 -222 -1249 294
rect -1215 -222 -1209 294
rect -1255 -234 -1209 -222
rect -947 294 -901 306
rect -947 -222 -941 294
rect -907 -222 -901 294
rect -947 -234 -901 -222
rect -639 294 -593 306
rect -639 -222 -633 294
rect -599 -222 -593 294
rect -639 -234 -593 -222
rect -331 294 -285 306
rect -331 -222 -325 294
rect -291 -222 -285 294
rect -331 -234 -285 -222
rect -23 294 23 306
rect -23 -222 -17 294
rect 17 -222 23 294
rect -23 -234 23 -222
rect 285 294 331 306
rect 285 -222 291 294
rect 325 -222 331 294
rect 285 -234 331 -222
rect 593 294 639 306
rect 593 -222 599 294
rect 633 -222 639 294
rect 593 -234 639 -222
rect 901 294 947 306
rect 901 -222 907 294
rect 941 -222 947 294
rect 901 -234 947 -222
rect 1209 294 1255 306
rect 1209 -222 1215 294
rect 1249 -222 1255 294
rect 1209 -234 1255 -222
rect -1199 -281 -957 -275
rect -1199 -315 -1187 -281
rect -969 -315 -957 -281
rect -1199 -321 -957 -315
rect -891 -281 -649 -275
rect -891 -315 -879 -281
rect -661 -315 -649 -281
rect -891 -321 -649 -315
rect -583 -281 -341 -275
rect -583 -315 -571 -281
rect -353 -315 -341 -281
rect -583 -321 -341 -315
rect -275 -281 -33 -275
rect -275 -315 -263 -281
rect -45 -315 -33 -281
rect -275 -321 -33 -315
rect 33 -281 275 -275
rect 33 -315 45 -281
rect 263 -315 275 -281
rect 33 -321 275 -315
rect 341 -281 583 -275
rect 341 -315 353 -281
rect 571 -315 583 -281
rect 341 -321 583 -315
rect 649 -281 891 -275
rect 649 -315 661 -281
rect 879 -315 891 -281
rect 649 -321 891 -315
rect 957 -281 1199 -275
rect 957 -315 969 -281
rect 1187 -315 1199 -281
rect 957 -321 1199 -315
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.7 l 1.25 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
