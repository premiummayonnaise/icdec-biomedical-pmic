magic
tech sky130A
magscale 1 2
timestamp 1769931968
<< pwell >>
rect -278 -733 278 733
<< mvnmos >>
rect -50 -475 50 475
<< mvndiff >>
rect -108 463 -50 475
rect -108 -463 -96 463
rect -62 -463 -50 463
rect -108 -475 -50 -463
rect 50 463 108 475
rect 50 -463 62 463
rect 96 -463 108 463
rect 50 -475 108 -463
<< mvndiffc >>
rect -96 -463 -62 463
rect 62 -463 96 463
<< mvpsubdiff >>
rect -242 685 242 697
rect -242 651 -134 685
rect 134 651 242 685
rect -242 639 242 651
rect -242 589 -184 639
rect -242 -589 -230 589
rect -196 -589 -184 589
rect 184 589 242 639
rect -242 -639 -184 -589
rect 184 -589 196 589
rect 230 -589 242 589
rect 184 -639 242 -589
rect -242 -651 242 -639
rect -242 -685 -134 -651
rect 134 -685 242 -651
rect -242 -697 242 -685
<< mvpsubdiffcont >>
rect -134 651 134 685
rect -230 -589 -196 589
rect 196 -589 230 589
rect -134 -685 134 -651
<< poly >>
rect -50 547 50 563
rect -50 513 -34 547
rect 34 513 50 547
rect -50 475 50 513
rect -50 -513 50 -475
rect -50 -547 -34 -513
rect 34 -547 50 -513
rect -50 -563 50 -547
<< polycont >>
rect -34 513 34 547
rect -34 -547 34 -513
<< locali >>
rect -230 651 -134 685
rect 134 651 230 685
rect -230 589 -196 651
rect 196 589 230 651
rect -50 513 -34 547
rect 34 513 50 547
rect -96 463 -62 479
rect -96 -479 -62 -463
rect 62 463 96 479
rect 62 -479 96 -463
rect -50 -547 -34 -513
rect 34 -547 50 -513
rect -230 -651 -196 -589
rect 196 -651 230 -589
rect -230 -685 -134 -651
rect 134 -685 230 -651
<< viali >>
rect -34 513 34 547
rect -96 -463 -62 463
rect 62 -463 96 463
rect -34 -547 34 -513
<< metal1 >>
rect -46 547 46 553
rect -46 513 -34 547
rect 34 513 46 547
rect -46 507 46 513
rect -102 463 -56 475
rect -102 -463 -96 463
rect -62 -463 -56 463
rect -102 -475 -56 -463
rect 56 463 102 475
rect 56 -463 62 463
rect 96 -463 102 463
rect 56 -475 102 -463
rect -46 -513 46 -507
rect -46 -547 -34 -513
rect 34 -547 46 -513
rect -46 -553 46 -547
<< properties >>
string FIXED_BBOX -213 -668 213 668
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.75 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
