magic
tech sky130A
magscale 1 2
timestamp 1769931968
<< pwell >>
rect -357 -2158 357 2158
<< mvnmos >>
rect -129 -1900 -29 1900
rect 29 -1900 129 1900
<< mvndiff >>
rect -187 1888 -129 1900
rect -187 -1888 -175 1888
rect -141 -1888 -129 1888
rect -187 -1900 -129 -1888
rect -29 1888 29 1900
rect -29 -1888 -17 1888
rect 17 -1888 29 1888
rect -29 -1900 29 -1888
rect 129 1888 187 1900
rect 129 -1888 141 1888
rect 175 -1888 187 1888
rect 129 -1900 187 -1888
<< mvndiffc >>
rect -175 -1888 -141 1888
rect -17 -1888 17 1888
rect 141 -1888 175 1888
<< mvpsubdiff >>
rect -321 2110 321 2122
rect -321 2076 -213 2110
rect 213 2076 321 2110
rect -321 2064 321 2076
rect -321 2014 -263 2064
rect -321 -2014 -309 2014
rect -275 -2014 -263 2014
rect 263 2014 321 2064
rect -321 -2064 -263 -2014
rect 263 -2014 275 2014
rect 309 -2014 321 2014
rect 263 -2064 321 -2014
rect -321 -2076 321 -2064
rect -321 -2110 -213 -2076
rect 213 -2110 321 -2076
rect -321 -2122 321 -2110
<< mvpsubdiffcont >>
rect -213 2076 213 2110
rect -309 -2014 -275 2014
rect 275 -2014 309 2014
rect -213 -2110 213 -2076
<< poly >>
rect -129 1972 -29 1988
rect -129 1938 -113 1972
rect -45 1938 -29 1972
rect -129 1900 -29 1938
rect 29 1972 129 1988
rect 29 1938 45 1972
rect 113 1938 129 1972
rect 29 1900 129 1938
rect -129 -1938 -29 -1900
rect -129 -1972 -113 -1938
rect -45 -1972 -29 -1938
rect -129 -1988 -29 -1972
rect 29 -1938 129 -1900
rect 29 -1972 45 -1938
rect 113 -1972 129 -1938
rect 29 -1988 129 -1972
<< polycont >>
rect -113 1938 -45 1972
rect 45 1938 113 1972
rect -113 -1972 -45 -1938
rect 45 -1972 113 -1938
<< locali >>
rect -309 2076 -213 2110
rect 213 2076 309 2110
rect -309 2014 -275 2076
rect 275 2014 309 2076
rect -129 1938 -113 1972
rect -45 1938 -29 1972
rect 29 1938 45 1972
rect 113 1938 129 1972
rect -175 1888 -141 1904
rect -175 -1904 -141 -1888
rect -17 1888 17 1904
rect -17 -1904 17 -1888
rect 141 1888 175 1904
rect 141 -1904 175 -1888
rect -129 -1972 -113 -1938
rect -45 -1972 -29 -1938
rect 29 -1972 45 -1938
rect 113 -1972 129 -1938
rect -309 -2076 -275 -2014
rect 275 -2076 309 -2014
rect -309 -2110 -213 -2076
rect 213 -2110 309 -2076
<< viali >>
rect -113 1938 -45 1972
rect 45 1938 113 1972
rect -175 -1888 -141 1888
rect -17 -1888 17 1888
rect 141 -1888 175 1888
rect -113 -1972 -45 -1938
rect 45 -1972 113 -1938
<< metal1 >>
rect -125 1972 -33 1978
rect -125 1938 -113 1972
rect -45 1938 -33 1972
rect -125 1932 -33 1938
rect 33 1972 125 1978
rect 33 1938 45 1972
rect 113 1938 125 1972
rect 33 1932 125 1938
rect -181 1888 -135 1900
rect -181 -1888 -175 1888
rect -141 -1888 -135 1888
rect -181 -1900 -135 -1888
rect -23 1888 23 1900
rect -23 -1888 -17 1888
rect 17 -1888 23 1888
rect -23 -1900 23 -1888
rect 135 1888 181 1900
rect 135 -1888 141 1888
rect 175 -1888 181 1888
rect 135 -1900 181 -1888
rect -125 -1938 -33 -1932
rect -125 -1972 -113 -1938
rect -45 -1972 -33 -1938
rect -125 -1978 -33 -1972
rect 33 -1938 125 -1932
rect 33 -1972 45 -1938
rect 113 -1972 125 -1938
rect 33 -1978 125 -1972
<< properties >>
string FIXED_BBOX -292 -2093 292 2093
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 19.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
