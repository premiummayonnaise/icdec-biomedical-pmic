magic
tech sky130A
magscale 1 2
timestamp 1769529800
<< pwell >>
rect -831 -729 831 729
<< mvnmos >>
rect -603 -471 -503 471
rect -445 -471 -345 471
rect -287 -471 -187 471
rect -129 -471 -29 471
rect 29 -471 129 471
rect 187 -471 287 471
rect 345 -471 445 471
rect 503 -471 603 471
<< mvndiff >>
rect -661 459 -603 471
rect -661 -459 -649 459
rect -615 -459 -603 459
rect -661 -471 -603 -459
rect -503 459 -445 471
rect -503 -459 -491 459
rect -457 -459 -445 459
rect -503 -471 -445 -459
rect -345 459 -287 471
rect -345 -459 -333 459
rect -299 -459 -287 459
rect -345 -471 -287 -459
rect -187 459 -129 471
rect -187 -459 -175 459
rect -141 -459 -129 459
rect -187 -471 -129 -459
rect -29 459 29 471
rect -29 -459 -17 459
rect 17 -459 29 459
rect -29 -471 29 -459
rect 129 459 187 471
rect 129 -459 141 459
rect 175 -459 187 459
rect 129 -471 187 -459
rect 287 459 345 471
rect 287 -459 299 459
rect 333 -459 345 459
rect 287 -471 345 -459
rect 445 459 503 471
rect 445 -459 457 459
rect 491 -459 503 459
rect 445 -471 503 -459
rect 603 459 661 471
rect 603 -459 615 459
rect 649 -459 661 459
rect 603 -471 661 -459
<< mvndiffc >>
rect -649 -459 -615 459
rect -491 -459 -457 459
rect -333 -459 -299 459
rect -175 -459 -141 459
rect -17 -459 17 459
rect 141 -459 175 459
rect 299 -459 333 459
rect 457 -459 491 459
rect 615 -459 649 459
<< mvpsubdiff >>
rect -795 681 795 693
rect -795 647 -687 681
rect 687 647 795 681
rect -795 635 795 647
rect -795 585 -737 635
rect -795 -585 -783 585
rect -749 -585 -737 585
rect 737 585 795 635
rect -795 -635 -737 -585
rect 737 -585 749 585
rect 783 -585 795 585
rect 737 -635 795 -585
rect -795 -647 795 -635
rect -795 -681 -687 -647
rect 687 -681 795 -647
rect -795 -693 795 -681
<< mvpsubdiffcont >>
rect -687 647 687 681
rect -783 -585 -749 585
rect 749 -585 783 585
rect -687 -681 687 -647
<< poly >>
rect -603 543 -503 559
rect -603 509 -587 543
rect -519 509 -503 543
rect -603 471 -503 509
rect -445 543 -345 559
rect -445 509 -429 543
rect -361 509 -345 543
rect -445 471 -345 509
rect -287 543 -187 559
rect -287 509 -271 543
rect -203 509 -187 543
rect -287 471 -187 509
rect -129 543 -29 559
rect -129 509 -113 543
rect -45 509 -29 543
rect -129 471 -29 509
rect 29 543 129 559
rect 29 509 45 543
rect 113 509 129 543
rect 29 471 129 509
rect 187 543 287 559
rect 187 509 203 543
rect 271 509 287 543
rect 187 471 287 509
rect 345 543 445 559
rect 345 509 361 543
rect 429 509 445 543
rect 345 471 445 509
rect 503 543 603 559
rect 503 509 519 543
rect 587 509 603 543
rect 503 471 603 509
rect -603 -509 -503 -471
rect -603 -543 -587 -509
rect -519 -543 -503 -509
rect -603 -559 -503 -543
rect -445 -509 -345 -471
rect -445 -543 -429 -509
rect -361 -543 -345 -509
rect -445 -559 -345 -543
rect -287 -509 -187 -471
rect -287 -543 -271 -509
rect -203 -543 -187 -509
rect -287 -559 -187 -543
rect -129 -509 -29 -471
rect -129 -543 -113 -509
rect -45 -543 -29 -509
rect -129 -559 -29 -543
rect 29 -509 129 -471
rect 29 -543 45 -509
rect 113 -543 129 -509
rect 29 -559 129 -543
rect 187 -509 287 -471
rect 187 -543 203 -509
rect 271 -543 287 -509
rect 187 -559 287 -543
rect 345 -509 445 -471
rect 345 -543 361 -509
rect 429 -543 445 -509
rect 345 -559 445 -543
rect 503 -509 603 -471
rect 503 -543 519 -509
rect 587 -543 603 -509
rect 503 -559 603 -543
<< polycont >>
rect -587 509 -519 543
rect -429 509 -361 543
rect -271 509 -203 543
rect -113 509 -45 543
rect 45 509 113 543
rect 203 509 271 543
rect 361 509 429 543
rect 519 509 587 543
rect -587 -543 -519 -509
rect -429 -543 -361 -509
rect -271 -543 -203 -509
rect -113 -543 -45 -509
rect 45 -543 113 -509
rect 203 -543 271 -509
rect 361 -543 429 -509
rect 519 -543 587 -509
<< locali >>
rect -783 647 -687 681
rect 687 647 783 681
rect -783 585 -749 647
rect 749 585 783 647
rect -603 509 -587 543
rect -519 509 -503 543
rect -445 509 -429 543
rect -361 509 -345 543
rect -287 509 -271 543
rect -203 509 -187 543
rect -129 509 -113 543
rect -45 509 -29 543
rect 29 509 45 543
rect 113 509 129 543
rect 187 509 203 543
rect 271 509 287 543
rect 345 509 361 543
rect 429 509 445 543
rect 503 509 519 543
rect 587 509 603 543
rect -649 459 -615 475
rect -649 -475 -615 -459
rect -491 459 -457 475
rect -491 -475 -457 -459
rect -333 459 -299 475
rect -333 -475 -299 -459
rect -175 459 -141 475
rect -175 -475 -141 -459
rect -17 459 17 475
rect -17 -475 17 -459
rect 141 459 175 475
rect 141 -475 175 -459
rect 299 459 333 475
rect 299 -475 333 -459
rect 457 459 491 475
rect 457 -475 491 -459
rect 615 459 649 475
rect 615 -475 649 -459
rect -603 -543 -587 -509
rect -519 -543 -503 -509
rect -445 -543 -429 -509
rect -361 -543 -345 -509
rect -287 -543 -271 -509
rect -203 -543 -187 -509
rect -129 -543 -113 -509
rect -45 -543 -29 -509
rect 29 -543 45 -509
rect 113 -543 129 -509
rect 187 -543 203 -509
rect 271 -543 287 -509
rect 345 -543 361 -509
rect 429 -543 445 -509
rect 503 -543 519 -509
rect 587 -543 603 -509
rect -783 -647 -749 -585
rect 749 -647 783 -585
rect -783 -681 -687 -647
rect 687 -681 783 -647
<< viali >>
rect -587 509 -519 543
rect -429 509 -361 543
rect -271 509 -203 543
rect -113 509 -45 543
rect 45 509 113 543
rect 203 509 271 543
rect 361 509 429 543
rect 519 509 587 543
rect -649 -459 -615 459
rect -491 -459 -457 459
rect -333 -459 -299 459
rect -175 -459 -141 459
rect -17 -459 17 459
rect 141 -459 175 459
rect 299 -459 333 459
rect 457 -459 491 459
rect 615 -459 649 459
rect -587 -543 -519 -509
rect -429 -543 -361 -509
rect -271 -543 -203 -509
rect -113 -543 -45 -509
rect 45 -543 113 -509
rect 203 -543 271 -509
rect 361 -543 429 -509
rect 519 -543 587 -509
<< metal1 >>
rect -599 543 -507 549
rect -599 509 -587 543
rect -519 509 -507 543
rect -599 503 -507 509
rect -441 543 -349 549
rect -441 509 -429 543
rect -361 509 -349 543
rect -441 503 -349 509
rect -283 543 -191 549
rect -283 509 -271 543
rect -203 509 -191 543
rect -283 503 -191 509
rect -125 543 -33 549
rect -125 509 -113 543
rect -45 509 -33 543
rect -125 503 -33 509
rect 33 543 125 549
rect 33 509 45 543
rect 113 509 125 543
rect 33 503 125 509
rect 191 543 283 549
rect 191 509 203 543
rect 271 509 283 543
rect 191 503 283 509
rect 349 543 441 549
rect 349 509 361 543
rect 429 509 441 543
rect 349 503 441 509
rect 507 543 599 549
rect 507 509 519 543
rect 587 509 599 543
rect 507 503 599 509
rect -655 459 -609 471
rect -655 -459 -649 459
rect -615 -459 -609 459
rect -655 -471 -609 -459
rect -497 459 -451 471
rect -497 -459 -491 459
rect -457 -459 -451 459
rect -497 -471 -451 -459
rect -339 459 -293 471
rect -339 -459 -333 459
rect -299 -459 -293 459
rect -339 -471 -293 -459
rect -181 459 -135 471
rect -181 -459 -175 459
rect -141 -459 -135 459
rect -181 -471 -135 -459
rect -23 459 23 471
rect -23 -459 -17 459
rect 17 -459 23 459
rect -23 -471 23 -459
rect 135 459 181 471
rect 135 -459 141 459
rect 175 -459 181 459
rect 135 -471 181 -459
rect 293 459 339 471
rect 293 -459 299 459
rect 333 -459 339 459
rect 293 -471 339 -459
rect 451 459 497 471
rect 451 -459 457 459
rect 491 -459 497 459
rect 451 -471 497 -459
rect 609 459 655 471
rect 609 -459 615 459
rect 649 -459 655 459
rect 609 -471 655 -459
rect -599 -509 -507 -503
rect -599 -543 -587 -509
rect -519 -543 -507 -509
rect -599 -549 -507 -543
rect -441 -509 -349 -503
rect -441 -543 -429 -509
rect -361 -543 -349 -509
rect -441 -549 -349 -543
rect -283 -509 -191 -503
rect -283 -543 -271 -509
rect -203 -543 -191 -509
rect -283 -549 -191 -543
rect -125 -509 -33 -503
rect -125 -543 -113 -509
rect -45 -543 -33 -509
rect -125 -549 -33 -543
rect 33 -509 125 -503
rect 33 -543 45 -509
rect 113 -543 125 -509
rect 33 -549 125 -543
rect 191 -509 283 -503
rect 191 -543 203 -509
rect 271 -543 283 -509
rect 191 -549 283 -543
rect 349 -509 441 -503
rect 349 -543 361 -509
rect 429 -543 441 -509
rect 349 -549 441 -543
rect 507 -509 599 -503
rect 507 -543 519 -509
rect 587 -543 599 -509
rect 507 -549 599 -543
<< properties >>
string FIXED_BBOX -766 -664 766 664
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.7125 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
