magic
tech sky130A
magscale 1 2
timestamp 1769089966
<< nwell >>
rect -4514 -5598 1006 -4068
<< pwell >>
rect -4460 -7501 940 -5598
rect -4474 -7530 943 -7501
rect -4475 -7870 943 -7530
rect -4475 -7899 942 -7870
<< psubdiff >>
rect -2700 -5720 -800 -5700
rect -2700 -5780 -2580 -5720
rect -2440 -5780 -2400 -5720
rect -2260 -5780 -2220 -5720
rect -2080 -5780 -2040 -5720
rect -1900 -5780 -1860 -5720
rect -1720 -5780 -1680 -5720
rect -1540 -5780 -1500 -5720
rect -1360 -5780 -1320 -5720
rect -1180 -5780 -1140 -5720
rect -1000 -5780 -960 -5720
rect -840 -5780 -800 -5720
rect -2700 -5800 -800 -5780
rect -2700 -5900 -2600 -5800
rect -2700 -6040 -2680 -5900
rect -2620 -6040 -2600 -5900
rect -2700 -6080 -2600 -6040
rect -2700 -6220 -2680 -6080
rect -2620 -6220 -2600 -6080
rect -2700 -6260 -2600 -6220
rect -2700 -6400 -2680 -6260
rect -2620 -6400 -2600 -6260
rect -2700 -6440 -2600 -6400
rect -2700 -6580 -2680 -6440
rect -2620 -6580 -2600 -6440
rect -2700 -6600 -2600 -6580
rect -900 -5900 -800 -5800
rect -900 -6040 -880 -5900
rect -820 -6040 -800 -5900
rect -900 -6080 -800 -6040
rect -900 -6220 -880 -6080
rect -820 -6220 -800 -6080
rect -900 -6260 -800 -6220
rect -900 -6400 -880 -6260
rect -820 -6400 -800 -6260
rect -900 -6440 -800 -6400
rect -900 -6580 -880 -6440
rect -820 -6580 -800 -6440
rect -900 -6600 -800 -6580
rect -3700 -6620 200 -6600
rect -3700 -6680 -3600 -6620
rect -3240 -6680 -3200 -6620
rect -3060 -6680 -3020 -6620
rect -2880 -6680 -2840 -6620
rect -2700 -6680 -2660 -6620
rect -2520 -6680 -2480 -6620
rect -2340 -6680 -2300 -6620
rect -2160 -6680 -2120 -6620
rect -1980 -6680 -1940 -6620
rect -1800 -6680 -1760 -6620
rect -1620 -6680 -1580 -6620
rect -1440 -6680 -1400 -6620
rect -1260 -6680 -1220 -6620
rect -1080 -6680 -1040 -6620
rect -900 -6680 -860 -6620
rect -720 -6680 -680 -6620
rect -540 -6680 -500 -6620
rect -360 -6680 -320 -6620
rect -180 -6680 -140 -6620
rect 100 -6680 200 -6620
rect -3700 -6700 200 -6680
rect -3700 -6760 -3600 -6700
rect -3700 -6900 -3680 -6760
rect -3620 -6900 -3600 -6760
rect -3700 -6940 -3600 -6900
rect -3700 -7080 -3680 -6940
rect -3620 -7080 -3600 -6940
rect -3700 -7120 -3600 -7080
rect -3700 -7260 -3680 -7120
rect -3620 -7260 -3600 -7120
rect -3700 -7300 -3600 -7260
rect -3700 -7440 -3680 -7300
rect -3620 -7440 -3600 -7300
rect -3700 -7480 -3600 -7440
rect -3700 -7620 -3680 -7480
rect -3620 -7620 -3600 -7480
rect -3700 -7660 -3600 -7620
rect -3700 -7880 -3680 -7660
rect -3620 -7800 -3600 -7660
rect -2700 -6740 -2600 -6700
rect -2700 -6880 -2680 -6740
rect -2620 -6880 -2600 -6740
rect -2700 -6920 -2600 -6880
rect -2700 -7060 -2680 -6920
rect -2620 -7060 -2600 -6920
rect -2700 -7100 -2600 -7060
rect -2700 -7240 -2680 -7100
rect -2620 -7240 -2600 -7100
rect -2700 -7280 -2600 -7240
rect -2700 -7420 -2680 -7280
rect -2620 -7420 -2600 -7280
rect -2700 -7460 -2600 -7420
rect -2700 -7600 -2680 -7460
rect -2620 -7600 -2600 -7460
rect -2700 -7640 -2600 -7600
rect -2700 -7780 -2680 -7640
rect -2620 -7780 -2600 -7640
rect -2700 -7800 -2600 -7780
rect -900 -6740 -800 -6700
rect -900 -6880 -880 -6740
rect -820 -6880 -800 -6740
rect -900 -6920 -800 -6880
rect -900 -7060 -880 -6920
rect -820 -7060 -800 -6920
rect -900 -7100 -800 -7060
rect -900 -7240 -880 -7100
rect -820 -7240 -800 -7100
rect -900 -7280 -800 -7240
rect -900 -7420 -880 -7280
rect -820 -7420 -800 -7280
rect -900 -7460 -800 -7420
rect -900 -7600 -880 -7460
rect -820 -7600 -800 -7460
rect -900 -7640 -800 -7600
rect -900 -7780 -880 -7640
rect -820 -7780 -800 -7640
rect -900 -7800 -800 -7780
rect -3620 -7804 -800 -7800
rect 100 -6760 200 -6700
rect 100 -6900 120 -6760
rect 180 -6900 200 -6760
rect 100 -6940 200 -6900
rect 100 -7080 120 -6940
rect 180 -7080 200 -6940
rect 100 -7120 200 -7080
rect 100 -7260 120 -7120
rect 180 -7260 200 -7120
rect 100 -7300 200 -7260
rect 100 -7440 120 -7300
rect 180 -7440 200 -7300
rect 100 -7480 200 -7440
rect 100 -7620 120 -7480
rect 180 -7620 200 -7480
rect 100 -7660 200 -7620
rect 100 -7804 120 -7660
rect -3620 -7820 120 -7804
rect -3420 -7880 -3380 -7820
rect -3240 -7880 -3200 -7820
rect -3060 -7880 -3020 -7820
rect -2880 -7880 -2840 -7820
rect -2700 -7880 -2660 -7820
rect -2520 -7880 -2480 -7820
rect -2340 -7880 -2300 -7820
rect -2160 -7880 -2120 -7820
rect -1980 -7880 -1940 -7820
rect -1800 -7880 -1760 -7820
rect -1620 -7880 -1580 -7820
rect -1440 -7880 -1400 -7820
rect -1260 -7880 -1220 -7820
rect -1080 -7880 -1040 -7820
rect -900 -7880 -860 -7820
rect -720 -7880 -680 -7820
rect -540 -7880 -500 -7820
rect -360 -7880 -320 -7820
rect -180 -7880 -140 -7820
rect 180 -7880 200 -7660
rect -3700 -7896 200 -7880
rect -3700 -7970 -3500 -7896
rect -2700 -7900 200 -7896
rect -3700 -8000 -3600 -7970
rect -2700 -8000 -2600 -7900
rect -900 -8000 -800 -7900
rect 100 -8000 200 -7900
<< nsubdiff >>
rect -4452 -4140 -4352 -4106
rect -4452 -4200 -4440 -4140
rect -4460 -4300 -4440 -4200
rect -4380 -4200 -4352 -4140
rect -3452 -4140 -3352 -4106
rect -3452 -4200 -3440 -4140
rect -4380 -4220 -3440 -4200
rect -3380 -4200 -3352 -4140
rect -1859 -4140 -1653 -4106
rect -1859 -4200 -1820 -4140
rect -3380 -4220 -1820 -4200
rect -1680 -4200 -1653 -4140
rect -151 -4140 -47 -4106
rect -151 -4200 -140 -4140
rect -1680 -4220 -140 -4200
rect -80 -4200 -47 -4140
rect 848 -4140 948 -4106
rect 848 -4200 860 -4140
rect -80 -4220 860 -4200
rect 920 -4200 948 -4140
rect -4100 -4280 -4060 -4220
rect -3840 -4280 -3800 -4220
rect -3580 -4280 -3520 -4220
rect -3300 -4280 -3260 -4220
rect -3040 -4280 -2980 -4220
rect -2760 -4280 -2720 -4220
rect -2500 -4280 -2460 -4220
rect -2240 -4280 -2200 -4220
rect -1980 -4280 -1940 -4220
rect -1460 -4280 -1420 -4220
rect -1200 -4280 -1160 -4220
rect -940 -4280 -900 -4220
rect -680 -4280 -640 -4220
rect -420 -4280 -340 -4220
rect 120 -4280 160 -4220
rect 300 -4280 340 -4220
rect 480 -4280 520 -4220
rect 660 -4280 700 -4220
rect 920 -4280 960 -4200
rect -4452 -4460 -4440 -4300
rect -4380 -4300 -1820 -4280
rect -4380 -4460 -4352 -4300
rect -4452 -4500 -4352 -4460
rect -4452 -4640 -4440 -4500
rect -4380 -4640 -4352 -4500
rect -4452 -4680 -4352 -4640
rect -4452 -4820 -4440 -4680
rect -4380 -4820 -4352 -4680
rect -4452 -4860 -4352 -4820
rect -4452 -5000 -4440 -4860
rect -4380 -5000 -4352 -4860
rect -4452 -5040 -4352 -5000
rect -4452 -5180 -4440 -5040
rect -4380 -5180 -4352 -5040
rect -4452 -5220 -4352 -5180
rect -4452 -5460 -4440 -5220
rect -4380 -5386 -4352 -5220
rect -3452 -4320 -3352 -4300
rect -3452 -4460 -3440 -4320
rect -3380 -4460 -3352 -4320
rect -3452 -4500 -3352 -4460
rect -3452 -4640 -3440 -4500
rect -3380 -4640 -3352 -4500
rect -3452 -4680 -3352 -4640
rect -3452 -4820 -3440 -4680
rect -3380 -4820 -3352 -4680
rect -3452 -4860 -3352 -4820
rect -1859 -4420 -1820 -4300
rect -1680 -4300 960 -4280
rect -1680 -4386 -1653 -4300
rect -151 -4320 -47 -4300
rect -151 -4386 -140 -4320
rect -1680 -4420 -1652 -4386
rect -1859 -4460 -1652 -4420
rect -1859 -4740 -1820 -4460
rect -1680 -4740 -1652 -4460
rect -1859 -4780 -1652 -4740
rect -1859 -4829 -1820 -4780
rect -3452 -5000 -3440 -4860
rect -3380 -5000 -3352 -4860
rect -3452 -5040 -3352 -5000
rect -3452 -5180 -3440 -5040
rect -3380 -5180 -3352 -5040
rect -3452 -5220 -3352 -5180
rect -3452 -5360 -3440 -5220
rect -3380 -5360 -3352 -5220
rect -3452 -5386 -3352 -5360
rect -1852 -5060 -1820 -4829
rect -1680 -5060 -1652 -4780
rect -1852 -5100 -1652 -5060
rect -1852 -5386 -1820 -5100
rect -4380 -5400 -1820 -5386
rect -1680 -5386 -1652 -5100
rect -152 -4460 -140 -4386
rect -80 -4460 -47 -4320
rect -152 -4500 -47 -4460
rect -152 -4640 -140 -4500
rect -80 -4640 -47 -4500
rect -152 -4680 -47 -4640
rect -152 -4820 -140 -4680
rect -80 -4820 -47 -4680
rect -152 -4857 -47 -4820
rect 848 -4320 948 -4300
rect 848 -4460 860 -4320
rect 920 -4460 948 -4320
rect 848 -4500 948 -4460
rect 848 -4640 860 -4500
rect 920 -4640 948 -4500
rect 848 -4680 948 -4640
rect 848 -4820 860 -4680
rect 920 -4820 948 -4680
rect -152 -4860 -52 -4857
rect -152 -5000 -140 -4860
rect -80 -5000 -52 -4860
rect -152 -5040 -52 -5000
rect -152 -5180 -140 -5040
rect -80 -5180 -52 -5040
rect -152 -5220 -52 -5180
rect -152 -5360 -140 -5220
rect -80 -5360 -52 -5220
rect -152 -5386 -52 -5360
rect 848 -4860 948 -4820
rect 848 -5000 860 -4860
rect 920 -5000 948 -4860
rect 848 -5040 948 -5000
rect 848 -5180 860 -5040
rect 920 -5180 948 -5040
rect 848 -5220 948 -5180
rect 848 -5386 860 -5220
rect -1680 -5400 860 -5386
rect -4120 -5460 -4080 -5400
rect -3860 -5460 -3820 -5400
rect -3600 -5460 -3560 -5400
rect -3340 -5460 -3300 -5400
rect -3080 -5460 -3040 -5400
rect -2820 -5460 -2780 -5400
rect -2560 -5460 -2520 -5400
rect -2300 -5460 -2260 -5400
rect -2040 -5460 -2000 -5400
rect -1500 -5460 -1460 -5400
rect -1240 -5460 -1200 -5400
rect -980 -5460 -940 -5400
rect -720 -5460 -680 -5400
rect -460 -5460 -420 -5400
rect -200 -5460 -160 -5400
rect 60 -5460 100 -5400
rect 320 -5460 360 -5400
rect 580 -5460 620 -5400
rect 920 -5460 948 -5220
rect -4452 -5486 948 -5460
<< psubdiffcont >>
rect -2580 -5780 -2440 -5720
rect -2400 -5780 -2260 -5720
rect -2220 -5780 -2080 -5720
rect -2040 -5780 -1900 -5720
rect -1860 -5780 -1720 -5720
rect -1680 -5780 -1540 -5720
rect -1500 -5780 -1360 -5720
rect -1320 -5780 -1180 -5720
rect -1140 -5780 -1000 -5720
rect -960 -5780 -840 -5720
rect -2680 -6040 -2620 -5900
rect -2680 -6220 -2620 -6080
rect -2680 -6400 -2620 -6260
rect -2680 -6580 -2620 -6440
rect -880 -6040 -820 -5900
rect -880 -6220 -820 -6080
rect -880 -6400 -820 -6260
rect -880 -6580 -820 -6440
rect -3600 -6680 -3240 -6620
rect -3200 -6680 -3060 -6620
rect -3020 -6680 -2880 -6620
rect -2840 -6680 -2700 -6620
rect -2660 -6680 -2520 -6620
rect -2480 -6680 -2340 -6620
rect -2300 -6680 -2160 -6620
rect -2120 -6680 -1980 -6620
rect -1940 -6680 -1800 -6620
rect -1760 -6680 -1620 -6620
rect -1580 -6680 -1440 -6620
rect -1400 -6680 -1260 -6620
rect -1220 -6680 -1080 -6620
rect -1040 -6680 -900 -6620
rect -860 -6680 -720 -6620
rect -680 -6680 -540 -6620
rect -500 -6680 -360 -6620
rect -320 -6680 -180 -6620
rect -140 -6680 100 -6620
rect -3680 -6900 -3620 -6760
rect -3680 -7080 -3620 -6940
rect -3680 -7260 -3620 -7120
rect -3680 -7440 -3620 -7300
rect -3680 -7620 -3620 -7480
rect -3680 -7820 -3620 -7660
rect -2680 -6880 -2620 -6740
rect -2680 -7060 -2620 -6920
rect -2680 -7240 -2620 -7100
rect -2680 -7420 -2620 -7280
rect -2680 -7600 -2620 -7460
rect -2680 -7780 -2620 -7640
rect -880 -6880 -820 -6740
rect -880 -7060 -820 -6920
rect -880 -7240 -820 -7100
rect -880 -7420 -820 -7280
rect -880 -7600 -820 -7460
rect -880 -7780 -820 -7640
rect 120 -6900 180 -6760
rect 120 -7080 180 -6940
rect 120 -7260 180 -7120
rect 120 -7440 180 -7300
rect 120 -7620 180 -7480
rect 120 -7820 180 -7660
rect -3680 -7880 -3420 -7820
rect -3380 -7880 -3240 -7820
rect -3200 -7880 -3060 -7820
rect -3020 -7880 -2880 -7820
rect -2840 -7880 -2700 -7820
rect -2660 -7880 -2520 -7820
rect -2480 -7880 -2340 -7820
rect -2300 -7880 -2160 -7820
rect -2120 -7880 -1980 -7820
rect -1940 -7880 -1800 -7820
rect -1760 -7880 -1620 -7820
rect -1580 -7880 -1440 -7820
rect -1400 -7880 -1260 -7820
rect -1220 -7880 -1080 -7820
rect -1040 -7880 -900 -7820
rect -860 -7880 -720 -7820
rect -680 -7880 -540 -7820
rect -500 -7880 -360 -7820
rect -320 -7880 -180 -7820
rect -140 -7880 180 -7820
<< nsubdiffcont >>
rect -4440 -4220 -4380 -4140
rect -3440 -4220 -3380 -4140
rect -1820 -4220 -1680 -4140
rect -140 -4220 -80 -4140
rect 860 -4220 920 -4140
rect -4440 -4280 -4100 -4220
rect -4060 -4280 -3840 -4220
rect -3800 -4280 -3580 -4220
rect -3520 -4280 -3300 -4220
rect -3260 -4280 -3040 -4220
rect -2980 -4280 -2760 -4220
rect -2720 -4280 -2500 -4220
rect -2460 -4280 -2240 -4220
rect -2200 -4280 -1980 -4220
rect -1940 -4280 -1460 -4220
rect -1420 -4280 -1200 -4220
rect -1160 -4280 -940 -4220
rect -900 -4280 -680 -4220
rect -640 -4280 -420 -4220
rect -340 -4280 120 -4220
rect 160 -4280 300 -4220
rect 340 -4280 480 -4220
rect 520 -4280 660 -4220
rect 700 -4280 920 -4220
rect -4440 -4460 -4380 -4280
rect -4440 -4640 -4380 -4500
rect -4440 -4820 -4380 -4680
rect -4440 -5000 -4380 -4860
rect -4440 -5180 -4380 -5040
rect -4440 -5400 -4380 -5220
rect -3440 -4460 -3380 -4320
rect -3440 -4640 -3380 -4500
rect -3440 -4820 -3380 -4680
rect -1820 -4420 -1680 -4280
rect -1820 -4740 -1680 -4460
rect -3440 -5000 -3380 -4860
rect -3440 -5180 -3380 -5040
rect -3440 -5360 -3380 -5220
rect -1820 -5060 -1680 -4780
rect -1820 -5400 -1680 -5100
rect -140 -4460 -80 -4320
rect -140 -4640 -80 -4500
rect -140 -4820 -80 -4680
rect 860 -4460 920 -4320
rect 860 -4640 920 -4500
rect 860 -4820 920 -4680
rect -140 -5000 -80 -4860
rect -140 -5180 -80 -5040
rect -140 -5360 -80 -5220
rect 860 -5000 920 -4860
rect 860 -5180 920 -5040
rect 860 -5400 920 -5220
rect -4440 -5460 -4120 -5400
rect -4080 -5460 -3860 -5400
rect -3820 -5460 -3600 -5400
rect -3560 -5460 -3340 -5400
rect -3300 -5460 -3080 -5400
rect -3040 -5460 -2820 -5400
rect -2780 -5460 -2560 -5400
rect -2520 -5460 -2300 -5400
rect -2260 -5460 -2040 -5400
rect -2000 -5460 -1500 -5400
rect -1460 -5460 -1240 -5400
rect -1200 -5460 -980 -5400
rect -940 -5460 -720 -5400
rect -680 -5460 -460 -5400
rect -420 -5460 -200 -5400
rect -160 -5460 60 -5400
rect 100 -5460 320 -5400
rect 360 -5460 580 -5400
rect 620 -5460 920 -5400
<< locali >>
rect -4492 -4120 1008 -4106
rect -4492 -4180 -4480 -4120
rect -4420 -4140 -4380 -4120
rect -4320 -4180 -4280 -4120
rect -4220 -4180 -4180 -4120
rect -4120 -4180 -4080 -4120
rect -4020 -4180 -3980 -4120
rect -3920 -4180 -3880 -4120
rect -3820 -4180 -3780 -4120
rect -3720 -4180 -3680 -4120
rect -3620 -4180 -3580 -4120
rect -3520 -4180 -3480 -4120
rect -3420 -4140 -3380 -4120
rect -3320 -4180 -3280 -4120
rect -3220 -4180 -3180 -4120
rect -3120 -4180 -3080 -4120
rect -3020 -4180 -2980 -4120
rect -2920 -4180 -2880 -4120
rect -2820 -4180 -2780 -4120
rect -2720 -4180 -2680 -4120
rect -2620 -4180 -2580 -4120
rect -2520 -4180 -2480 -4120
rect -2420 -4180 -2380 -4120
rect -2320 -4180 -2280 -4120
rect -2220 -4180 -2180 -4120
rect -2120 -4180 -2080 -4120
rect -2020 -4180 -1980 -4120
rect -1920 -4180 -1880 -4120
rect -1820 -4140 -1780 -4120
rect -1720 -4140 -1680 -4120
rect -1620 -4180 -1580 -4120
rect -1520 -4180 -1480 -4120
rect -1420 -4180 -1380 -4120
rect -1320 -4180 -1280 -4120
rect -1220 -4180 -1180 -4120
rect -1120 -4180 -1080 -4120
rect -1020 -4180 -980 -4120
rect -920 -4180 -880 -4120
rect -820 -4180 -780 -4120
rect -720 -4180 -680 -4120
rect -620 -4180 -580 -4120
rect -520 -4180 -480 -4120
rect -420 -4180 -380 -4120
rect -320 -4180 -280 -4120
rect -220 -4180 -180 -4120
rect -120 -4140 -80 -4120
rect -20 -4180 20 -4120
rect 80 -4180 120 -4120
rect 180 -4180 220 -4120
rect 280 -4180 320 -4120
rect 380 -4180 420 -4120
rect 480 -4180 520 -4120
rect 580 -4180 620 -4120
rect 680 -4180 720 -4120
rect 780 -4180 820 -4120
rect 880 -4140 920 -4120
rect 980 -4180 1008 -4120
rect -4492 -4220 -4440 -4180
rect -4380 -4220 -3440 -4180
rect -3380 -4220 -1820 -4180
rect -1680 -4220 -140 -4180
rect -80 -4220 860 -4180
rect 920 -4220 1008 -4180
rect -4492 -4280 -4480 -4220
rect -4100 -4280 -4080 -4220
rect -3820 -4280 -3800 -4220
rect -3300 -4280 -3280 -4220
rect -3020 -4280 -2980 -4220
rect -2500 -4280 -2480 -4220
rect -2220 -4280 -2200 -4220
rect -1200 -4280 -1180 -4220
rect -920 -4280 -900 -4220
rect -420 -4280 -380 -4220
rect 300 -4280 320 -4220
rect 480 -4280 520 -4220
rect 680 -4280 700 -4220
rect 980 -4280 1008 -4220
rect -4492 -4306 -4440 -4280
rect -4455 -4460 -4440 -4306
rect -4380 -4306 -1820 -4280
rect -4380 -4460 -4349 -4306
rect -4455 -4500 -4349 -4460
rect -4455 -4640 -4440 -4500
rect -4380 -4640 -4349 -4500
rect -4455 -4680 -4349 -4640
rect -4455 -4696 -4440 -4680
rect -4452 -4820 -4440 -4696
rect -4380 -4696 -4349 -4680
rect -4380 -4820 -4352 -4696
rect -4452 -4860 -4352 -4820
rect -4452 -5000 -4440 -4860
rect -4380 -5000 -4352 -4860
rect -4452 -5040 -4352 -5000
rect -4452 -5180 -4440 -5040
rect -4380 -5180 -4352 -5040
rect -3940 -5180 -3820 -4306
rect -3454 -4320 -3348 -4306
rect -3454 -4460 -3440 -4320
rect -3380 -4460 -3348 -4320
rect -3454 -4500 -3348 -4460
rect -3454 -4640 -3440 -4500
rect -3380 -4640 -3348 -4500
rect -3454 -4680 -3348 -4640
rect -3454 -4707 -3440 -4680
rect -3452 -4820 -3440 -4707
rect -3380 -4707 -3348 -4680
rect -3380 -4820 -3352 -4707
rect -3452 -4860 -3352 -4820
rect -3452 -5000 -3440 -4860
rect -3380 -5000 -3352 -4860
rect -3452 -5040 -3352 -5000
rect -3452 -5180 -3440 -5040
rect -3380 -5180 -3352 -5040
rect -3000 -5180 -2880 -4306
rect -2360 -5180 -2240 -4306
rect -1859 -4420 -1820 -4306
rect -1680 -4306 1008 -4280
rect -1680 -4386 -1653 -4306
rect -1680 -4420 -1652 -4386
rect -1859 -4460 -1652 -4420
rect -1859 -4740 -1820 -4460
rect -1680 -4740 -1652 -4460
rect -1859 -4780 -1652 -4740
rect -1859 -4829 -1820 -4780
rect -1852 -5060 -1820 -4829
rect -1680 -5060 -1652 -4780
rect -1852 -5100 -1652 -5060
rect -4452 -5220 -4352 -5180
rect -4452 -5460 -4440 -5220
rect -4380 -5386 -4352 -5220
rect -3452 -5220 -3352 -5180
rect -3452 -5360 -3440 -5220
rect -3380 -5360 -3352 -5220
rect -3452 -5386 -3352 -5360
rect -1852 -5386 -1820 -5100
rect -4380 -5400 -1820 -5386
rect -1680 -5386 -1652 -5100
rect -1260 -5180 -1140 -4306
rect -600 -5180 -480 -4306
rect -151 -4320 -47 -4306
rect -151 -4386 -140 -4320
rect -152 -4460 -140 -4386
rect -80 -4460 -47 -4320
rect -152 -4500 -47 -4460
rect -152 -4640 -140 -4500
rect -80 -4640 -47 -4500
rect -152 -4680 -47 -4640
rect -152 -4820 -140 -4680
rect -80 -4820 -47 -4680
rect -152 -4857 -47 -4820
rect -152 -4860 -52 -4857
rect -152 -5000 -140 -4860
rect -80 -5000 -52 -4860
rect -152 -5040 -52 -5000
rect -152 -5180 -140 -5040
rect -80 -5180 -52 -5040
rect 360 -5180 480 -4306
rect 848 -4320 952 -4306
rect 848 -4460 860 -4320
rect 920 -4460 952 -4320
rect 848 -4500 952 -4460
rect 848 -4640 860 -4500
rect 920 -4640 952 -4500
rect 848 -4680 952 -4640
rect 848 -4820 860 -4680
rect 920 -4820 952 -4680
rect 848 -4835 952 -4820
rect 848 -4860 948 -4835
rect 848 -5000 860 -4860
rect 920 -5000 948 -4860
rect 848 -5040 948 -5000
rect 848 -5180 860 -5040
rect 920 -5180 948 -5040
rect -152 -5220 -52 -5180
rect -152 -5360 -140 -5220
rect -80 -5360 -52 -5220
rect -152 -5386 -52 -5360
rect 848 -5220 948 -5180
rect 848 -5386 860 -5220
rect -1680 -5400 860 -5386
rect -4120 -5460 -4080 -5400
rect -3860 -5460 -3820 -5400
rect -3600 -5460 -3560 -5400
rect -3340 -5460 -3300 -5400
rect -3080 -5460 -3040 -5400
rect -2820 -5460 -2780 -5400
rect -2560 -5460 -2520 -5400
rect -2300 -5460 -2260 -5400
rect -2040 -5460 -2000 -5400
rect -1500 -5460 -1460 -5400
rect -1240 -5460 -1200 -5400
rect -980 -5460 -940 -5400
rect -720 -5460 -680 -5400
rect -460 -5460 -420 -5400
rect -200 -5460 -160 -5400
rect 60 -5460 100 -5400
rect 320 -5460 360 -5400
rect 580 -5460 620 -5400
rect 920 -5460 948 -5220
rect -4452 -5486 948 -5460
rect -2700 -5720 -800 -5700
rect -2700 -5780 -2580 -5720
rect -2440 -5780 -2400 -5720
rect -2260 -5780 -2220 -5720
rect -2080 -5780 -2040 -5720
rect -1900 -5780 -1860 -5720
rect -1720 -5780 -1680 -5720
rect -1540 -5780 -1500 -5720
rect -1360 -5780 -1320 -5720
rect -1180 -5780 -1140 -5720
rect -1000 -5780 -960 -5720
rect -840 -5780 -800 -5720
rect -2700 -5800 -800 -5780
rect -2700 -5900 -2600 -5800
rect -2700 -6040 -2680 -5900
rect -2620 -6040 -2600 -5900
rect -2700 -6080 -2600 -6040
rect -2700 -6220 -2680 -6080
rect -2620 -6220 -2600 -6080
rect -2700 -6260 -2600 -6220
rect -2700 -6400 -2680 -6260
rect -2620 -6400 -2600 -6260
rect -2700 -6440 -2600 -6400
rect -2700 -6580 -2680 -6440
rect -2620 -6580 -2600 -6440
rect -2700 -6600 -2600 -6580
rect -900 -5900 -800 -5800
rect -900 -6040 -880 -5900
rect -820 -6040 -800 -5900
rect -900 -6080 -800 -6040
rect -900 -6220 -880 -6080
rect -820 -6220 -800 -6080
rect -900 -6260 -800 -6220
rect -900 -6400 -880 -6260
rect -820 -6400 -800 -6260
rect -900 -6440 -800 -6400
rect -900 -6580 -880 -6440
rect -820 -6580 -800 -6440
rect -900 -6600 -800 -6580
rect -3700 -6620 200 -6600
rect -3700 -6680 -3600 -6620
rect -3240 -6680 -3200 -6620
rect -3060 -6680 -3020 -6620
rect -2880 -6680 -2840 -6620
rect -2700 -6680 -2660 -6620
rect -2520 -6680 -2480 -6620
rect -2340 -6680 -2300 -6620
rect -2160 -6680 -2120 -6620
rect -1980 -6680 -1940 -6620
rect -1800 -6680 -1760 -6620
rect -1620 -6680 -1580 -6620
rect -1440 -6680 -1400 -6620
rect -1260 -6680 -1220 -6620
rect -1080 -6680 -1040 -6620
rect -900 -6680 -860 -6620
rect -720 -6680 -680 -6620
rect -540 -6680 -500 -6620
rect -360 -6680 -320 -6620
rect -180 -6680 -140 -6620
rect 100 -6680 200 -6620
rect -3700 -6700 200 -6680
rect -3700 -6760 -3600 -6700
rect -3700 -6900 -3680 -6760
rect -3620 -6900 -3600 -6760
rect -3700 -6940 -3600 -6900
rect -3700 -7080 -3680 -6940
rect -3620 -7080 -3600 -6940
rect -2700 -6740 -2600 -6700
rect -2700 -6880 -2680 -6740
rect -2620 -6880 -2600 -6740
rect -2700 -6920 -2600 -6880
rect -3700 -7120 -3600 -7080
rect -3700 -7260 -3680 -7120
rect -3620 -7260 -3600 -7120
rect -3700 -7300 -3600 -7260
rect -3700 -7440 -3680 -7300
rect -3620 -7440 -3600 -7300
rect -3700 -7480 -3600 -7440
rect -3700 -7620 -3680 -7480
rect -3620 -7620 -3600 -7480
rect -3700 -7660 -3600 -7620
rect -3700 -7800 -3680 -7660
rect -4500 -7820 -3680 -7800
rect -3620 -7800 -3600 -7660
rect -3160 -7800 -3040 -7000
rect -2700 -7060 -2680 -6920
rect -2620 -7060 -2600 -6920
rect -2700 -7100 -2600 -7060
rect -2700 -7240 -2680 -7100
rect -2620 -7240 -2600 -7100
rect -2700 -7280 -2600 -7240
rect -2700 -7420 -2680 -7280
rect -2620 -7420 -2600 -7280
rect -2700 -7460 -2600 -7420
rect -2700 -7600 -2680 -7460
rect -2620 -7600 -2600 -7460
rect -2700 -7640 -2600 -7600
rect -2700 -7780 -2680 -7640
rect -2620 -7780 -2600 -7640
rect -2700 -7800 -2600 -7780
rect -900 -6740 -800 -6700
rect -900 -6880 -880 -6740
rect -820 -6880 -800 -6740
rect -900 -6920 -800 -6880
rect -900 -7060 -880 -6920
rect -820 -7060 -800 -6920
rect 100 -6760 200 -6700
rect 100 -6900 120 -6760
rect 180 -6900 200 -6760
rect 100 -6940 200 -6900
rect -900 -7100 -800 -7060
rect -900 -7240 -880 -7100
rect -820 -7240 -800 -7100
rect -900 -7280 -800 -7240
rect -900 -7420 -880 -7280
rect -820 -7420 -800 -7280
rect -900 -7460 -800 -7420
rect -900 -7600 -880 -7460
rect -820 -7600 -800 -7460
rect -900 -7640 -800 -7600
rect -900 -7780 -880 -7640
rect -820 -7780 -800 -7640
rect -900 -7800 -800 -7780
rect -360 -7800 -240 -7000
rect 100 -7080 120 -6940
rect 180 -7080 200 -6940
rect 100 -7120 200 -7080
rect 100 -7260 120 -7120
rect 180 -7260 200 -7120
rect 100 -7300 200 -7260
rect 100 -7440 120 -7300
rect 180 -7440 200 -7300
rect 100 -7480 200 -7440
rect 100 -7620 120 -7480
rect 180 -7620 200 -7480
rect 100 -7660 200 -7620
rect 100 -7800 120 -7660
rect -3620 -7820 120 -7800
rect 180 -7800 200 -7660
rect 180 -7820 1000 -7800
rect -4500 -7880 -4480 -7820
rect -4420 -7880 -4380 -7820
rect -4320 -7880 -4280 -7820
rect -4220 -7880 -4180 -7820
rect -4120 -7880 -4080 -7820
rect -4020 -7880 -3980 -7820
rect -3920 -7880 -3880 -7820
rect -3820 -7880 -3780 -7820
rect -3720 -7880 -3680 -7820
rect -3420 -7880 -3380 -7820
rect -3220 -7880 -3200 -7820
rect -2700 -7880 -2680 -7820
rect -2520 -7880 -2480 -7820
rect -2320 -7880 -2300 -7820
rect -1800 -7880 -1780 -7820
rect -1620 -7880 -1580 -7820
rect -1420 -7880 -1400 -7820
rect -900 -7880 -880 -7820
rect -720 -7880 -680 -7820
rect -520 -7880 -500 -7820
rect 180 -7880 220 -7820
rect 280 -7880 320 -7820
rect 380 -7880 420 -7820
rect 480 -7880 520 -7820
rect 580 -7880 620 -7820
rect 680 -7880 720 -7820
rect 780 -7880 820 -7820
rect 880 -7880 920 -7820
rect 980 -7880 1000 -7820
rect -4500 -7920 1000 -7880
rect -4500 -7980 -4480 -7920
rect -4420 -7980 -4380 -7920
rect -4320 -7980 -4280 -7920
rect -4220 -7980 -4180 -7920
rect -4120 -7980 -4080 -7920
rect -4020 -7980 -3980 -7920
rect -3920 -7980 -3880 -7920
rect -3820 -7980 -3780 -7920
rect -3720 -7980 -3680 -7920
rect -3620 -7980 -3580 -7920
rect -3520 -7980 -3480 -7920
rect -3420 -7980 -3380 -7920
rect -3320 -7980 -3280 -7920
rect -3220 -7980 -3180 -7920
rect -3120 -7980 -3080 -7920
rect -3020 -7980 -2980 -7920
rect -2920 -7980 -2880 -7920
rect -2820 -7980 -2780 -7920
rect -2720 -7980 -2680 -7920
rect -2620 -7980 -2580 -7920
rect -2520 -7980 -2480 -7920
rect -2420 -7980 -2380 -7920
rect -2320 -7980 -2280 -7920
rect -2220 -7980 -2180 -7920
rect -2120 -7980 -2080 -7920
rect -2020 -7980 -1980 -7920
rect -1920 -7980 -1880 -7920
rect -1820 -7980 -1780 -7920
rect -1720 -7980 -1680 -7920
rect -1620 -7980 -1580 -7920
rect -1520 -7980 -1480 -7920
rect -1420 -7980 -1380 -7920
rect -1320 -7980 -1280 -7920
rect -1220 -7980 -1180 -7920
rect -1120 -7980 -1080 -7920
rect -1020 -7980 -980 -7920
rect -920 -7980 -880 -7920
rect -820 -7980 -780 -7920
rect -720 -7980 -680 -7920
rect -620 -7980 -580 -7920
rect -520 -7980 -480 -7920
rect -420 -7980 -380 -7920
rect -320 -7980 -280 -7920
rect -220 -7980 -180 -7920
rect -120 -7980 -80 -7920
rect -20 -7980 20 -7920
rect 80 -7980 120 -7920
rect 180 -7980 220 -7920
rect 280 -7980 320 -7920
rect 380 -7980 420 -7920
rect 480 -7980 520 -7920
rect 580 -7980 620 -7920
rect 680 -7980 720 -7920
rect 780 -7980 820 -7920
rect 880 -7980 920 -7920
rect 980 -7980 1000 -7920
rect -4500 -8000 1000 -7980
<< viali >>
rect -4480 -4140 -4420 -4120
rect -4480 -4180 -4440 -4140
rect -4440 -4180 -4420 -4140
rect -4380 -4180 -4320 -4120
rect -4280 -4180 -4220 -4120
rect -4180 -4180 -4120 -4120
rect -4080 -4180 -4020 -4120
rect -3980 -4180 -3920 -4120
rect -3880 -4180 -3820 -4120
rect -3780 -4180 -3720 -4120
rect -3680 -4180 -3620 -4120
rect -3580 -4180 -3520 -4120
rect -3480 -4140 -3420 -4120
rect -3480 -4180 -3440 -4140
rect -3440 -4180 -3420 -4140
rect -3380 -4180 -3320 -4120
rect -3280 -4180 -3220 -4120
rect -3180 -4180 -3120 -4120
rect -3080 -4180 -3020 -4120
rect -2980 -4180 -2920 -4120
rect -2880 -4180 -2820 -4120
rect -2780 -4180 -2720 -4120
rect -2680 -4180 -2620 -4120
rect -2580 -4180 -2520 -4120
rect -2480 -4180 -2420 -4120
rect -2380 -4180 -2320 -4120
rect -2280 -4180 -2220 -4120
rect -2180 -4180 -2120 -4120
rect -2080 -4180 -2020 -4120
rect -1980 -4180 -1920 -4120
rect -1880 -4180 -1820 -4120
rect -1780 -4140 -1720 -4120
rect -1780 -4180 -1720 -4140
rect -1680 -4180 -1620 -4120
rect -1580 -4180 -1520 -4120
rect -1480 -4180 -1420 -4120
rect -1380 -4180 -1320 -4120
rect -1280 -4180 -1220 -4120
rect -1180 -4180 -1120 -4120
rect -1080 -4180 -1020 -4120
rect -980 -4180 -920 -4120
rect -880 -4180 -820 -4120
rect -780 -4180 -720 -4120
rect -680 -4180 -620 -4120
rect -580 -4180 -520 -4120
rect -480 -4180 -420 -4120
rect -380 -4180 -320 -4120
rect -280 -4180 -220 -4120
rect -180 -4140 -120 -4120
rect -180 -4180 -140 -4140
rect -140 -4180 -120 -4140
rect -80 -4180 -20 -4120
rect 20 -4180 80 -4120
rect 120 -4180 180 -4120
rect 220 -4180 280 -4120
rect 320 -4180 380 -4120
rect 420 -4180 480 -4120
rect 520 -4180 580 -4120
rect 620 -4180 680 -4120
rect 720 -4180 780 -4120
rect 820 -4140 880 -4120
rect 820 -4180 860 -4140
rect 860 -4180 880 -4140
rect 920 -4180 980 -4120
rect -4480 -4280 -4440 -4220
rect -4440 -4280 -4420 -4220
rect -4380 -4280 -4320 -4220
rect -4280 -4280 -4220 -4220
rect -4180 -4280 -4120 -4220
rect -4080 -4280 -4060 -4220
rect -4060 -4280 -4020 -4220
rect -3980 -4280 -3920 -4220
rect -3880 -4280 -3840 -4220
rect -3840 -4280 -3820 -4220
rect -3780 -4280 -3720 -4220
rect -3680 -4280 -3620 -4220
rect -3580 -4280 -3520 -4220
rect -3480 -4280 -3420 -4220
rect -3380 -4280 -3320 -4220
rect -3280 -4280 -3260 -4220
rect -3260 -4280 -3220 -4220
rect -3180 -4280 -3120 -4220
rect -3080 -4280 -3040 -4220
rect -3040 -4280 -3020 -4220
rect -2980 -4280 -2920 -4220
rect -2880 -4280 -2820 -4220
rect -2780 -4280 -2760 -4220
rect -2760 -4280 -2720 -4220
rect -2680 -4280 -2620 -4220
rect -2580 -4280 -2520 -4220
rect -2480 -4280 -2460 -4220
rect -2460 -4280 -2420 -4220
rect -2380 -4280 -2320 -4220
rect -2280 -4280 -2240 -4220
rect -2240 -4280 -2220 -4220
rect -2180 -4280 -2120 -4220
rect -2080 -4280 -2020 -4220
rect -1980 -4280 -1940 -4220
rect -1940 -4280 -1920 -4220
rect -1880 -4280 -1820 -4220
rect -1780 -4280 -1720 -4220
rect -1680 -4280 -1620 -4220
rect -1580 -4280 -1520 -4220
rect -1480 -4280 -1460 -4220
rect -1460 -4280 -1420 -4220
rect -1380 -4280 -1320 -4220
rect -1280 -4280 -1220 -4220
rect -1180 -4280 -1160 -4220
rect -1160 -4280 -1120 -4220
rect -1080 -4280 -1020 -4220
rect -980 -4280 -940 -4220
rect -940 -4280 -920 -4220
rect -880 -4280 -820 -4220
rect -780 -4280 -720 -4220
rect -680 -4280 -640 -4220
rect -640 -4280 -620 -4220
rect -580 -4280 -520 -4220
rect -480 -4280 -420 -4220
rect -380 -4280 -340 -4220
rect -340 -4280 -320 -4220
rect -280 -4280 -220 -4220
rect -180 -4280 -120 -4220
rect -80 -4280 -20 -4220
rect 20 -4280 80 -4220
rect 120 -4280 160 -4220
rect 160 -4280 180 -4220
rect 220 -4280 280 -4220
rect 320 -4280 340 -4220
rect 340 -4280 380 -4220
rect 420 -4280 480 -4220
rect 520 -4280 580 -4220
rect 620 -4280 660 -4220
rect 660 -4280 680 -4220
rect 720 -4280 780 -4220
rect 820 -4280 880 -4220
rect 920 -4280 980 -4220
rect -4480 -7880 -4420 -7820
rect -4380 -7880 -4320 -7820
rect -4280 -7880 -4220 -7820
rect -4180 -7880 -4120 -7820
rect -4080 -7880 -4020 -7820
rect -3980 -7880 -3920 -7820
rect -3880 -7880 -3820 -7820
rect -3780 -7880 -3720 -7820
rect -3680 -7880 -3620 -7820
rect -3580 -7880 -3520 -7820
rect -3480 -7880 -3420 -7820
rect -3380 -7880 -3320 -7820
rect -3280 -7880 -3240 -7820
rect -3240 -7880 -3220 -7820
rect -3180 -7880 -3120 -7820
rect -3080 -7880 -3060 -7820
rect -3060 -7880 -3020 -7820
rect -2980 -7880 -2920 -7820
rect -2880 -7880 -2840 -7820
rect -2840 -7880 -2820 -7820
rect -2780 -7880 -2720 -7820
rect -2680 -7880 -2660 -7820
rect -2660 -7880 -2620 -7820
rect -2580 -7880 -2520 -7820
rect -2480 -7880 -2420 -7820
rect -2380 -7880 -2340 -7820
rect -2340 -7880 -2320 -7820
rect -2280 -7880 -2220 -7820
rect -2180 -7880 -2160 -7820
rect -2160 -7880 -2120 -7820
rect -2080 -7880 -2020 -7820
rect -1980 -7880 -1940 -7820
rect -1940 -7880 -1920 -7820
rect -1880 -7880 -1820 -7820
rect -1780 -7880 -1760 -7820
rect -1760 -7880 -1720 -7820
rect -1680 -7880 -1620 -7820
rect -1580 -7880 -1520 -7820
rect -1480 -7880 -1440 -7820
rect -1440 -7880 -1420 -7820
rect -1380 -7880 -1320 -7820
rect -1280 -7880 -1260 -7820
rect -1260 -7880 -1220 -7820
rect -1180 -7880 -1120 -7820
rect -1080 -7880 -1040 -7820
rect -1040 -7880 -1020 -7820
rect -980 -7880 -920 -7820
rect -880 -7880 -860 -7820
rect -860 -7880 -820 -7820
rect -780 -7880 -720 -7820
rect -680 -7880 -620 -7820
rect -580 -7880 -540 -7820
rect -540 -7880 -520 -7820
rect -480 -7880 -420 -7820
rect -380 -7880 -360 -7820
rect -360 -7880 -320 -7820
rect -280 -7880 -220 -7820
rect -180 -7880 -140 -7820
rect -140 -7880 -120 -7820
rect -80 -7880 -20 -7820
rect 20 -7880 80 -7820
rect 120 -7880 180 -7820
rect 220 -7880 280 -7820
rect 320 -7880 380 -7820
rect 420 -7880 480 -7820
rect 520 -7880 580 -7820
rect 620 -7880 680 -7820
rect 720 -7880 780 -7820
rect 820 -7880 880 -7820
rect 920 -7880 980 -7820
rect -4480 -7980 -4420 -7920
rect -4380 -7980 -4320 -7920
rect -4280 -7980 -4220 -7920
rect -4180 -7980 -4120 -7920
rect -4080 -7980 -4020 -7920
rect -3980 -7980 -3920 -7920
rect -3880 -7980 -3820 -7920
rect -3780 -7980 -3720 -7920
rect -3680 -7980 -3620 -7920
rect -3580 -7980 -3520 -7920
rect -3480 -7980 -3420 -7920
rect -3380 -7980 -3320 -7920
rect -3280 -7980 -3220 -7920
rect -3180 -7980 -3120 -7920
rect -3080 -7980 -3020 -7920
rect -2980 -7980 -2920 -7920
rect -2880 -7980 -2820 -7920
rect -2780 -7980 -2720 -7920
rect -2680 -7980 -2620 -7920
rect -2580 -7980 -2520 -7920
rect -2480 -7980 -2420 -7920
rect -2380 -7980 -2320 -7920
rect -2280 -7980 -2220 -7920
rect -2180 -7980 -2120 -7920
rect -2080 -7980 -2020 -7920
rect -1980 -7980 -1920 -7920
rect -1880 -7980 -1820 -7920
rect -1780 -7980 -1720 -7920
rect -1680 -7980 -1620 -7920
rect -1580 -7980 -1520 -7920
rect -1480 -7980 -1420 -7920
rect -1380 -7980 -1320 -7920
rect -1280 -7980 -1220 -7920
rect -1180 -7980 -1120 -7920
rect -1080 -7980 -1020 -7920
rect -980 -7980 -920 -7920
rect -880 -7980 -820 -7920
rect -780 -7980 -720 -7920
rect -680 -7980 -620 -7920
rect -580 -7980 -520 -7920
rect -480 -7980 -420 -7920
rect -380 -7980 -320 -7920
rect -280 -7980 -220 -7920
rect -180 -7980 -120 -7920
rect -80 -7980 -20 -7920
rect 20 -7980 80 -7920
rect 120 -7980 180 -7920
rect 220 -7980 280 -7920
rect 320 -7980 380 -7920
rect 420 -7980 480 -7920
rect 520 -7980 580 -7920
rect 620 -7980 680 -7920
rect 720 -7980 780 -7920
rect 820 -7980 880 -7920
rect 920 -7980 980 -7920
<< metal1 >>
rect -4492 -4120 1008 -4106
rect -4492 -4180 -4480 -4120
rect -4420 -4180 -4380 -4120
rect -4320 -4180 -4280 -4120
rect -4220 -4180 -4180 -4120
rect -4120 -4180 -4080 -4120
rect -4020 -4180 -3980 -4120
rect -3920 -4180 -3880 -4120
rect -3820 -4180 -3780 -4120
rect -3720 -4180 -3680 -4120
rect -3620 -4180 -3580 -4120
rect -3520 -4180 -3480 -4120
rect -3420 -4180 -3380 -4120
rect -3320 -4180 -3280 -4120
rect -3220 -4180 -3180 -4120
rect -3120 -4180 -3080 -4120
rect -3020 -4180 -2980 -4120
rect -2920 -4180 -2880 -4120
rect -2820 -4180 -2780 -4120
rect -2720 -4180 -2680 -4120
rect -2620 -4180 -2580 -4120
rect -2520 -4180 -2480 -4120
rect -2420 -4180 -2380 -4120
rect -2320 -4180 -2280 -4120
rect -2220 -4180 -2180 -4120
rect -2120 -4180 -2080 -4120
rect -2020 -4180 -1980 -4120
rect -1920 -4180 -1880 -4120
rect -1820 -4180 -1780 -4120
rect -1720 -4180 -1680 -4120
rect -1620 -4180 -1580 -4120
rect -1520 -4180 -1480 -4120
rect -1420 -4180 -1380 -4120
rect -1320 -4180 -1280 -4120
rect -1220 -4180 -1180 -4120
rect -1120 -4180 -1080 -4120
rect -1020 -4180 -980 -4120
rect -920 -4180 -880 -4120
rect -820 -4180 -780 -4120
rect -720 -4180 -680 -4120
rect -620 -4180 -580 -4120
rect -520 -4180 -480 -4120
rect -420 -4180 -380 -4120
rect -320 -4180 -280 -4120
rect -220 -4180 -180 -4120
rect -120 -4180 -80 -4120
rect -20 -4180 20 -4120
rect 80 -4180 120 -4120
rect 180 -4180 220 -4120
rect 280 -4180 320 -4120
rect 380 -4180 420 -4120
rect 480 -4180 520 -4120
rect 580 -4180 620 -4120
rect 680 -4180 720 -4120
rect 780 -4180 820 -4120
rect 880 -4180 920 -4120
rect 980 -4180 1008 -4120
rect -4492 -4220 1008 -4180
rect -4492 -4280 -4480 -4220
rect -4420 -4280 -4380 -4220
rect -4320 -4280 -4280 -4220
rect -4220 -4280 -4180 -4220
rect -4120 -4280 -4080 -4220
rect -4020 -4280 -3980 -4220
rect -3920 -4280 -3880 -4220
rect -3820 -4280 -3780 -4220
rect -3720 -4280 -3680 -4220
rect -3620 -4280 -3580 -4220
rect -3520 -4280 -3480 -4220
rect -3420 -4280 -3380 -4220
rect -3320 -4280 -3280 -4220
rect -3220 -4280 -3180 -4220
rect -3120 -4280 -3080 -4220
rect -3020 -4280 -2980 -4220
rect -2920 -4280 -2880 -4220
rect -2820 -4280 -2780 -4220
rect -2720 -4280 -2680 -4220
rect -2620 -4280 -2580 -4220
rect -2520 -4280 -2480 -4220
rect -2420 -4280 -2380 -4220
rect -2320 -4280 -2280 -4220
rect -2220 -4280 -2180 -4220
rect -2120 -4280 -2080 -4220
rect -2020 -4280 -1980 -4220
rect -1920 -4280 -1880 -4220
rect -1820 -4280 -1780 -4220
rect -1720 -4280 -1680 -4220
rect -1620 -4280 -1580 -4220
rect -1520 -4280 -1480 -4220
rect -1420 -4280 -1380 -4220
rect -1320 -4280 -1280 -4220
rect -1220 -4280 -1180 -4220
rect -1120 -4280 -1080 -4220
rect -1020 -4280 -980 -4220
rect -920 -4280 -880 -4220
rect -820 -4280 -780 -4220
rect -720 -4280 -680 -4220
rect -620 -4280 -580 -4220
rect -520 -4280 -480 -4220
rect -420 -4280 -380 -4220
rect -320 -4280 -280 -4220
rect -220 -4280 -180 -4220
rect -120 -4280 -80 -4220
rect -20 -4280 20 -4220
rect 80 -4280 120 -4220
rect 180 -4280 220 -4220
rect 280 -4280 320 -4220
rect 380 -4280 420 -4220
rect 480 -4280 520 -4220
rect 580 -4280 620 -4220
rect 680 -4280 720 -4220
rect 780 -4280 820 -4220
rect 880 -4280 920 -4220
rect 980 -4280 1008 -4220
rect -4492 -4306 1008 -4280
rect -4260 -4500 -4140 -4420
rect -4260 -4560 -4240 -4500
rect -4180 -4560 -4140 -4500
rect -4260 -4600 -4140 -4560
rect -4260 -4660 -4240 -4600
rect -4180 -4660 -4140 -4600
rect -4260 -4700 -4140 -4660
rect -4260 -4760 -4240 -4700
rect -4180 -4760 -4140 -4700
rect -4260 -4800 -4140 -4760
rect -4260 -4860 -4240 -4800
rect -4180 -4860 -4140 -4800
rect -4260 -4900 -4140 -4860
rect -4260 -4960 -4240 -4900
rect -4180 -4960 -4140 -4900
rect -4260 -5000 -4140 -4960
rect -4260 -5060 -4240 -5000
rect -4180 -5060 -4140 -5000
rect -4260 -5100 -4140 -5060
rect -4260 -5160 -4240 -5100
rect -4180 -5160 -4140 -5100
rect -4260 -5180 -4140 -5160
rect -3660 -4500 -3540 -4420
rect -3660 -4560 -3620 -4500
rect -3560 -4560 -3540 -4500
rect -3660 -4600 -3540 -4560
rect -3660 -4660 -3620 -4600
rect -3560 -4660 -3540 -4600
rect -3660 -4700 -3540 -4660
rect -3660 -4760 -3620 -4700
rect -3560 -4760 -3540 -4700
rect -3660 -4800 -3540 -4760
rect -3660 -4860 -3620 -4800
rect -3560 -4860 -3540 -4800
rect -3660 -4900 -3540 -4860
rect -3660 -4960 -3620 -4900
rect -3560 -4960 -3540 -4900
rect -3660 -5000 -3540 -4960
rect -3660 -5060 -3620 -5000
rect -3560 -5060 -3540 -5000
rect -3660 -5100 -3540 -5060
rect -3660 -5160 -3620 -5100
rect -3560 -5160 -3540 -5100
rect -3660 -5180 -3540 -5160
rect -3320 -4500 -3200 -4420
rect -3320 -4560 -3300 -4500
rect -3240 -4560 -3200 -4500
rect -3320 -4600 -3200 -4560
rect -3320 -4660 -3300 -4600
rect -3240 -4660 -3200 -4600
rect -3320 -4700 -3200 -4660
rect -3320 -4760 -3300 -4700
rect -3240 -4760 -3200 -4700
rect -2680 -4760 -2560 -4460
rect -3320 -4800 -3200 -4760
rect -3320 -4860 -3300 -4800
rect -3240 -4860 -3200 -4800
rect -3320 -4900 -3200 -4860
rect -3320 -4960 -3300 -4900
rect -3240 -4960 -3200 -4900
rect -3320 -5000 -3200 -4960
rect -3320 -5060 -3300 -5000
rect -3240 -5060 -3200 -5000
rect -3320 -5100 -3200 -5060
rect -3320 -5160 -3300 -5100
rect -3240 -5160 -3200 -5100
rect -3320 -5180 -3200 -5160
rect -2700 -5220 -2560 -4760
rect -2060 -4500 -1940 -4420
rect -2060 -4560 -2020 -4500
rect -1960 -4560 -1940 -4500
rect -2060 -4600 -1940 -4560
rect -2060 -4660 -2020 -4600
rect -1960 -4660 -1940 -4600
rect -2060 -4700 -1940 -4660
rect -2060 -4760 -2020 -4700
rect -1960 -4760 -1940 -4700
rect -2060 -4800 -1940 -4760
rect -2060 -4860 -2020 -4800
rect -1960 -4860 -1940 -4800
rect -2060 -4900 -1940 -4860
rect -2060 -4960 -2020 -4900
rect -1960 -4960 -1940 -4900
rect -2060 -5000 -1940 -4960
rect -2060 -5060 -2020 -5000
rect -1960 -5060 -1940 -5000
rect -2060 -5100 -1940 -5060
rect -2060 -5160 -2020 -5100
rect -1960 -5160 -1940 -5100
rect -2060 -5180 -1940 -5160
rect -1560 -4500 -1440 -4420
rect -1560 -4560 -1540 -4500
rect -1480 -4560 -1440 -4500
rect -1560 -4600 -1440 -4560
rect -1560 -4660 -1540 -4600
rect -1480 -4660 -1440 -4600
rect -1560 -4700 -1440 -4660
rect -1560 -4760 -1540 -4700
rect -1480 -4760 -1440 -4700
rect -1560 -4800 -1440 -4760
rect -1560 -4860 -1540 -4800
rect -1480 -4860 -1440 -4800
rect -1560 -4900 -1440 -4860
rect -1560 -4960 -1540 -4900
rect -1480 -4960 -1440 -4900
rect -1560 -5000 -1440 -4960
rect -1560 -5060 -1540 -5000
rect -1480 -5060 -1440 -5000
rect -1560 -5100 -1440 -5060
rect -1560 -5160 -1540 -5100
rect -1480 -5160 -1440 -5100
rect -1560 -5180 -1440 -5160
rect -920 -5220 -800 -4440
rect -300 -4500 -180 -4420
rect -300 -4560 -260 -4500
rect -200 -4560 -180 -4500
rect -300 -4600 -180 -4560
rect -300 -4660 -260 -4600
rect -200 -4660 -180 -4600
rect -300 -4700 -180 -4660
rect -300 -4760 -260 -4700
rect -200 -4760 -180 -4700
rect -300 -4800 -180 -4760
rect -300 -4860 -260 -4800
rect -200 -4860 -180 -4800
rect -300 -4900 -180 -4860
rect -300 -4960 -260 -4900
rect -200 -4960 -180 -4900
rect -300 -5000 -180 -4960
rect -300 -5060 -260 -5000
rect -200 -5060 -180 -5000
rect -300 -5100 -180 -5060
rect -300 -5160 -260 -5100
rect -200 -5160 -180 -5100
rect -300 -5180 -180 -5160
rect 40 -4500 160 -4420
rect 40 -4560 60 -4500
rect 120 -4560 160 -4500
rect 40 -4600 160 -4560
rect 40 -4660 60 -4600
rect 120 -4660 160 -4600
rect 40 -4700 160 -4660
rect 40 -4760 60 -4700
rect 120 -4760 160 -4700
rect 40 -4800 160 -4760
rect 40 -4860 60 -4800
rect 120 -4860 160 -4800
rect 40 -4900 160 -4860
rect 40 -4960 60 -4900
rect 120 -4960 160 -4900
rect 40 -5000 160 -4960
rect 40 -5060 60 -5000
rect 120 -5060 160 -5000
rect 40 -5100 160 -5060
rect 40 -5160 60 -5100
rect 120 -5160 160 -5100
rect 40 -5180 160 -5160
rect 660 -4500 780 -4420
rect 660 -4560 700 -4500
rect 760 -4560 780 -4500
rect 660 -4600 780 -4560
rect 660 -4660 700 -4600
rect 760 -4660 780 -4600
rect 660 -4700 780 -4660
rect 660 -4760 700 -4700
rect 760 -4760 780 -4700
rect 660 -4800 780 -4760
rect 660 -4860 700 -4800
rect 760 -4860 780 -4800
rect 660 -4900 780 -4860
rect 660 -4960 700 -4900
rect 760 -4960 780 -4900
rect 660 -5000 780 -4960
rect 660 -5060 700 -5000
rect 760 -5060 780 -5000
rect 660 -5100 780 -5060
rect 660 -5160 700 -5100
rect 760 -5160 780 -5100
rect 660 -5180 780 -5160
rect -4140 -5300 -2020 -5220
rect -1460 -5300 680 -5220
rect -2700 -5760 -2580 -5300
rect -920 -5600 -800 -5300
rect -2060 -5620 -800 -5600
rect -2060 -5680 -2040 -5620
rect -1980 -5680 -1940 -5620
rect -1880 -5680 -1840 -5620
rect -1780 -5680 -800 -5620
rect -2060 -5700 -800 -5680
rect -2700 -5840 -2680 -5760
rect -2600 -5840 -2580 -5760
rect -2700 -5860 -2580 -5840
rect -2320 -5780 -2220 -5740
rect -2320 -5840 -2300 -5780
rect -2240 -5840 -2220 -5780
rect -2320 -5880 -2220 -5840
rect -2320 -5940 -2300 -5880
rect -2240 -5940 -2220 -5880
rect -2320 -5980 -2220 -5940
rect -2320 -6040 -2300 -5980
rect -2240 -6040 -2220 -5980
rect -2320 -6080 -2220 -6040
rect -2320 -6140 -2300 -6080
rect -2240 -6140 -2220 -6080
rect -2320 -6180 -2220 -6140
rect -2320 -6240 -2300 -6180
rect -2240 -6240 -2220 -6180
rect -2320 -6320 -2220 -6240
rect -2460 -6380 -2100 -6360
rect -2460 -6440 -2440 -6380
rect -2380 -6440 -2320 -6380
rect -2260 -6440 -2180 -6380
rect -2120 -6440 -2100 -6380
rect -2460 -6460 -2100 -6440
rect -2060 -6600 -1960 -5920
rect -1780 -6340 -1680 -5700
rect -1240 -5780 -1140 -5740
rect -1240 -5840 -1220 -5780
rect -1160 -5840 -1140 -5780
rect -1240 -5880 -1140 -5840
rect -1920 -6380 -1820 -6360
rect -1920 -6440 -1900 -6380
rect -1840 -6440 -1820 -6380
rect -1920 -6460 -1820 -6440
rect -1640 -6380 -1540 -6360
rect -1640 -6440 -1620 -6380
rect -1560 -6440 -1540 -6380
rect -1640 -6460 -1540 -6440
rect -1500 -6600 -1400 -5920
rect -1240 -5940 -1220 -5880
rect -1160 -5940 -1140 -5880
rect -1240 -5980 -1140 -5940
rect -1240 -6040 -1220 -5980
rect -1160 -6040 -1140 -5980
rect -1240 -6080 -1140 -6040
rect -1240 -6140 -1220 -6080
rect -1160 -6140 -1140 -6080
rect -1240 -6180 -1140 -6140
rect -1240 -6240 -1220 -6180
rect -1160 -6240 -1140 -6180
rect -1240 -6320 -1140 -6240
rect -1360 -6380 -1040 -6360
rect -1360 -6440 -1340 -6380
rect -1280 -6440 -1220 -6380
rect -1160 -6440 -1120 -6380
rect -1060 -6440 -1040 -6380
rect -1360 -6460 -1040 -6440
rect -2060 -6700 -1320 -6600
rect -3320 -6860 -2900 -6840
rect -3320 -6920 -3300 -6860
rect -3240 -6920 -3200 -6860
rect -3140 -6920 -3080 -6860
rect -3020 -6920 -2980 -6860
rect -2920 -6920 -2900 -6860
rect -3320 -6940 -2900 -6920
rect -3480 -7000 -3360 -6980
rect -3480 -7060 -3460 -7000
rect -3400 -7060 -3360 -7000
rect -3480 -7100 -3360 -7060
rect -3480 -7160 -3460 -7100
rect -3400 -7160 -3360 -7100
rect -3480 -7200 -3360 -7160
rect -3480 -7260 -3460 -7200
rect -3400 -7260 -3360 -7200
rect -3480 -7300 -3360 -7260
rect -3480 -7360 -3460 -7300
rect -3400 -7360 -3360 -7300
rect -3480 -7400 -3360 -7360
rect -3480 -7460 -3460 -7400
rect -3400 -7460 -3360 -7400
rect -3480 -7500 -3360 -7460
rect -3480 -7560 -3460 -7500
rect -3400 -7560 -3360 -7500
rect -3480 -7580 -3360 -7560
rect -2860 -7000 -2740 -6980
rect -2860 -7060 -2820 -7000
rect -2760 -7060 -2740 -7000
rect -2860 -7100 -2740 -7060
rect -2860 -7160 -2820 -7100
rect -2760 -7160 -2740 -7100
rect -2860 -7200 -2740 -7160
rect -2860 -7260 -2820 -7200
rect -2760 -7260 -2740 -7200
rect -2860 -7300 -2740 -7260
rect -2860 -7360 -2820 -7300
rect -2760 -7360 -2740 -7300
rect -2860 -7400 -2740 -7360
rect -2860 -7460 -2820 -7400
rect -2760 -7460 -2740 -7400
rect -2860 -7500 -2740 -7460
rect -2860 -7560 -2820 -7500
rect -2760 -7560 -2740 -7500
rect -2860 -7580 -2740 -7560
rect -2060 -7580 -1960 -6700
rect -1920 -7620 -1780 -7520
rect -2180 -7660 -1780 -7620
rect -2180 -7720 -2160 -7660
rect -2100 -7720 -2060 -7660
rect -2000 -7720 -1960 -7660
rect -1900 -7720 -1860 -7660
rect -1800 -7720 -1780 -7660
rect -2180 -7760 -1780 -7720
rect -1740 -7800 -1620 -6900
rect -1580 -7600 -1460 -7520
rect -1420 -7580 -1320 -6700
rect -520 -6860 -80 -6840
rect -520 -6920 -500 -6860
rect -440 -6920 -400 -6860
rect -340 -6920 -260 -6860
rect -200 -6920 -160 -6860
rect -100 -6920 -80 -6860
rect -520 -6940 -80 -6920
rect -700 -7000 -540 -6980
rect -700 -7060 -660 -7000
rect -600 -7060 -540 -7000
rect -700 -7100 -540 -7060
rect -700 -7160 -660 -7100
rect -600 -7160 -540 -7100
rect -700 -7200 -540 -7160
rect -700 -7260 -660 -7200
rect -600 -7260 -540 -7200
rect -700 -7300 -540 -7260
rect -700 -7360 -660 -7300
rect -600 -7360 -540 -7300
rect -700 -7400 -540 -7360
rect -700 -7460 -660 -7400
rect -600 -7460 -540 -7400
rect -700 -7500 -540 -7460
rect -700 -7560 -660 -7500
rect -600 -7560 -540 -7500
rect -700 -7580 -540 -7560
rect -60 -7000 100 -6980
rect -60 -7060 0 -7000
rect 60 -7060 100 -7000
rect -60 -7100 100 -7060
rect -60 -7160 0 -7100
rect 60 -7160 100 -7100
rect -60 -7200 100 -7160
rect -60 -7260 0 -7200
rect 60 -7260 100 -7200
rect -60 -7300 100 -7260
rect -60 -7360 0 -7300
rect 60 -7360 100 -7300
rect -60 -7400 100 -7360
rect -60 -7460 0 -7400
rect 60 -7460 100 -7400
rect -60 -7500 100 -7460
rect -60 -7560 0 -7500
rect 60 -7560 100 -7500
rect -60 -7580 100 -7560
rect -1580 -7620 -1440 -7600
rect -1580 -7660 -1200 -7620
rect -1580 -7720 -1560 -7660
rect -1500 -7720 -1460 -7660
rect -1400 -7720 -1360 -7660
rect -1300 -7720 -1280 -7660
rect -1220 -7720 -1200 -7660
rect -1580 -7760 -1200 -7720
rect -4500 -7820 1000 -7800
rect -4500 -7880 -4480 -7820
rect -4420 -7880 -4380 -7820
rect -4320 -7880 -4280 -7820
rect -4220 -7880 -4180 -7820
rect -4120 -7880 -4080 -7820
rect -4020 -7880 -3980 -7820
rect -3920 -7880 -3880 -7820
rect -3820 -7880 -3780 -7820
rect -3720 -7880 -3680 -7820
rect -3620 -7880 -3580 -7820
rect -3520 -7880 -3480 -7820
rect -3420 -7880 -3380 -7820
rect -3320 -7880 -3280 -7820
rect -3220 -7880 -3180 -7820
rect -3120 -7880 -3080 -7820
rect -3020 -7880 -2980 -7820
rect -2920 -7880 -2880 -7820
rect -2820 -7880 -2780 -7820
rect -2720 -7880 -2680 -7820
rect -2620 -7880 -2580 -7820
rect -2520 -7880 -2480 -7820
rect -2420 -7880 -2380 -7820
rect -2320 -7880 -2280 -7820
rect -2220 -7880 -2180 -7820
rect -2120 -7880 -2080 -7820
rect -2020 -7880 -1980 -7820
rect -1920 -7880 -1880 -7820
rect -1820 -7880 -1780 -7820
rect -1720 -7880 -1680 -7820
rect -1620 -7880 -1580 -7820
rect -1520 -7880 -1480 -7820
rect -1420 -7880 -1380 -7820
rect -1320 -7880 -1280 -7820
rect -1220 -7880 -1180 -7820
rect -1120 -7880 -1080 -7820
rect -1020 -7880 -980 -7820
rect -920 -7880 -880 -7820
rect -820 -7880 -780 -7820
rect -720 -7880 -680 -7820
rect -620 -7880 -580 -7820
rect -520 -7880 -480 -7820
rect -420 -7880 -380 -7820
rect -320 -7880 -280 -7820
rect -220 -7880 -180 -7820
rect -120 -7880 -80 -7820
rect -20 -7880 20 -7820
rect 80 -7880 120 -7820
rect 180 -7880 220 -7820
rect 280 -7880 320 -7820
rect 380 -7880 420 -7820
rect 480 -7880 520 -7820
rect 580 -7880 620 -7820
rect 680 -7880 720 -7820
rect 780 -7880 820 -7820
rect 880 -7880 920 -7820
rect 980 -7880 1000 -7820
rect -4500 -7920 1000 -7880
rect -4500 -7980 -4480 -7920
rect -4420 -7980 -4380 -7920
rect -4320 -7980 -4280 -7920
rect -4220 -7980 -4180 -7920
rect -4120 -7980 -4080 -7920
rect -4020 -7980 -3980 -7920
rect -3920 -7980 -3880 -7920
rect -3820 -7980 -3780 -7920
rect -3720 -7980 -3680 -7920
rect -3620 -7980 -3580 -7920
rect -3520 -7980 -3480 -7920
rect -3420 -7980 -3380 -7920
rect -3320 -7980 -3280 -7920
rect -3220 -7980 -3180 -7920
rect -3120 -7980 -3080 -7920
rect -3020 -7980 -2980 -7920
rect -2920 -7980 -2880 -7920
rect -2820 -7980 -2780 -7920
rect -2720 -7980 -2680 -7920
rect -2620 -7980 -2580 -7920
rect -2520 -7980 -2480 -7920
rect -2420 -7980 -2380 -7920
rect -2320 -7980 -2280 -7920
rect -2220 -7980 -2180 -7920
rect -2120 -7980 -2080 -7920
rect -2020 -7980 -1980 -7920
rect -1920 -7980 -1880 -7920
rect -1820 -7980 -1780 -7920
rect -1720 -7980 -1680 -7920
rect -1620 -7980 -1580 -7920
rect -1520 -7980 -1480 -7920
rect -1420 -7980 -1380 -7920
rect -1320 -7980 -1280 -7920
rect -1220 -7980 -1180 -7920
rect -1120 -7980 -1080 -7920
rect -1020 -7980 -980 -7920
rect -920 -7980 -880 -7920
rect -820 -7980 -780 -7920
rect -720 -7980 -680 -7920
rect -620 -7980 -580 -7920
rect -520 -7980 -480 -7920
rect -420 -7980 -380 -7920
rect -320 -7980 -280 -7920
rect -220 -7980 -180 -7920
rect -120 -7980 -80 -7920
rect -20 -7980 20 -7920
rect 80 -7980 120 -7920
rect 180 -7980 220 -7920
rect 280 -7980 320 -7920
rect 380 -7980 420 -7920
rect 480 -7980 520 -7920
rect 580 -7980 620 -7920
rect 680 -7980 720 -7920
rect 780 -7980 820 -7920
rect 880 -7980 920 -7920
rect 980 -7980 1000 -7920
rect -4500 -8000 1000 -7980
rect -4000 -8220 -3800 -8200
rect -4000 -8280 -3980 -8220
rect -3920 -8280 -3880 -8220
rect -3820 -8280 -3800 -8220
rect -4000 -8320 -3800 -8280
rect -4000 -8380 -3980 -8320
rect -3920 -8380 -3880 -8320
rect -3820 -8380 -3800 -8320
rect -4000 -8400 -3800 -8380
rect -2700 -8220 -2500 -8200
rect -2700 -8280 -2680 -8220
rect -2620 -8280 -2580 -8220
rect -2520 -8280 -2500 -8220
rect -2700 -8320 -2500 -8280
rect -2700 -8380 -2680 -8320
rect -2620 -8380 -2580 -8320
rect -2520 -8380 -2500 -8320
rect -2700 -8400 -2500 -8380
rect -1780 -8220 -1580 -8200
rect -1780 -8280 -1760 -8220
rect -1700 -8280 -1660 -8220
rect -1600 -8280 -1580 -8220
rect -1780 -8320 -1580 -8280
rect -1780 -8380 -1760 -8320
rect -1700 -8380 -1660 -8320
rect -1600 -8380 -1580 -8320
rect -1780 -8400 -1580 -8380
rect -1000 -8220 -800 -8200
rect -1000 -8280 -980 -8220
rect -920 -8280 -880 -8220
rect -820 -8280 -800 -8220
rect -1000 -8320 -800 -8280
rect -1000 -8380 -980 -8320
rect -920 -8380 -880 -8320
rect -820 -8380 -800 -8320
rect -1000 -8400 -800 -8380
rect 280 -8220 480 -8200
rect 280 -8280 300 -8220
rect 360 -8280 400 -8220
rect 460 -8280 480 -8220
rect 280 -8320 480 -8280
rect 280 -8380 300 -8320
rect 360 -8380 400 -8320
rect 460 -8380 480 -8320
rect 280 -8400 480 -8380
<< via1 >>
rect -4240 -4560 -4180 -4500
rect -4240 -4660 -4180 -4600
rect -4240 -4760 -4180 -4700
rect -4240 -4860 -4180 -4800
rect -4240 -4960 -4180 -4900
rect -4240 -5060 -4180 -5000
rect -4240 -5160 -4180 -5100
rect -3620 -4560 -3560 -4500
rect -3620 -4660 -3560 -4600
rect -3620 -4760 -3560 -4700
rect -3620 -4860 -3560 -4800
rect -3620 -4960 -3560 -4900
rect -3620 -5060 -3560 -5000
rect -3620 -5160 -3560 -5100
rect -3300 -4560 -3240 -4500
rect -3300 -4660 -3240 -4600
rect -3300 -4760 -3240 -4700
rect -3300 -4860 -3240 -4800
rect -3300 -4960 -3240 -4900
rect -3300 -5060 -3240 -5000
rect -3300 -5160 -3240 -5100
rect -2020 -4560 -1960 -4500
rect -2020 -4660 -1960 -4600
rect -2020 -4760 -1960 -4700
rect -2020 -4860 -1960 -4800
rect -2020 -4960 -1960 -4900
rect -2020 -5060 -1960 -5000
rect -2020 -5160 -1960 -5100
rect -1540 -4560 -1480 -4500
rect -1540 -4660 -1480 -4600
rect -1540 -4760 -1480 -4700
rect -1540 -4860 -1480 -4800
rect -1540 -4960 -1480 -4900
rect -1540 -5060 -1480 -5000
rect -1540 -5160 -1480 -5100
rect -260 -4560 -200 -4500
rect -260 -4660 -200 -4600
rect -260 -4760 -200 -4700
rect -260 -4860 -200 -4800
rect -260 -4960 -200 -4900
rect -260 -5060 -200 -5000
rect -260 -5160 -200 -5100
rect 60 -4560 120 -4500
rect 60 -4660 120 -4600
rect 60 -4760 120 -4700
rect 60 -4860 120 -4800
rect 60 -4960 120 -4900
rect 60 -5060 120 -5000
rect 60 -5160 120 -5100
rect 700 -4560 760 -4500
rect 700 -4660 760 -4600
rect 700 -4760 760 -4700
rect 700 -4860 760 -4800
rect 700 -4960 760 -4900
rect 700 -5060 760 -5000
rect 700 -5160 760 -5100
rect -2040 -5680 -1980 -5620
rect -1940 -5680 -1880 -5620
rect -1840 -5680 -1780 -5620
rect -2680 -5840 -2600 -5760
rect -2300 -5840 -2240 -5780
rect -2300 -5940 -2240 -5880
rect -2300 -6040 -2240 -5980
rect -2300 -6140 -2240 -6080
rect -2300 -6240 -2240 -6180
rect -2440 -6440 -2380 -6380
rect -2320 -6440 -2260 -6380
rect -2180 -6440 -2120 -6380
rect -1220 -5840 -1160 -5780
rect -1900 -6440 -1840 -6380
rect -1620 -6440 -1560 -6380
rect -1220 -5940 -1160 -5880
rect -1220 -6040 -1160 -5980
rect -1220 -6140 -1160 -6080
rect -1220 -6240 -1160 -6180
rect -1340 -6440 -1280 -6380
rect -1220 -6440 -1160 -6380
rect -1120 -6440 -1060 -6380
rect -3300 -6920 -3240 -6860
rect -3200 -6920 -3140 -6860
rect -3080 -6920 -3020 -6860
rect -2980 -6920 -2920 -6860
rect -3460 -7060 -3400 -7000
rect -3460 -7160 -3400 -7100
rect -3460 -7260 -3400 -7200
rect -3460 -7360 -3400 -7300
rect -3460 -7460 -3400 -7400
rect -3460 -7560 -3400 -7500
rect -2820 -7060 -2760 -7000
rect -2820 -7160 -2760 -7100
rect -2820 -7260 -2760 -7200
rect -2820 -7360 -2760 -7300
rect -2820 -7460 -2760 -7400
rect -2820 -7560 -2760 -7500
rect -2160 -7720 -2100 -7660
rect -2060 -7720 -2000 -7660
rect -1960 -7720 -1900 -7660
rect -1860 -7720 -1800 -7660
rect -500 -6920 -440 -6860
rect -400 -6920 -340 -6860
rect -260 -6920 -200 -6860
rect -160 -6920 -100 -6860
rect -660 -7060 -600 -7000
rect -660 -7160 -600 -7100
rect -660 -7260 -600 -7200
rect -660 -7360 -600 -7300
rect -660 -7460 -600 -7400
rect -660 -7560 -600 -7500
rect 0 -7060 60 -7000
rect 0 -7160 60 -7100
rect 0 -7260 60 -7200
rect 0 -7360 60 -7300
rect 0 -7460 60 -7400
rect 0 -7560 60 -7500
rect -1560 -7720 -1500 -7660
rect -1460 -7720 -1400 -7660
rect -1360 -7720 -1300 -7660
rect -1280 -7720 -1220 -7660
rect -3980 -8280 -3920 -8220
rect -3880 -8280 -3820 -8220
rect -3980 -8380 -3920 -8320
rect -3880 -8380 -3820 -8320
rect -2680 -8280 -2620 -8220
rect -2580 -8280 -2520 -8220
rect -2680 -8380 -2620 -8320
rect -2580 -8380 -2520 -8320
rect -1760 -8280 -1700 -8220
rect -1660 -8280 -1600 -8220
rect -1760 -8380 -1700 -8320
rect -1660 -8380 -1600 -8320
rect -980 -8280 -920 -8220
rect -880 -8280 -820 -8220
rect -980 -8380 -920 -8320
rect -880 -8380 -820 -8320
rect 300 -8280 360 -8220
rect 400 -8280 460 -8220
rect 300 -8380 360 -8320
rect 400 -8380 460 -8320
<< metal2 >>
rect -4260 -4500 -4140 -4420
rect -4260 -4560 -4240 -4500
rect -4180 -4560 -4140 -4500
rect -4260 -4600 -4140 -4560
rect -4260 -4660 -4240 -4600
rect -4180 -4660 -4140 -4600
rect -4260 -4700 -4140 -4660
rect -4260 -4760 -4240 -4700
rect -4180 -4760 -4140 -4700
rect -4260 -4800 -4140 -4760
rect -4260 -4860 -4240 -4800
rect -4180 -4860 -4140 -4800
rect -4260 -4900 -4140 -4860
rect -4260 -4960 -4240 -4900
rect -4180 -4960 -4140 -4900
rect -4260 -5000 -4140 -4960
rect -4260 -5060 -4240 -5000
rect -4180 -5060 -4140 -5000
rect -4260 -5100 -4140 -5060
rect -4260 -5160 -4240 -5100
rect -4180 -5160 -4140 -5100
rect -4260 -6100 -4140 -5160
rect -3660 -4500 -3540 -4420
rect -3660 -4560 -3620 -4500
rect -3560 -4560 -3540 -4500
rect -3660 -4600 -3540 -4560
rect -3660 -4660 -3620 -4600
rect -3560 -4660 -3540 -4600
rect -3660 -4700 -3540 -4660
rect -3660 -4760 -3620 -4700
rect -3560 -4760 -3540 -4700
rect -3660 -4800 -3540 -4760
rect -3660 -4860 -3620 -4800
rect -3560 -4860 -3540 -4800
rect -3660 -4900 -3540 -4860
rect -3660 -4960 -3620 -4900
rect -3560 -4960 -3540 -4900
rect -3660 -5000 -3540 -4960
rect -3660 -5060 -3620 -5000
rect -3560 -5060 -3540 -5000
rect -3660 -5100 -3540 -5060
rect -3660 -5160 -3620 -5100
rect -3560 -5160 -3540 -5100
rect -3660 -6100 -3540 -5160
rect -3320 -4500 -3200 -4420
rect -3320 -4560 -3300 -4500
rect -3240 -4560 -3200 -4500
rect -3320 -4600 -3200 -4560
rect -3320 -4660 -3300 -4600
rect -3240 -4660 -3200 -4600
rect -3320 -4700 -3200 -4660
rect -3320 -4760 -3300 -4700
rect -3240 -4760 -3200 -4700
rect -3320 -4800 -3200 -4760
rect -3320 -4860 -3300 -4800
rect -3240 -4860 -3200 -4800
rect -3320 -4900 -3200 -4860
rect -3320 -4960 -3300 -4900
rect -3240 -4960 -3200 -4900
rect -3320 -5000 -3200 -4960
rect -3320 -5060 -3300 -5000
rect -3240 -5060 -3200 -5000
rect -3320 -5100 -3200 -5060
rect -3320 -5160 -3300 -5100
rect -3240 -5160 -3200 -5100
rect -3320 -5440 -3200 -5160
rect -3320 -5520 -3300 -5440
rect -3220 -5520 -3200 -5440
rect -3320 -5540 -3200 -5520
rect -2060 -4500 -1940 -4420
rect -2060 -4560 -2020 -4500
rect -1960 -4560 -1940 -4500
rect -2060 -4600 -1940 -4560
rect -2060 -4660 -2020 -4600
rect -1960 -4660 -1940 -4600
rect -2060 -4700 -1940 -4660
rect -2060 -4760 -2020 -4700
rect -1960 -4760 -1940 -4700
rect -2060 -4800 -1940 -4760
rect -2060 -4860 -2020 -4800
rect -1960 -4860 -1940 -4800
rect -2060 -4900 -1940 -4860
rect -2060 -4960 -2020 -4900
rect -1960 -4960 -1940 -4900
rect -2060 -5000 -1940 -4960
rect -2060 -5060 -2020 -5000
rect -1960 -5060 -1940 -5000
rect -2060 -5100 -1940 -5060
rect -2060 -5160 -2020 -5100
rect -1960 -5160 -1940 -5100
rect -2060 -5440 -1940 -5160
rect -2060 -5520 -2040 -5440
rect -1960 -5520 -1940 -5440
rect -2060 -5540 -1940 -5520
rect -1560 -4500 -1440 -4420
rect -1560 -4560 -1540 -4500
rect -1480 -4560 -1440 -4500
rect -1560 -4600 -1440 -4560
rect -1560 -4660 -1540 -4600
rect -1480 -4660 -1440 -4600
rect -1560 -4700 -1440 -4660
rect -1560 -4760 -1540 -4700
rect -1480 -4760 -1440 -4700
rect -1560 -4800 -1440 -4760
rect -1560 -4860 -1540 -4800
rect -1480 -4860 -1440 -4800
rect -1560 -4900 -1440 -4860
rect -1560 -4960 -1540 -4900
rect -1480 -4960 -1440 -4900
rect -1560 -5000 -1440 -4960
rect -1560 -5060 -1540 -5000
rect -1480 -5060 -1440 -5000
rect -1560 -5100 -1440 -5060
rect -1560 -5160 -1540 -5100
rect -1480 -5160 -1440 -5100
rect -1560 -5440 -1440 -5160
rect -1560 -5520 -1540 -5440
rect -1460 -5520 -1440 -5440
rect -1560 -5540 -1440 -5520
rect -300 -4500 -180 -4400
rect -300 -4560 -260 -4500
rect -200 -4560 -180 -4500
rect -300 -4600 -180 -4560
rect -300 -4660 -260 -4600
rect -200 -4660 -180 -4600
rect -300 -4700 -180 -4660
rect -300 -4760 -260 -4700
rect -200 -4760 -180 -4700
rect -300 -4800 -180 -4760
rect -300 -4860 -260 -4800
rect -200 -4860 -180 -4800
rect -300 -4900 -180 -4860
rect -300 -4960 -260 -4900
rect -200 -4960 -180 -4900
rect -300 -5000 -180 -4960
rect -300 -5060 -260 -5000
rect -200 -5060 -180 -5000
rect -300 -5100 -180 -5060
rect -300 -5160 -260 -5100
rect -200 -5160 -180 -5100
rect -300 -5440 -180 -5160
rect -300 -5520 -280 -5440
rect -200 -5520 -180 -5440
rect -300 -5540 -180 -5520
rect 40 -4500 160 -4420
rect 40 -4560 60 -4500
rect 120 -4560 160 -4500
rect 40 -4600 160 -4560
rect 40 -4660 60 -4600
rect 120 -4660 160 -4600
rect 40 -4700 160 -4660
rect 40 -4760 60 -4700
rect 120 -4760 160 -4700
rect 40 -4800 160 -4760
rect 40 -4860 60 -4800
rect 120 -4860 160 -4800
rect 40 -4900 160 -4860
rect 40 -4960 60 -4900
rect 120 -4960 160 -4900
rect 40 -5000 160 -4960
rect 40 -5060 60 -5000
rect 120 -5060 160 -5000
rect 40 -5100 160 -5060
rect 40 -5160 60 -5100
rect 120 -5160 160 -5100
rect -2060 -5620 -1680 -5600
rect -2060 -5680 -2040 -5620
rect -1980 -5680 -1940 -5620
rect -1880 -5680 -1840 -5620
rect -1780 -5680 -1680 -5620
rect -2060 -5700 -1680 -5680
rect -2700 -5760 -580 -5740
rect -2700 -5840 -2680 -5760
rect -2600 -5780 -1080 -5760
rect -2600 -5840 -2300 -5780
rect -2240 -5840 -1220 -5780
rect -1160 -5840 -1080 -5780
rect -1000 -5840 -960 -5760
rect -880 -5840 -840 -5760
rect -760 -5840 -720 -5760
rect -640 -5840 -580 -5760
rect -2700 -5860 -580 -5840
rect -2320 -5880 -2220 -5860
rect -2320 -5940 -2300 -5880
rect -2240 -5940 -2220 -5880
rect -2320 -5980 -2220 -5940
rect -2320 -6040 -2300 -5980
rect -2240 -6040 -2220 -5980
rect -2320 -6080 -2220 -6040
rect -4460 -6220 -2740 -6100
rect -2320 -6140 -2300 -6080
rect -2240 -6140 -2220 -6080
rect -2320 -6180 -2220 -6140
rect -4000 -6860 -3800 -6840
rect -4000 -6920 -3980 -6860
rect -3920 -6920 -3880 -6860
rect -3820 -6920 -3800 -6860
rect -4000 -6960 -3800 -6920
rect -4000 -7020 -3980 -6960
rect -3920 -7020 -3880 -6960
rect -3820 -7020 -3800 -6960
rect -4000 -8220 -3800 -7020
rect -3480 -7000 -3360 -6220
rect -3320 -6860 -2900 -6840
rect -3320 -6920 -3300 -6860
rect -3240 -6920 -3200 -6860
rect -3140 -6920 -3080 -6860
rect -3020 -6920 -2980 -6860
rect -2920 -6920 -2900 -6860
rect -3320 -6940 -2900 -6920
rect -3480 -7060 -3460 -7000
rect -3400 -7060 -3360 -7000
rect -3480 -7100 -3360 -7060
rect -3480 -7160 -3460 -7100
rect -3400 -7160 -3360 -7100
rect -3480 -7200 -3360 -7160
rect -3480 -7260 -3460 -7200
rect -3400 -7260 -3360 -7200
rect -3480 -7300 -3360 -7260
rect -3480 -7360 -3460 -7300
rect -3400 -7360 -3360 -7300
rect -3480 -7400 -3360 -7360
rect -3480 -7460 -3460 -7400
rect -3400 -7460 -3360 -7400
rect -3480 -7500 -3360 -7460
rect -3480 -7560 -3460 -7500
rect -3400 -7560 -3360 -7500
rect -3480 -7580 -3360 -7560
rect -2860 -7000 -2740 -6220
rect -2860 -7060 -2820 -7000
rect -2760 -7060 -2740 -7000
rect -2860 -7100 -2740 -7060
rect -2860 -7160 -2820 -7100
rect -2760 -7160 -2740 -7100
rect -2860 -7200 -2740 -7160
rect -2860 -7260 -2820 -7200
rect -2760 -7260 -2740 -7200
rect -2860 -7300 -2740 -7260
rect -2860 -7360 -2820 -7300
rect -2760 -7360 -2740 -7300
rect -2860 -7400 -2740 -7360
rect -2860 -7460 -2820 -7400
rect -2760 -7460 -2740 -7400
rect -2860 -7500 -2740 -7460
rect -2860 -7560 -2820 -7500
rect -2760 -7560 -2740 -7500
rect -2860 -7580 -2740 -7560
rect -2700 -6500 -2500 -6200
rect -2320 -6240 -2300 -6180
rect -2240 -6240 -2220 -6180
rect -2320 -6320 -2220 -6240
rect -1240 -5880 -1140 -5860
rect -1240 -5940 -1220 -5880
rect -1160 -5940 -1140 -5880
rect -1240 -5980 -1140 -5940
rect -1240 -6040 -1220 -5980
rect -1160 -6040 -1140 -5980
rect -1240 -6080 -1140 -6040
rect -1240 -6140 -1220 -6080
rect -1160 -6140 -1140 -6080
rect 40 -6100 160 -5160
rect 660 -4500 780 -4420
rect 660 -4560 700 -4500
rect 760 -4560 780 -4500
rect 660 -4600 780 -4560
rect 660 -4660 700 -4600
rect 760 -4660 780 -4600
rect 660 -4700 780 -4660
rect 660 -4760 700 -4700
rect 760 -4760 780 -4700
rect 660 -4800 780 -4760
rect 660 -4860 700 -4800
rect 760 -4860 780 -4800
rect 660 -4900 780 -4860
rect 660 -4960 700 -4900
rect 760 -4960 780 -4900
rect 660 -5000 780 -4960
rect 660 -5060 700 -5000
rect 760 -5060 780 -5000
rect 660 -5100 780 -5060
rect 660 -5160 700 -5100
rect 760 -5160 780 -5100
rect 280 -6100 483 -6097
rect 660 -6100 780 -5160
rect -1240 -6180 -1140 -6140
rect -1240 -6240 -1220 -6180
rect -1160 -6240 -1140 -6180
rect -1240 -6320 -1140 -6240
rect -2460 -6380 -2100 -6360
rect -2460 -6440 -2440 -6380
rect -2380 -6440 -2320 -6380
rect -2260 -6440 -2180 -6380
rect -2120 -6440 -2100 -6380
rect -2460 -6460 -2100 -6440
rect -1920 -6380 -1820 -6360
rect -1920 -6440 -1900 -6380
rect -1840 -6440 -1820 -6380
rect -1920 -6500 -1820 -6440
rect -1640 -6380 -1540 -6360
rect -1640 -6440 -1620 -6380
rect -1560 -6440 -1540 -6380
rect -1640 -6500 -1540 -6440
rect -1360 -6380 -1040 -6360
rect -1360 -6440 -1340 -6380
rect -1280 -6440 -1220 -6380
rect -1160 -6440 -1120 -6380
rect -1060 -6440 -1040 -6380
rect -1360 -6460 -1040 -6440
rect -2700 -6600 -1140 -6500
rect -4000 -8280 -3980 -8220
rect -3920 -8280 -3880 -8220
rect -3820 -8280 -3800 -8220
rect -4000 -8320 -3800 -8280
rect -4000 -8380 -3980 -8320
rect -3920 -8380 -3880 -8320
rect -3820 -8380 -3800 -8320
rect -4000 -8400 -3800 -8380
rect -2700 -8220 -2500 -6600
rect -1000 -6660 -800 -6200
rect -2320 -6680 -800 -6660
rect -2320 -6740 -2300 -6680
rect -2240 -6740 -2180 -6680
rect -2120 -6740 -2040 -6680
rect -1980 -6740 -1480 -6680
rect -1420 -6740 -1340 -6680
rect -1280 -6740 -1220 -6680
rect -1160 -6740 -800 -6680
rect -2320 -6760 -800 -6740
rect -2180 -7660 -1200 -7600
rect -2180 -7720 -2160 -7660
rect -2100 -7720 -2060 -7660
rect -2000 -7720 -1960 -7660
rect -1900 -7720 -1860 -7660
rect -1800 -7720 -1560 -7660
rect -1500 -7720 -1460 -7660
rect -1400 -7720 -1360 -7660
rect -1300 -7720 -1280 -7660
rect -1220 -7720 -1200 -7660
rect -2180 -7760 -1200 -7720
rect -2700 -8280 -2680 -8220
rect -2620 -8280 -2580 -8220
rect -2520 -8280 -2500 -8220
rect -2700 -8320 -2500 -8280
rect -2700 -8380 -2680 -8320
rect -2620 -8380 -2580 -8320
rect -2520 -8380 -2500 -8320
rect -2700 -8400 -2500 -8380
rect -1780 -8220 -1580 -7760
rect -1780 -8280 -1760 -8220
rect -1700 -8280 -1660 -8220
rect -1600 -8280 -1580 -8220
rect -1780 -8320 -1580 -8280
rect -1780 -8380 -1760 -8320
rect -1700 -8380 -1660 -8320
rect -1600 -8380 -1580 -8320
rect -1780 -8400 -1580 -8380
rect -1000 -8220 -800 -6760
rect -700 -6220 940 -6100
rect -700 -6980 -580 -6220
rect -520 -6860 -80 -6840
rect -520 -6920 -500 -6860
rect -440 -6920 -400 -6860
rect -340 -6920 -260 -6860
rect -200 -6920 -160 -6860
rect -100 -6920 -80 -6860
rect -520 -6940 -80 -6920
rect -20 -6980 100 -6220
rect -700 -7000 -540 -6980
rect -700 -7060 -660 -7000
rect -600 -7060 -540 -7000
rect -700 -7100 -540 -7060
rect -700 -7160 -660 -7100
rect -600 -7160 -540 -7100
rect -700 -7200 -540 -7160
rect -700 -7260 -660 -7200
rect -600 -7260 -540 -7200
rect -700 -7300 -540 -7260
rect -700 -7360 -660 -7300
rect -600 -7360 -540 -7300
rect -700 -7400 -540 -7360
rect -700 -7460 -660 -7400
rect -600 -7460 -540 -7400
rect -700 -7500 -540 -7460
rect -700 -7560 -660 -7500
rect -600 -7560 -540 -7500
rect -700 -7580 -540 -7560
rect -60 -7000 100 -6980
rect -60 -7060 0 -7000
rect 60 -7060 100 -7000
rect -60 -7100 100 -7060
rect -60 -7160 0 -7100
rect 60 -7160 100 -7100
rect -60 -7200 100 -7160
rect -60 -7260 0 -7200
rect 60 -7260 100 -7200
rect -60 -7300 100 -7260
rect -60 -7360 0 -7300
rect 60 -7360 100 -7300
rect -60 -7400 100 -7360
rect -60 -7460 0 -7400
rect 60 -7460 100 -7400
rect -60 -7500 100 -7460
rect -60 -7560 0 -7500
rect 60 -7560 100 -7500
rect -60 -7580 100 -7560
rect -1000 -8280 -980 -8220
rect -920 -8280 -880 -8220
rect -820 -8280 -800 -8220
rect -1000 -8320 -800 -8280
rect -1000 -8380 -980 -8320
rect -920 -8380 -880 -8320
rect -820 -8380 -800 -8320
rect -1000 -8400 -800 -8380
rect 280 -8220 483 -6220
rect 280 -8280 300 -8220
rect 360 -8280 400 -8220
rect 460 -8280 483 -8220
rect 280 -8320 483 -8280
rect 280 -8380 300 -8320
rect 360 -8380 400 -8320
rect 460 -8380 483 -8320
rect 280 -8399 483 -8380
rect 280 -8400 480 -8399
<< via2 >>
rect -3300 -5520 -3220 -5440
rect -2040 -5520 -1960 -5440
rect -1540 -5520 -1460 -5440
rect -280 -5520 -200 -5440
rect -2040 -5680 -1980 -5620
rect -1940 -5680 -1880 -5620
rect -1840 -5680 -1780 -5620
rect -1080 -5840 -1000 -5760
rect -960 -5840 -880 -5760
rect -840 -5840 -760 -5760
rect -720 -5840 -640 -5760
rect -3980 -6920 -3920 -6860
rect -3880 -6920 -3820 -6860
rect -3980 -7020 -3920 -6960
rect -3880 -7020 -3820 -6960
rect -3300 -6920 -3240 -6860
rect -3200 -6920 -3140 -6860
rect -3080 -6920 -3020 -6860
rect -2980 -6920 -2920 -6860
rect -2440 -6440 -2380 -6380
rect -2320 -6440 -2260 -6380
rect -2180 -6440 -2120 -6380
rect -1340 -6440 -1280 -6380
rect -1220 -6440 -1160 -6380
rect -1120 -6440 -1060 -6380
rect -2300 -6740 -2240 -6680
rect -2180 -6740 -2120 -6680
rect -2040 -6740 -1980 -6680
rect -1480 -6740 -1420 -6680
rect -1340 -6740 -1280 -6680
rect -1220 -6740 -1160 -6680
rect -500 -6920 -440 -6860
rect -400 -6920 -340 -6860
rect -260 -6920 -200 -6860
rect -160 -6920 -100 -6860
<< metal3 >>
rect -3320 -5440 -1940 -5420
rect -3320 -5520 -3300 -5440
rect -3220 -5520 -2040 -5440
rect -1960 -5520 -1940 -5440
rect -3320 -5540 -1940 -5520
rect -1560 -5440 -180 -5420
rect -1560 -5520 -1540 -5440
rect -1460 -5520 -280 -5440
rect -200 -5520 -180 -5440
rect -1560 -5540 -180 -5520
rect -2860 -5600 -2740 -5540
rect -2860 -5620 -1680 -5600
rect -2860 -5680 -2040 -5620
rect -1980 -5680 -1940 -5620
rect -1880 -5680 -1840 -5620
rect -1780 -5680 -1680 -5620
rect -2860 -5700 -1680 -5680
rect -760 -5740 -640 -5540
rect -1100 -5760 -580 -5740
rect -1100 -5840 -1080 -5760
rect -1000 -5840 -960 -5760
rect -880 -5840 -840 -5760
rect -760 -5840 -720 -5760
rect -640 -5840 -580 -5760
rect -1100 -5860 -580 -5840
rect -2460 -6380 -2100 -6360
rect -2460 -6440 -2440 -6380
rect -2380 -6440 -2320 -6380
rect -2260 -6440 -2180 -6380
rect -2120 -6440 -2100 -6380
rect -2460 -6460 -2100 -6440
rect -2200 -6660 -2100 -6460
rect -1360 -6380 -1040 -6360
rect -1360 -6440 -1340 -6380
rect -1280 -6440 -1220 -6380
rect -1160 -6440 -1120 -6380
rect -1060 -6440 -1040 -6380
rect -1360 -6460 -1040 -6440
rect -1360 -6660 -1260 -6460
rect -2320 -6680 -1960 -6660
rect -2320 -6740 -2300 -6680
rect -2240 -6740 -2180 -6680
rect -2120 -6740 -2040 -6680
rect -1980 -6740 -1960 -6680
rect -2320 -6760 -1960 -6740
rect -1500 -6680 -1140 -6660
rect -1500 -6740 -1480 -6680
rect -1420 -6740 -1340 -6680
rect -1280 -6740 -1220 -6680
rect -1160 -6740 -1140 -6680
rect -1500 -6760 -1140 -6740
rect -4000 -6860 -40 -6840
rect -4000 -6920 -3980 -6860
rect -3920 -6920 -3880 -6860
rect -3820 -6920 -3300 -6860
rect -3240 -6920 -3200 -6860
rect -3140 -6920 -3080 -6860
rect -3020 -6920 -2980 -6860
rect -2920 -6920 -500 -6860
rect -440 -6920 -400 -6860
rect -340 -6920 -260 -6860
rect -200 -6920 -160 -6860
rect -100 -6920 -40 -6860
rect -4000 -6940 -40 -6920
rect -4000 -6960 -3800 -6940
rect -4000 -7020 -3980 -6960
rect -3920 -7020 -3880 -6960
rect -3820 -7020 -3800 -6960
rect -4000 -7040 -3800 -7020
use sky130_fd_pr__nfet_g5v0d10v5_KHGXMS  sky130_fd_pr__nfet_g5v0d10v5_KHGXMS_0
timestamp 1769077132
transform 1 0 -3103 0 1 -7243
box -297 -357 297 357
use sky130_fd_pr__nfet_g5v0d10v5_KHGXMS  sky130_fd_pr__nfet_g5v0d10v5_KHGXMS_1
timestamp 1769077132
transform 1 0 -303 0 1 -7243
box -297 -357 297 357
use sky130_fd_pr__pfet_g5v0d10v5_S3L597  sky130_fd_pr__pfet_g5v0d10v5_S3L597_0
timestamp 1769076474
transform 1 0 -861 0 1 -4847
box -691 -439 691 477
use sky130_fd_pr__pfet_g5v0d10v5_S3L597  sky130_fd_pr__pfet_g5v0d10v5_S3L597_1
timestamp 1769076474
transform 1 0 -2621 0 1 -4847
box -691 -439 691 477
use sky130_fd_pr__pfet_g5v0d10v5_SXU6V5  sky130_fd_pr__pfet_g5v0d10v5_SXU6V5_0
timestamp 1769076474
transform 1 0 411 0 1 -4847
box -363 -439 363 477
use sky130_fd_pr__pfet_g5v0d10v5_SXU6V5  sky130_fd_pr__pfet_g5v0d10v5_SXU6V5_1
timestamp 1769076474
transform 1 0 -3889 0 1 -4847
box -363 -439 363 477
use sky130_fd_pr__nfet_g5v0d10v5_P5847U  XM2
timestamp 1769077132
transform 1 0 -1735 0 1 -6155
box -525 -265 525 265
use sky130_fd_pr__nfet_g5v0d10v5_3ZGXMS  XM8
timestamp 1769084796
transform 1 0 -1683 0 1 -7223
box -297 -357 297 357
<< labels >>
flabel metal1 -1900 -8000 -1700 -7800 0 FreeSans 256 0 0 0 VSS
port 6 nsew
flabel metal1 -4000 -8400 -3800 -8200 0 FreeSans 256 0 0 0 B2
port 5 nsew
flabel metal1 -1892 -4306 -1692 -4106 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -1000 -8400 -800 -8200 0 FreeSans 256 0 0 0 REF
port 1 nsew
flabel metal1 -2700 -8400 -2500 -8200 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal1 -1780 -8400 -1580 -8200 0 FreeSans 256 0 0 0 B1
port 4 nsew
flabel metal1 280 -8400 480 -8200 0 FreeSans 256 0 0 0 OUT
port 3 nsew
<< end >>
