magic
tech sky130A
magscale 1 2
timestamp 1770083657
<< pwell >>
rect 1274 3474 6926 3626
rect 1274 3274 3926 3474
rect 1274 2026 1726 3274
rect 2574 2026 2926 3274
rect 3774 2026 3926 3274
rect 1274 1874 3926 2026
rect 4274 3274 6926 3474
rect 4274 2026 4426 3274
rect 5274 2026 5626 3274
rect 6474 2026 6926 3274
rect 4274 1874 6926 2026
rect 1274 1426 1426 1874
rect 6774 1426 6926 1874
rect 1274 1274 3926 1426
rect 1274 26 1726 1274
rect 2574 26 2926 1274
rect 3774 26 3926 1274
rect 1274 -174 3926 26
rect 4274 1274 6926 1426
rect 4274 26 4426 1274
rect 5274 26 5626 1274
rect 6474 26 6926 1274
rect 4274 -174 6926 26
rect 1274 -326 6926 -174
<< psubdiff >>
rect 1300 3567 6900 3600
rect 1300 3533 1441 3567
rect 1475 3533 1509 3567
rect 1543 3533 1577 3567
rect 1611 3533 1645 3567
rect 1679 3533 1713 3567
rect 1747 3533 1781 3567
rect 1815 3533 1849 3567
rect 1883 3533 1917 3567
rect 1951 3533 1985 3567
rect 2019 3533 2053 3567
rect 2087 3533 2121 3567
rect 2155 3533 2189 3567
rect 2223 3533 2257 3567
rect 2291 3533 2325 3567
rect 2359 3533 2393 3567
rect 2427 3533 2461 3567
rect 2495 3533 2529 3567
rect 2563 3533 2597 3567
rect 2631 3533 2665 3567
rect 2699 3533 2733 3567
rect 2767 3533 2801 3567
rect 2835 3533 2869 3567
rect 2903 3533 2937 3567
rect 2971 3533 3005 3567
rect 3039 3533 3073 3567
rect 3107 3533 3141 3567
rect 3175 3533 3209 3567
rect 3243 3533 3277 3567
rect 3311 3533 3345 3567
rect 3379 3533 3413 3567
rect 3447 3533 3481 3567
rect 3515 3533 3549 3567
rect 3583 3533 3617 3567
rect 3651 3533 3685 3567
rect 3719 3533 3753 3567
rect 3787 3533 3821 3567
rect 3855 3533 3889 3567
rect 3923 3533 3957 3567
rect 3991 3533 4025 3567
rect 4059 3533 4093 3567
rect 4127 3533 4161 3567
rect 4195 3533 4229 3567
rect 4263 3533 4297 3567
rect 4331 3533 4365 3567
rect 4399 3533 4433 3567
rect 4467 3533 4501 3567
rect 4535 3533 4569 3567
rect 4603 3533 4637 3567
rect 4671 3533 4705 3567
rect 4739 3533 4773 3567
rect 4807 3533 4841 3567
rect 4875 3533 4909 3567
rect 4943 3533 4977 3567
rect 5011 3533 5045 3567
rect 5079 3533 5113 3567
rect 5147 3533 5181 3567
rect 5215 3533 5249 3567
rect 5283 3533 5317 3567
rect 5351 3533 5385 3567
rect 5419 3533 5453 3567
rect 5487 3533 5521 3567
rect 5555 3533 5589 3567
rect 5623 3533 5657 3567
rect 5691 3533 5725 3567
rect 5759 3533 5793 3567
rect 5827 3533 5861 3567
rect 5895 3533 5929 3567
rect 5963 3533 5997 3567
rect 6031 3533 6065 3567
rect 6099 3533 6133 3567
rect 6167 3533 6201 3567
rect 6235 3533 6269 3567
rect 6303 3533 6337 3567
rect 6371 3533 6405 3567
rect 6439 3533 6473 3567
rect 6507 3533 6541 3567
rect 6575 3533 6609 3567
rect 6643 3533 6677 3567
rect 6711 3533 6745 3567
rect 6779 3533 6900 3567
rect 1300 3500 6900 3533
rect 1300 3469 1400 3500
rect 1300 3435 1333 3469
rect 1367 3435 1400 3469
rect 1300 3401 1400 3435
rect 1300 3367 1333 3401
rect 1367 3367 1400 3401
rect 6800 3464 6900 3500
rect 6800 3430 6833 3464
rect 6867 3430 6900 3464
rect 1300 3333 1400 3367
rect 1300 3299 1333 3333
rect 1367 3299 1400 3333
rect 1300 3265 1400 3299
rect 1300 3231 1333 3265
rect 1367 3231 1400 3265
rect 1300 3197 1400 3231
rect 1300 3163 1333 3197
rect 1367 3163 1400 3197
rect 1300 3129 1400 3163
rect 1300 3095 1333 3129
rect 1367 3095 1400 3129
rect 1300 3061 1400 3095
rect 1300 3027 1333 3061
rect 1367 3027 1400 3061
rect 1300 2993 1400 3027
rect 1300 2959 1333 2993
rect 1367 2959 1400 2993
rect 1300 2925 1400 2959
rect 1300 2891 1333 2925
rect 1367 2891 1400 2925
rect 1300 2857 1400 2891
rect 1300 2823 1333 2857
rect 1367 2823 1400 2857
rect 1300 2789 1400 2823
rect 1300 2755 1333 2789
rect 1367 2755 1400 2789
rect 1300 2721 1400 2755
rect 1300 2687 1333 2721
rect 1367 2687 1400 2721
rect 1300 2653 1400 2687
rect 1300 2619 1333 2653
rect 1367 2619 1400 2653
rect 1300 2585 1400 2619
rect 1300 2551 1333 2585
rect 1367 2551 1400 2585
rect 1300 2517 1400 2551
rect 1300 2483 1333 2517
rect 1367 2483 1400 2517
rect 1300 2449 1400 2483
rect 1300 2415 1333 2449
rect 1367 2415 1400 2449
rect 1300 2381 1400 2415
rect 1300 2347 1333 2381
rect 1367 2347 1400 2381
rect 1300 2313 1400 2347
rect 1300 2279 1333 2313
rect 1367 2279 1400 2313
rect 1300 2245 1400 2279
rect 1300 2211 1333 2245
rect 1367 2211 1400 2245
rect 1300 2177 1400 2211
rect 1300 2143 1333 2177
rect 1367 2143 1400 2177
rect 1300 2109 1400 2143
rect 1300 2075 1333 2109
rect 1367 2075 1400 2109
rect 1300 2041 1400 2075
rect 1300 2007 1333 2041
rect 1367 2007 1400 2041
rect 1300 1973 1400 2007
rect 1300 1939 1333 1973
rect 1367 1939 1400 1973
rect 1300 1905 1400 1939
rect 1300 1871 1333 1905
rect 1367 1871 1400 1905
rect 1600 3367 2700 3400
rect 1600 3333 1623 3367
rect 1657 3333 1691 3367
rect 1725 3333 1759 3367
rect 1793 3333 1827 3367
rect 1861 3333 1895 3367
rect 1929 3333 1963 3367
rect 1997 3333 2031 3367
rect 2065 3333 2099 3367
rect 2133 3333 2167 3367
rect 2201 3333 2235 3367
rect 2269 3333 2303 3367
rect 2337 3333 2371 3367
rect 2405 3333 2439 3367
rect 2473 3333 2507 3367
rect 2541 3333 2575 3367
rect 2609 3333 2643 3367
rect 2677 3333 2700 3367
rect 1600 3300 2700 3333
rect 1600 2000 1700 3300
rect 2600 2000 2700 3300
rect 1600 1900 2700 2000
rect 2800 3367 3900 3400
rect 2800 3333 2823 3367
rect 2857 3333 2891 3367
rect 2925 3333 2959 3367
rect 2993 3333 3027 3367
rect 3061 3333 3095 3367
rect 3129 3333 3163 3367
rect 3197 3333 3231 3367
rect 3265 3333 3299 3367
rect 3333 3333 3367 3367
rect 3401 3333 3435 3367
rect 3469 3333 3503 3367
rect 3537 3333 3571 3367
rect 3605 3333 3639 3367
rect 3673 3333 3707 3367
rect 3741 3333 3775 3367
rect 3809 3333 3843 3367
rect 3877 3333 3900 3367
rect 2800 3300 3900 3333
rect 2800 2000 2900 3300
rect 3800 2000 3900 3300
rect 2800 1900 3900 2000
rect 4300 3367 5400 3400
rect 4300 3333 4323 3367
rect 4357 3333 4391 3367
rect 4425 3333 4459 3367
rect 4493 3333 4527 3367
rect 4561 3333 4595 3367
rect 4629 3333 4663 3367
rect 4697 3333 4731 3367
rect 4765 3333 4799 3367
rect 4833 3333 4867 3367
rect 4901 3333 4935 3367
rect 4969 3333 5003 3367
rect 5037 3333 5071 3367
rect 5105 3333 5139 3367
rect 5173 3333 5207 3367
rect 5241 3333 5275 3367
rect 5309 3333 5343 3367
rect 5377 3333 5400 3367
rect 4300 3300 5400 3333
rect 4300 2000 4400 3300
rect 5300 2000 5400 3300
rect 4300 1900 5400 2000
rect 5500 3367 6600 3400
rect 5500 3333 5523 3367
rect 5557 3333 5591 3367
rect 5625 3333 5659 3367
rect 5693 3333 5727 3367
rect 5761 3333 5795 3367
rect 5829 3333 5863 3367
rect 5897 3333 5931 3367
rect 5965 3333 5999 3367
rect 6033 3333 6067 3367
rect 6101 3333 6135 3367
rect 6169 3333 6203 3367
rect 6237 3333 6271 3367
rect 6305 3333 6339 3367
rect 6373 3333 6407 3367
rect 6441 3333 6475 3367
rect 6509 3333 6543 3367
rect 6577 3333 6600 3367
rect 5500 3300 6600 3333
rect 5500 2000 5600 3300
rect 6500 2000 6600 3300
rect 5500 1900 6600 2000
rect 6800 3396 6900 3430
rect 6800 3362 6833 3396
rect 6867 3362 6900 3396
rect 6800 3328 6900 3362
rect 6800 3294 6833 3328
rect 6867 3294 6900 3328
rect 6800 3260 6900 3294
rect 6800 3226 6833 3260
rect 6867 3226 6900 3260
rect 6800 3192 6900 3226
rect 6800 3158 6833 3192
rect 6867 3158 6900 3192
rect 6800 3124 6900 3158
rect 6800 3090 6833 3124
rect 6867 3090 6900 3124
rect 6800 3056 6900 3090
rect 6800 3022 6833 3056
rect 6867 3022 6900 3056
rect 6800 2988 6900 3022
rect 6800 2954 6833 2988
rect 6867 2954 6900 2988
rect 6800 2920 6900 2954
rect 6800 2886 6833 2920
rect 6867 2886 6900 2920
rect 6800 2852 6900 2886
rect 6800 2818 6833 2852
rect 6867 2818 6900 2852
rect 6800 2784 6900 2818
rect 6800 2750 6833 2784
rect 6867 2750 6900 2784
rect 6800 2716 6900 2750
rect 6800 2682 6833 2716
rect 6867 2682 6900 2716
rect 6800 2648 6900 2682
rect 6800 2614 6833 2648
rect 6867 2614 6900 2648
rect 6800 2580 6900 2614
rect 6800 2546 6833 2580
rect 6867 2546 6900 2580
rect 6800 2512 6900 2546
rect 6800 2478 6833 2512
rect 6867 2478 6900 2512
rect 6800 2444 6900 2478
rect 6800 2410 6833 2444
rect 6867 2410 6900 2444
rect 6800 2376 6900 2410
rect 6800 2342 6833 2376
rect 6867 2342 6900 2376
rect 6800 2308 6900 2342
rect 6800 2274 6833 2308
rect 6867 2274 6900 2308
rect 6800 2240 6900 2274
rect 6800 2206 6833 2240
rect 6867 2206 6900 2240
rect 6800 2172 6900 2206
rect 6800 2138 6833 2172
rect 6867 2138 6900 2172
rect 6800 2104 6900 2138
rect 6800 2070 6833 2104
rect 6867 2070 6900 2104
rect 6800 2036 6900 2070
rect 6800 2002 6833 2036
rect 6867 2002 6900 2036
rect 6800 1968 6900 2002
rect 6800 1934 6833 1968
rect 6867 1934 6900 1968
rect 6800 1900 6900 1934
rect 1300 1837 1400 1871
rect 1300 1803 1333 1837
rect 1367 1803 1400 1837
rect 1300 1769 1400 1803
rect 1300 1735 1333 1769
rect 1367 1735 1400 1769
rect 1300 1701 1400 1735
rect 1300 1667 1333 1701
rect 1367 1667 1400 1701
rect 1300 1633 1400 1667
rect 1300 1599 1333 1633
rect 1367 1599 1400 1633
rect 1300 1565 1400 1599
rect 1300 1531 1333 1565
rect 1367 1531 1400 1565
rect 1300 1497 1400 1531
rect 1300 1463 1333 1497
rect 1367 1463 1400 1497
rect 1300 1429 1400 1463
rect 1300 1395 1333 1429
rect 1367 1395 1400 1429
rect 6800 1866 6833 1900
rect 6867 1866 6900 1900
rect 6800 1832 6900 1866
rect 6800 1798 6833 1832
rect 6867 1798 6900 1832
rect 6800 1764 6900 1798
rect 6800 1730 6833 1764
rect 6867 1730 6900 1764
rect 6800 1696 6900 1730
rect 6800 1662 6833 1696
rect 6867 1662 6900 1696
rect 6800 1628 6900 1662
rect 6800 1594 6833 1628
rect 6867 1594 6900 1628
rect 6800 1560 6900 1594
rect 6800 1526 6833 1560
rect 6867 1526 6900 1560
rect 6800 1492 6900 1526
rect 6800 1458 6833 1492
rect 6867 1458 6900 1492
rect 6800 1424 6900 1458
rect 1300 1361 1400 1395
rect 1300 1327 1333 1361
rect 1367 1327 1400 1361
rect 1300 1293 1400 1327
rect 1300 1259 1333 1293
rect 1367 1259 1400 1293
rect 1300 1225 1400 1259
rect 1300 1191 1333 1225
rect 1367 1191 1400 1225
rect 1300 1157 1400 1191
rect 1300 1123 1333 1157
rect 1367 1123 1400 1157
rect 1300 1089 1400 1123
rect 1300 1055 1333 1089
rect 1367 1055 1400 1089
rect 1300 1021 1400 1055
rect 1300 987 1333 1021
rect 1367 987 1400 1021
rect 1300 953 1400 987
rect 1300 919 1333 953
rect 1367 919 1400 953
rect 1300 885 1400 919
rect 1300 851 1333 885
rect 1367 851 1400 885
rect 1300 817 1400 851
rect 1300 783 1333 817
rect 1367 783 1400 817
rect 1300 749 1400 783
rect 1300 715 1333 749
rect 1367 715 1400 749
rect 1300 681 1400 715
rect 1300 647 1333 681
rect 1367 647 1400 681
rect 1300 613 1400 647
rect 1300 579 1333 613
rect 1367 579 1400 613
rect 1300 545 1400 579
rect 1300 511 1333 545
rect 1367 511 1400 545
rect 1300 477 1400 511
rect 1300 443 1333 477
rect 1367 443 1400 477
rect 1300 409 1400 443
rect 1300 375 1333 409
rect 1367 375 1400 409
rect 1300 341 1400 375
rect 1300 307 1333 341
rect 1367 307 1400 341
rect 1300 273 1400 307
rect 1300 239 1333 273
rect 1367 239 1400 273
rect 1300 205 1400 239
rect 1300 171 1333 205
rect 1367 171 1400 205
rect 1300 137 1400 171
rect 1300 103 1333 137
rect 1367 103 1400 137
rect 1300 69 1400 103
rect 1300 35 1333 69
rect 1367 35 1400 69
rect 1300 1 1400 35
rect 1300 -33 1333 1
rect 1367 -33 1400 1
rect 1300 -67 1400 -33
rect 1300 -101 1333 -67
rect 1367 -101 1400 -67
rect 1600 1300 2700 1400
rect 1600 0 1700 1300
rect 2600 0 2700 1300
rect 1600 -33 2700 0
rect 1600 -67 1623 -33
rect 1657 -67 1691 -33
rect 1725 -67 1759 -33
rect 1793 -67 1827 -33
rect 1861 -67 1895 -33
rect 1929 -67 1963 -33
rect 1997 -67 2031 -33
rect 2065 -67 2099 -33
rect 2133 -67 2167 -33
rect 2201 -67 2235 -33
rect 2269 -67 2303 -33
rect 2337 -67 2371 -33
rect 2405 -67 2439 -33
rect 2473 -67 2507 -33
rect 2541 -67 2575 -33
rect 2609 -67 2643 -33
rect 2677 -67 2700 -33
rect 1600 -100 2700 -67
rect 2800 1300 3900 1400
rect 2800 0 2900 1300
rect 3800 0 3900 1300
rect 2800 -33 3900 0
rect 2800 -67 2823 -33
rect 2857 -67 2891 -33
rect 2925 -67 2959 -33
rect 2993 -67 3027 -33
rect 3061 -67 3095 -33
rect 3129 -67 3163 -33
rect 3197 -67 3231 -33
rect 3265 -67 3299 -33
rect 3333 -67 3367 -33
rect 3401 -67 3435 -33
rect 3469 -67 3503 -33
rect 3537 -67 3571 -33
rect 3605 -67 3639 -33
rect 3673 -67 3707 -33
rect 3741 -67 3775 -33
rect 3809 -67 3843 -33
rect 3877 -67 3900 -33
rect 2800 -100 3900 -67
rect 4300 1300 5400 1400
rect 4300 0 4400 1300
rect 5300 0 5400 1300
rect 4300 -33 5400 0
rect 4300 -67 4323 -33
rect 4357 -67 4391 -33
rect 4425 -67 4459 -33
rect 4493 -67 4527 -33
rect 4561 -67 4595 -33
rect 4629 -67 4663 -33
rect 4697 -67 4731 -33
rect 4765 -67 4799 -33
rect 4833 -67 4867 -33
rect 4901 -67 4935 -33
rect 4969 -67 5003 -33
rect 5037 -67 5071 -33
rect 5105 -67 5139 -33
rect 5173 -67 5207 -33
rect 5241 -67 5275 -33
rect 5309 -67 5343 -33
rect 5377 -67 5400 -33
rect 4300 -100 5400 -67
rect 5500 1300 6600 1400
rect 5500 0 5600 1300
rect 6500 0 6600 1300
rect 5500 -33 6600 0
rect 5500 -67 5523 -33
rect 5557 -67 5591 -33
rect 5625 -67 5659 -33
rect 5693 -67 5727 -33
rect 5761 -67 5795 -33
rect 5829 -67 5863 -33
rect 5897 -67 5931 -33
rect 5965 -67 5999 -33
rect 6033 -67 6067 -33
rect 6101 -67 6135 -33
rect 6169 -67 6203 -33
rect 6237 -67 6271 -33
rect 6305 -67 6339 -33
rect 6373 -67 6407 -33
rect 6441 -67 6475 -33
rect 6509 -67 6543 -33
rect 6577 -67 6600 -33
rect 5500 -100 6600 -67
rect 6800 1390 6833 1424
rect 6867 1390 6900 1424
rect 6800 1356 6900 1390
rect 6800 1322 6833 1356
rect 6867 1322 6900 1356
rect 6800 1288 6900 1322
rect 6800 1254 6833 1288
rect 6867 1254 6900 1288
rect 6800 1220 6900 1254
rect 6800 1186 6833 1220
rect 6867 1186 6900 1220
rect 6800 1152 6900 1186
rect 6800 1118 6833 1152
rect 6867 1118 6900 1152
rect 6800 1084 6900 1118
rect 6800 1050 6833 1084
rect 6867 1050 6900 1084
rect 6800 1016 6900 1050
rect 6800 982 6833 1016
rect 6867 982 6900 1016
rect 6800 948 6900 982
rect 6800 914 6833 948
rect 6867 914 6900 948
rect 6800 880 6900 914
rect 6800 846 6833 880
rect 6867 846 6900 880
rect 6800 812 6900 846
rect 6800 778 6833 812
rect 6867 778 6900 812
rect 6800 744 6900 778
rect 6800 710 6833 744
rect 6867 710 6900 744
rect 6800 676 6900 710
rect 6800 642 6833 676
rect 6867 642 6900 676
rect 6800 608 6900 642
rect 6800 574 6833 608
rect 6867 574 6900 608
rect 6800 540 6900 574
rect 6800 506 6833 540
rect 6867 506 6900 540
rect 6800 472 6900 506
rect 6800 438 6833 472
rect 6867 438 6900 472
rect 6800 404 6900 438
rect 6800 370 6833 404
rect 6867 370 6900 404
rect 6800 336 6900 370
rect 6800 302 6833 336
rect 6867 302 6900 336
rect 6800 268 6900 302
rect 6800 234 6833 268
rect 6867 234 6900 268
rect 6800 200 6900 234
rect 6800 166 6833 200
rect 6867 166 6900 200
rect 6800 132 6900 166
rect 6800 98 6833 132
rect 6867 98 6900 132
rect 6800 64 6900 98
rect 6800 30 6833 64
rect 6867 30 6900 64
rect 6800 -4 6900 30
rect 6800 -38 6833 -4
rect 6867 -38 6900 -4
rect 6800 -72 6900 -38
rect 1300 -135 1400 -101
rect 1300 -169 1333 -135
rect 1367 -169 1400 -135
rect 1300 -200 1400 -169
rect 6800 -106 6833 -72
rect 6867 -106 6900 -72
rect 6800 -140 6900 -106
rect 6800 -174 6833 -140
rect 6867 -174 6900 -140
rect 6800 -200 6900 -174
rect 1300 -233 6900 -200
rect 1300 -267 1431 -233
rect 1465 -267 1499 -233
rect 1533 -267 1567 -233
rect 1601 -267 1635 -233
rect 1669 -267 1703 -233
rect 1737 -267 1771 -233
rect 1805 -267 1839 -233
rect 1873 -267 1907 -233
rect 1941 -267 1975 -233
rect 2009 -267 2043 -233
rect 2077 -267 2111 -233
rect 2145 -267 2179 -233
rect 2213 -267 2247 -233
rect 2281 -267 2315 -233
rect 2349 -267 2383 -233
rect 2417 -267 2451 -233
rect 2485 -267 2519 -233
rect 2553 -267 2587 -233
rect 2621 -267 2655 -233
rect 2689 -267 2723 -233
rect 2757 -267 2791 -233
rect 2825 -267 2859 -233
rect 2893 -267 2927 -233
rect 2961 -267 2995 -233
rect 3029 -267 3063 -233
rect 3097 -267 3131 -233
rect 3165 -267 3199 -233
rect 3233 -267 3267 -233
rect 3301 -267 3335 -233
rect 3369 -267 3403 -233
rect 3437 -267 3471 -233
rect 3505 -267 3539 -233
rect 3573 -267 3607 -233
rect 3641 -267 3675 -233
rect 3709 -267 3743 -233
rect 3777 -267 3811 -233
rect 3845 -267 3879 -233
rect 3913 -267 3947 -233
rect 3981 -267 4015 -233
rect 4049 -267 4083 -233
rect 4117 -267 4151 -233
rect 4185 -267 4219 -233
rect 4253 -267 4287 -233
rect 4321 -267 4355 -233
rect 4389 -267 4423 -233
rect 4457 -267 4491 -233
rect 4525 -267 4559 -233
rect 4593 -267 4627 -233
rect 4661 -267 4695 -233
rect 4729 -267 4763 -233
rect 4797 -267 4831 -233
rect 4865 -267 4899 -233
rect 4933 -267 4967 -233
rect 5001 -267 5035 -233
rect 5069 -267 5103 -233
rect 5137 -267 5171 -233
rect 5205 -267 5239 -233
rect 5273 -267 5307 -233
rect 5341 -267 5375 -233
rect 5409 -267 5443 -233
rect 5477 -267 5511 -233
rect 5545 -267 5579 -233
rect 5613 -267 5647 -233
rect 5681 -267 5715 -233
rect 5749 -267 5783 -233
rect 5817 -267 5851 -233
rect 5885 -267 5919 -233
rect 5953 -267 5987 -233
rect 6021 -267 6055 -233
rect 6089 -267 6123 -233
rect 6157 -267 6191 -233
rect 6225 -267 6259 -233
rect 6293 -267 6327 -233
rect 6361 -267 6395 -233
rect 6429 -267 6463 -233
rect 6497 -267 6531 -233
rect 6565 -267 6599 -233
rect 6633 -267 6667 -233
rect 6701 -267 6735 -233
rect 6769 -267 6900 -233
rect 1300 -300 6900 -267
<< psubdiffcont >>
rect 1441 3533 1475 3567
rect 1509 3533 1543 3567
rect 1577 3533 1611 3567
rect 1645 3533 1679 3567
rect 1713 3533 1747 3567
rect 1781 3533 1815 3567
rect 1849 3533 1883 3567
rect 1917 3533 1951 3567
rect 1985 3533 2019 3567
rect 2053 3533 2087 3567
rect 2121 3533 2155 3567
rect 2189 3533 2223 3567
rect 2257 3533 2291 3567
rect 2325 3533 2359 3567
rect 2393 3533 2427 3567
rect 2461 3533 2495 3567
rect 2529 3533 2563 3567
rect 2597 3533 2631 3567
rect 2665 3533 2699 3567
rect 2733 3533 2767 3567
rect 2801 3533 2835 3567
rect 2869 3533 2903 3567
rect 2937 3533 2971 3567
rect 3005 3533 3039 3567
rect 3073 3533 3107 3567
rect 3141 3533 3175 3567
rect 3209 3533 3243 3567
rect 3277 3533 3311 3567
rect 3345 3533 3379 3567
rect 3413 3533 3447 3567
rect 3481 3533 3515 3567
rect 3549 3533 3583 3567
rect 3617 3533 3651 3567
rect 3685 3533 3719 3567
rect 3753 3533 3787 3567
rect 3821 3533 3855 3567
rect 3889 3533 3923 3567
rect 3957 3533 3991 3567
rect 4025 3533 4059 3567
rect 4093 3533 4127 3567
rect 4161 3533 4195 3567
rect 4229 3533 4263 3567
rect 4297 3533 4331 3567
rect 4365 3533 4399 3567
rect 4433 3533 4467 3567
rect 4501 3533 4535 3567
rect 4569 3533 4603 3567
rect 4637 3533 4671 3567
rect 4705 3533 4739 3567
rect 4773 3533 4807 3567
rect 4841 3533 4875 3567
rect 4909 3533 4943 3567
rect 4977 3533 5011 3567
rect 5045 3533 5079 3567
rect 5113 3533 5147 3567
rect 5181 3533 5215 3567
rect 5249 3533 5283 3567
rect 5317 3533 5351 3567
rect 5385 3533 5419 3567
rect 5453 3533 5487 3567
rect 5521 3533 5555 3567
rect 5589 3533 5623 3567
rect 5657 3533 5691 3567
rect 5725 3533 5759 3567
rect 5793 3533 5827 3567
rect 5861 3533 5895 3567
rect 5929 3533 5963 3567
rect 5997 3533 6031 3567
rect 6065 3533 6099 3567
rect 6133 3533 6167 3567
rect 6201 3533 6235 3567
rect 6269 3533 6303 3567
rect 6337 3533 6371 3567
rect 6405 3533 6439 3567
rect 6473 3533 6507 3567
rect 6541 3533 6575 3567
rect 6609 3533 6643 3567
rect 6677 3533 6711 3567
rect 6745 3533 6779 3567
rect 1333 3435 1367 3469
rect 1333 3367 1367 3401
rect 6833 3430 6867 3464
rect 1333 3299 1367 3333
rect 1333 3231 1367 3265
rect 1333 3163 1367 3197
rect 1333 3095 1367 3129
rect 1333 3027 1367 3061
rect 1333 2959 1367 2993
rect 1333 2891 1367 2925
rect 1333 2823 1367 2857
rect 1333 2755 1367 2789
rect 1333 2687 1367 2721
rect 1333 2619 1367 2653
rect 1333 2551 1367 2585
rect 1333 2483 1367 2517
rect 1333 2415 1367 2449
rect 1333 2347 1367 2381
rect 1333 2279 1367 2313
rect 1333 2211 1367 2245
rect 1333 2143 1367 2177
rect 1333 2075 1367 2109
rect 1333 2007 1367 2041
rect 1333 1939 1367 1973
rect 1333 1871 1367 1905
rect 1623 3333 1657 3367
rect 1691 3333 1725 3367
rect 1759 3333 1793 3367
rect 1827 3333 1861 3367
rect 1895 3333 1929 3367
rect 1963 3333 1997 3367
rect 2031 3333 2065 3367
rect 2099 3333 2133 3367
rect 2167 3333 2201 3367
rect 2235 3333 2269 3367
rect 2303 3333 2337 3367
rect 2371 3333 2405 3367
rect 2439 3333 2473 3367
rect 2507 3333 2541 3367
rect 2575 3333 2609 3367
rect 2643 3333 2677 3367
rect 2823 3333 2857 3367
rect 2891 3333 2925 3367
rect 2959 3333 2993 3367
rect 3027 3333 3061 3367
rect 3095 3333 3129 3367
rect 3163 3333 3197 3367
rect 3231 3333 3265 3367
rect 3299 3333 3333 3367
rect 3367 3333 3401 3367
rect 3435 3333 3469 3367
rect 3503 3333 3537 3367
rect 3571 3333 3605 3367
rect 3639 3333 3673 3367
rect 3707 3333 3741 3367
rect 3775 3333 3809 3367
rect 3843 3333 3877 3367
rect 4323 3333 4357 3367
rect 4391 3333 4425 3367
rect 4459 3333 4493 3367
rect 4527 3333 4561 3367
rect 4595 3333 4629 3367
rect 4663 3333 4697 3367
rect 4731 3333 4765 3367
rect 4799 3333 4833 3367
rect 4867 3333 4901 3367
rect 4935 3333 4969 3367
rect 5003 3333 5037 3367
rect 5071 3333 5105 3367
rect 5139 3333 5173 3367
rect 5207 3333 5241 3367
rect 5275 3333 5309 3367
rect 5343 3333 5377 3367
rect 5523 3333 5557 3367
rect 5591 3333 5625 3367
rect 5659 3333 5693 3367
rect 5727 3333 5761 3367
rect 5795 3333 5829 3367
rect 5863 3333 5897 3367
rect 5931 3333 5965 3367
rect 5999 3333 6033 3367
rect 6067 3333 6101 3367
rect 6135 3333 6169 3367
rect 6203 3333 6237 3367
rect 6271 3333 6305 3367
rect 6339 3333 6373 3367
rect 6407 3333 6441 3367
rect 6475 3333 6509 3367
rect 6543 3333 6577 3367
rect 6833 3362 6867 3396
rect 6833 3294 6867 3328
rect 6833 3226 6867 3260
rect 6833 3158 6867 3192
rect 6833 3090 6867 3124
rect 6833 3022 6867 3056
rect 6833 2954 6867 2988
rect 6833 2886 6867 2920
rect 6833 2818 6867 2852
rect 6833 2750 6867 2784
rect 6833 2682 6867 2716
rect 6833 2614 6867 2648
rect 6833 2546 6867 2580
rect 6833 2478 6867 2512
rect 6833 2410 6867 2444
rect 6833 2342 6867 2376
rect 6833 2274 6867 2308
rect 6833 2206 6867 2240
rect 6833 2138 6867 2172
rect 6833 2070 6867 2104
rect 6833 2002 6867 2036
rect 6833 1934 6867 1968
rect 1333 1803 1367 1837
rect 1333 1735 1367 1769
rect 1333 1667 1367 1701
rect 1333 1599 1367 1633
rect 1333 1531 1367 1565
rect 1333 1463 1367 1497
rect 1333 1395 1367 1429
rect 6833 1866 6867 1900
rect 6833 1798 6867 1832
rect 6833 1730 6867 1764
rect 6833 1662 6867 1696
rect 6833 1594 6867 1628
rect 6833 1526 6867 1560
rect 6833 1458 6867 1492
rect 1333 1327 1367 1361
rect 1333 1259 1367 1293
rect 1333 1191 1367 1225
rect 1333 1123 1367 1157
rect 1333 1055 1367 1089
rect 1333 987 1367 1021
rect 1333 919 1367 953
rect 1333 851 1367 885
rect 1333 783 1367 817
rect 1333 715 1367 749
rect 1333 647 1367 681
rect 1333 579 1367 613
rect 1333 511 1367 545
rect 1333 443 1367 477
rect 1333 375 1367 409
rect 1333 307 1367 341
rect 1333 239 1367 273
rect 1333 171 1367 205
rect 1333 103 1367 137
rect 1333 35 1367 69
rect 1333 -33 1367 1
rect 1333 -101 1367 -67
rect 1623 -67 1657 -33
rect 1691 -67 1725 -33
rect 1759 -67 1793 -33
rect 1827 -67 1861 -33
rect 1895 -67 1929 -33
rect 1963 -67 1997 -33
rect 2031 -67 2065 -33
rect 2099 -67 2133 -33
rect 2167 -67 2201 -33
rect 2235 -67 2269 -33
rect 2303 -67 2337 -33
rect 2371 -67 2405 -33
rect 2439 -67 2473 -33
rect 2507 -67 2541 -33
rect 2575 -67 2609 -33
rect 2643 -67 2677 -33
rect 2823 -67 2857 -33
rect 2891 -67 2925 -33
rect 2959 -67 2993 -33
rect 3027 -67 3061 -33
rect 3095 -67 3129 -33
rect 3163 -67 3197 -33
rect 3231 -67 3265 -33
rect 3299 -67 3333 -33
rect 3367 -67 3401 -33
rect 3435 -67 3469 -33
rect 3503 -67 3537 -33
rect 3571 -67 3605 -33
rect 3639 -67 3673 -33
rect 3707 -67 3741 -33
rect 3775 -67 3809 -33
rect 3843 -67 3877 -33
rect 4323 -67 4357 -33
rect 4391 -67 4425 -33
rect 4459 -67 4493 -33
rect 4527 -67 4561 -33
rect 4595 -67 4629 -33
rect 4663 -67 4697 -33
rect 4731 -67 4765 -33
rect 4799 -67 4833 -33
rect 4867 -67 4901 -33
rect 4935 -67 4969 -33
rect 5003 -67 5037 -33
rect 5071 -67 5105 -33
rect 5139 -67 5173 -33
rect 5207 -67 5241 -33
rect 5275 -67 5309 -33
rect 5343 -67 5377 -33
rect 5523 -67 5557 -33
rect 5591 -67 5625 -33
rect 5659 -67 5693 -33
rect 5727 -67 5761 -33
rect 5795 -67 5829 -33
rect 5863 -67 5897 -33
rect 5931 -67 5965 -33
rect 5999 -67 6033 -33
rect 6067 -67 6101 -33
rect 6135 -67 6169 -33
rect 6203 -67 6237 -33
rect 6271 -67 6305 -33
rect 6339 -67 6373 -33
rect 6407 -67 6441 -33
rect 6475 -67 6509 -33
rect 6543 -67 6577 -33
rect 6833 1390 6867 1424
rect 6833 1322 6867 1356
rect 6833 1254 6867 1288
rect 6833 1186 6867 1220
rect 6833 1118 6867 1152
rect 6833 1050 6867 1084
rect 6833 982 6867 1016
rect 6833 914 6867 948
rect 6833 846 6867 880
rect 6833 778 6867 812
rect 6833 710 6867 744
rect 6833 642 6867 676
rect 6833 574 6867 608
rect 6833 506 6867 540
rect 6833 438 6867 472
rect 6833 370 6867 404
rect 6833 302 6867 336
rect 6833 234 6867 268
rect 6833 166 6867 200
rect 6833 98 6867 132
rect 6833 30 6867 64
rect 6833 -38 6867 -4
rect 1333 -169 1367 -135
rect 6833 -106 6867 -72
rect 6833 -174 6867 -140
rect 1431 -267 1465 -233
rect 1499 -267 1533 -233
rect 1567 -267 1601 -233
rect 1635 -267 1669 -233
rect 1703 -267 1737 -233
rect 1771 -267 1805 -233
rect 1839 -267 1873 -233
rect 1907 -267 1941 -233
rect 1975 -267 2009 -233
rect 2043 -267 2077 -233
rect 2111 -267 2145 -233
rect 2179 -267 2213 -233
rect 2247 -267 2281 -233
rect 2315 -267 2349 -233
rect 2383 -267 2417 -233
rect 2451 -267 2485 -233
rect 2519 -267 2553 -233
rect 2587 -267 2621 -233
rect 2655 -267 2689 -233
rect 2723 -267 2757 -233
rect 2791 -267 2825 -233
rect 2859 -267 2893 -233
rect 2927 -267 2961 -233
rect 2995 -267 3029 -233
rect 3063 -267 3097 -233
rect 3131 -267 3165 -233
rect 3199 -267 3233 -233
rect 3267 -267 3301 -233
rect 3335 -267 3369 -233
rect 3403 -267 3437 -233
rect 3471 -267 3505 -233
rect 3539 -267 3573 -233
rect 3607 -267 3641 -233
rect 3675 -267 3709 -233
rect 3743 -267 3777 -233
rect 3811 -267 3845 -233
rect 3879 -267 3913 -233
rect 3947 -267 3981 -233
rect 4015 -267 4049 -233
rect 4083 -267 4117 -233
rect 4151 -267 4185 -233
rect 4219 -267 4253 -233
rect 4287 -267 4321 -233
rect 4355 -267 4389 -233
rect 4423 -267 4457 -233
rect 4491 -267 4525 -233
rect 4559 -267 4593 -233
rect 4627 -267 4661 -233
rect 4695 -267 4729 -233
rect 4763 -267 4797 -233
rect 4831 -267 4865 -233
rect 4899 -267 4933 -233
rect 4967 -267 5001 -233
rect 5035 -267 5069 -233
rect 5103 -267 5137 -233
rect 5171 -267 5205 -233
rect 5239 -267 5273 -233
rect 5307 -267 5341 -233
rect 5375 -267 5409 -233
rect 5443 -267 5477 -233
rect 5511 -267 5545 -233
rect 5579 -267 5613 -233
rect 5647 -267 5681 -233
rect 5715 -267 5749 -233
rect 5783 -267 5817 -233
rect 5851 -267 5885 -233
rect 5919 -267 5953 -233
rect 5987 -267 6021 -233
rect 6055 -267 6089 -233
rect 6123 -267 6157 -233
rect 6191 -267 6225 -233
rect 6259 -267 6293 -233
rect 6327 -267 6361 -233
rect 6395 -267 6429 -233
rect 6463 -267 6497 -233
rect 6531 -267 6565 -233
rect 6599 -267 6633 -233
rect 6667 -267 6701 -233
rect 6735 -267 6769 -233
<< poly >>
rect 1720 2100 1780 3120
rect 2510 2100 2570 3120
rect 2920 2100 2980 3120
rect 3710 2090 3770 3110
rect 4420 2100 4480 3120
rect 5210 2100 5270 3120
rect 5620 2100 5680 3120
rect 6410 2100 6470 3120
rect 1720 200 1780 1220
rect 2510 200 2570 1220
rect 2920 200 2980 1220
rect 3720 200 3780 1220
rect 4420 200 4480 1200
rect 5210 200 5270 1200
rect 5620 200 5680 1200
rect 6410 210 6470 1210
<< locali >>
rect 1300 3567 6900 3600
rect 1300 3533 1441 3567
rect 1475 3533 1509 3567
rect 1543 3533 1577 3567
rect 1611 3533 1645 3567
rect 1679 3533 1713 3567
rect 1747 3533 1781 3567
rect 1815 3533 1849 3567
rect 1883 3533 1917 3567
rect 1951 3533 1985 3567
rect 2019 3533 2053 3567
rect 2087 3533 2121 3567
rect 2155 3533 2189 3567
rect 2223 3533 2257 3567
rect 2291 3533 2325 3567
rect 2359 3533 2393 3567
rect 2427 3533 2461 3567
rect 2495 3533 2529 3567
rect 2563 3533 2597 3567
rect 2631 3533 2665 3567
rect 2699 3533 2733 3567
rect 2767 3533 2801 3567
rect 2835 3533 2869 3567
rect 2903 3533 2937 3567
rect 2971 3533 3005 3567
rect 3039 3533 3073 3567
rect 3107 3533 3141 3567
rect 3175 3533 3209 3567
rect 3243 3533 3277 3567
rect 3311 3533 3345 3567
rect 3379 3533 3413 3567
rect 3447 3533 3481 3567
rect 3515 3533 3549 3567
rect 3583 3533 3617 3567
rect 3651 3533 3685 3567
rect 3719 3533 3753 3567
rect 3787 3533 3821 3567
rect 3855 3533 3889 3567
rect 3923 3533 3957 3567
rect 3991 3533 4025 3567
rect 4059 3533 4093 3567
rect 4127 3533 4161 3567
rect 4195 3533 4229 3567
rect 4263 3533 4297 3567
rect 4331 3533 4365 3567
rect 4399 3533 4433 3567
rect 4467 3533 4501 3567
rect 4535 3533 4569 3567
rect 4603 3533 4637 3567
rect 4671 3533 4705 3567
rect 4739 3533 4773 3567
rect 4807 3533 4841 3567
rect 4875 3533 4909 3567
rect 4943 3533 4977 3567
rect 5011 3533 5045 3567
rect 5079 3533 5113 3567
rect 5147 3533 5181 3567
rect 5215 3533 5249 3567
rect 5283 3533 5317 3567
rect 5351 3533 5385 3567
rect 5419 3533 5453 3567
rect 5487 3533 5521 3567
rect 5555 3533 5589 3567
rect 5623 3533 5657 3567
rect 5691 3533 5725 3567
rect 5759 3533 5793 3567
rect 5827 3533 5861 3567
rect 5895 3533 5929 3567
rect 5963 3533 5997 3567
rect 6031 3533 6065 3567
rect 6099 3533 6133 3567
rect 6167 3533 6201 3567
rect 6235 3533 6269 3567
rect 6303 3533 6337 3567
rect 6371 3533 6405 3567
rect 6439 3533 6473 3567
rect 6507 3533 6541 3567
rect 6575 3533 6609 3567
rect 6643 3533 6677 3567
rect 6711 3533 6745 3567
rect 6779 3533 6900 3567
rect 1300 3500 6900 3533
rect 1300 3469 1400 3500
rect 1300 3435 1333 3469
rect 1367 3435 1400 3469
rect 1300 3402 1400 3435
rect 6800 3464 6900 3500
rect 6800 3430 6833 3464
rect 6867 3430 6900 3464
rect 6800 3402 6900 3430
rect 1300 3401 1720 3402
rect 1300 3367 1333 3401
rect 1367 3400 1720 3401
rect 6480 3400 6900 3402
rect 1367 3367 3900 3400
rect 1300 3333 1623 3367
rect 1657 3333 1691 3367
rect 1725 3333 1759 3367
rect 1793 3333 1827 3367
rect 1861 3333 1895 3367
rect 1929 3333 1963 3367
rect 1997 3333 2031 3367
rect 2065 3333 2099 3367
rect 2133 3333 2167 3367
rect 2201 3333 2235 3367
rect 2269 3333 2303 3367
rect 2337 3333 2371 3367
rect 2405 3333 2439 3367
rect 2473 3333 2507 3367
rect 2541 3333 2575 3367
rect 2609 3333 2643 3367
rect 2677 3333 2823 3367
rect 2857 3333 2891 3367
rect 2925 3333 2959 3367
rect 2993 3333 3027 3367
rect 3061 3333 3095 3367
rect 3129 3333 3163 3367
rect 3197 3333 3231 3367
rect 3265 3333 3299 3367
rect 3333 3333 3367 3367
rect 3401 3333 3435 3367
rect 3469 3333 3503 3367
rect 3537 3333 3571 3367
rect 3605 3333 3639 3367
rect 3673 3333 3707 3367
rect 3741 3333 3775 3367
rect 3809 3333 3843 3367
rect 3877 3333 3900 3367
rect 1300 3299 1333 3333
rect 1367 3300 3900 3333
rect 3960 3347 4240 3400
rect 3960 3313 4033 3347
rect 4067 3313 4133 3347
rect 4167 3313 4240 3347
rect 1367 3299 1400 3300
rect 1300 3265 1400 3299
rect 1300 3231 1333 3265
rect 1367 3231 1400 3265
rect 3960 3260 4240 3313
rect 4300 3396 6900 3400
rect 4300 3367 6833 3396
rect 4300 3333 4323 3367
rect 4357 3333 4391 3367
rect 4425 3333 4459 3367
rect 4493 3333 4527 3367
rect 4561 3333 4595 3367
rect 4629 3333 4663 3367
rect 4697 3333 4731 3367
rect 4765 3333 4799 3367
rect 4833 3333 4867 3367
rect 4901 3333 4935 3367
rect 4969 3333 5003 3367
rect 5037 3333 5071 3367
rect 5105 3333 5139 3367
rect 5173 3333 5207 3367
rect 5241 3333 5275 3367
rect 5309 3333 5343 3367
rect 5377 3333 5523 3367
rect 5557 3333 5591 3367
rect 5625 3333 5659 3367
rect 5693 3333 5727 3367
rect 5761 3333 5795 3367
rect 5829 3333 5863 3367
rect 5897 3333 5931 3367
rect 5965 3333 5999 3367
rect 6033 3333 6067 3367
rect 6101 3333 6135 3367
rect 6169 3333 6203 3367
rect 6237 3333 6271 3367
rect 6305 3333 6339 3367
rect 6373 3333 6407 3367
rect 6441 3333 6475 3367
rect 6509 3333 6543 3367
rect 6577 3362 6833 3367
rect 6867 3362 6900 3396
rect 6577 3333 6900 3362
rect 4300 3328 6900 3333
rect 4300 3300 6833 3328
rect 6800 3294 6833 3300
rect 6867 3294 6900 3328
rect 6800 3260 6900 3294
rect 1300 3197 1400 3231
rect 1300 3163 1333 3197
rect 1367 3163 1400 3197
rect 1300 3129 1400 3163
rect 3000 3247 5200 3260
rect 3000 3213 4033 3247
rect 4067 3213 4133 3247
rect 4167 3213 5200 3247
rect 3000 3160 5200 3213
rect 6800 3226 6833 3260
rect 6867 3226 6900 3260
rect 6800 3192 6900 3226
rect 1300 3095 1333 3129
rect 1367 3095 1400 3129
rect 1300 3061 1400 3095
rect 1300 3027 1333 3061
rect 1367 3027 1400 3061
rect 1300 2993 1400 3027
rect 1300 2959 1333 2993
rect 1367 2959 1400 2993
rect 1300 2925 1400 2959
rect 1300 2891 1333 2925
rect 1367 2891 1400 2925
rect 1300 2857 1400 2891
rect 1300 2823 1333 2857
rect 1367 2823 1400 2857
rect 1300 2789 1400 2823
rect 1300 2755 1333 2789
rect 1367 2755 1400 2789
rect 1300 2721 1400 2755
rect 1300 2687 1333 2721
rect 1367 2687 1400 2721
rect 1300 2653 1400 2687
rect 1300 2619 1333 2653
rect 1367 2619 1400 2653
rect 1300 2585 1400 2619
rect 1300 2551 1333 2585
rect 1367 2551 1400 2585
rect 1300 2517 1400 2551
rect 1300 2483 1333 2517
rect 1367 2483 1400 2517
rect 1300 2449 1400 2483
rect 1300 2415 1333 2449
rect 1367 2415 1400 2449
rect 1300 2381 1400 2415
rect 1300 2347 1333 2381
rect 1367 2347 1400 2381
rect 1300 2313 1400 2347
rect 1300 2279 1333 2313
rect 1367 2279 1400 2313
rect 1300 2245 1400 2279
rect 1300 2211 1333 2245
rect 1367 2211 1400 2245
rect 1300 2177 1400 2211
rect 1300 2143 1333 2177
rect 1367 2143 1400 2177
rect 1300 2109 1400 2143
rect 1300 2075 1333 2109
rect 1367 2075 1400 2109
rect 1300 2041 1400 2075
rect 1300 2007 1333 2041
rect 1367 2007 1400 2041
rect 1300 1973 1400 2007
rect 1300 1939 1333 1973
rect 1367 1939 1400 1973
rect 1300 1905 1400 1939
rect 1300 1871 1333 1905
rect 1367 1871 1400 1905
rect 1300 1837 1400 1871
rect 1300 1803 1333 1837
rect 1367 1803 1400 1837
rect 1300 1769 1400 1803
rect 2080 1800 2200 3020
rect 3280 2200 3400 3160
rect 3900 3147 4300 3160
rect 3900 3113 4033 3147
rect 4067 3113 4133 3147
rect 4167 3113 4300 3147
rect 3900 3047 4300 3113
rect 3900 3013 4033 3047
rect 4067 3013 4133 3047
rect 4167 3013 4300 3047
rect 3900 2947 4300 3013
rect 3900 2913 4033 2947
rect 4067 2913 4133 2947
rect 4167 2913 4300 2947
rect 3900 2847 4300 2913
rect 3900 2813 4033 2847
rect 4067 2813 4133 2847
rect 4167 2813 4300 2847
rect 3900 2747 4300 2813
rect 3900 2713 4033 2747
rect 4067 2713 4133 2747
rect 4167 2713 4300 2747
rect 3900 2647 4300 2713
rect 3900 2613 4033 2647
rect 4067 2613 4133 2647
rect 4167 2613 4300 2647
rect 3900 2547 4300 2613
rect 3900 2513 4033 2547
rect 4067 2513 4133 2547
rect 4167 2513 4300 2547
rect 3900 2447 4300 2513
rect 3900 2413 4033 2447
rect 4067 2413 4133 2447
rect 4167 2413 4300 2447
rect 3900 2347 4300 2413
rect 3900 2313 4033 2347
rect 4067 2313 4133 2347
rect 4167 2313 4300 2347
rect 3900 2247 4300 2313
rect 3900 2213 4033 2247
rect 4067 2213 4133 2247
rect 4167 2213 4300 2247
rect 3900 2147 4300 2213
rect 4780 2200 4900 3160
rect 6800 3158 6833 3192
rect 6867 3158 6900 3192
rect 6800 3124 6900 3158
rect 6800 3090 6833 3124
rect 6867 3090 6900 3124
rect 6800 3056 6900 3090
rect 6800 3022 6833 3056
rect 6867 3022 6900 3056
rect 3900 2113 4033 2147
rect 4067 2113 4133 2147
rect 4167 2113 4300 2147
rect 3900 1800 4300 2113
rect 5980 1800 6100 3020
rect 6800 2988 6900 3022
rect 6800 2954 6833 2988
rect 6867 2954 6900 2988
rect 6800 2920 6900 2954
rect 6800 2886 6833 2920
rect 6867 2886 6900 2920
rect 6800 2852 6900 2886
rect 6800 2818 6833 2852
rect 6867 2818 6900 2852
rect 6800 2784 6900 2818
rect 6800 2750 6833 2784
rect 6867 2750 6900 2784
rect 6800 2716 6900 2750
rect 6800 2682 6833 2716
rect 6867 2682 6900 2716
rect 6800 2648 6900 2682
rect 6800 2614 6833 2648
rect 6867 2614 6900 2648
rect 6800 2580 6900 2614
rect 6800 2546 6833 2580
rect 6867 2546 6900 2580
rect 6800 2512 6900 2546
rect 6800 2478 6833 2512
rect 6867 2478 6900 2512
rect 6800 2444 6900 2478
rect 6800 2410 6833 2444
rect 6867 2410 6900 2444
rect 6800 2376 6900 2410
rect 6800 2342 6833 2376
rect 6867 2342 6900 2376
rect 6800 2308 6900 2342
rect 6800 2274 6833 2308
rect 6867 2274 6900 2308
rect 6800 2240 6900 2274
rect 6800 2206 6833 2240
rect 6867 2206 6900 2240
rect 6800 2172 6900 2206
rect 6800 2138 6833 2172
rect 6867 2138 6900 2172
rect 6800 2104 6900 2138
rect 6800 2070 6833 2104
rect 6867 2070 6900 2104
rect 6800 2036 6900 2070
rect 6800 2002 6833 2036
rect 6867 2002 6900 2036
rect 6800 1968 6900 2002
rect 6800 1934 6833 1968
rect 6867 1934 6900 1968
rect 6800 1900 6900 1934
rect 6800 1866 6833 1900
rect 6867 1866 6900 1900
rect 6800 1832 6900 1866
rect 1300 1735 1333 1769
rect 1367 1735 1400 1769
rect 1300 1701 1400 1735
rect 1300 1667 1333 1701
rect 1367 1667 1400 1701
rect 1300 1633 1400 1667
rect 1300 1599 1333 1633
rect 1367 1599 1400 1633
rect 1300 1565 1400 1599
rect 1300 1531 1333 1565
rect 1367 1531 1400 1565
rect 1300 1497 1400 1531
rect 1500 1727 6700 1800
rect 1500 1693 1533 1727
rect 1567 1693 1633 1727
rect 1667 1693 1733 1727
rect 1767 1693 1833 1727
rect 1867 1693 1933 1727
rect 1967 1693 2033 1727
rect 2067 1693 2133 1727
rect 2167 1693 2233 1727
rect 2267 1693 2333 1727
rect 2367 1693 2433 1727
rect 2467 1693 2533 1727
rect 2567 1693 2633 1727
rect 2667 1693 2733 1727
rect 2767 1693 2833 1727
rect 2867 1693 2933 1727
rect 2967 1693 3033 1727
rect 3067 1693 3133 1727
rect 3167 1693 3233 1727
rect 3267 1693 3333 1727
rect 3367 1693 3433 1727
rect 3467 1693 3533 1727
rect 3567 1693 3633 1727
rect 3667 1693 3733 1727
rect 3767 1693 3833 1727
rect 3867 1693 3933 1727
rect 3967 1693 4033 1727
rect 4067 1693 4133 1727
rect 4167 1693 4233 1727
rect 4267 1693 4333 1727
rect 4367 1693 4433 1727
rect 4467 1693 4533 1727
rect 4567 1693 4633 1727
rect 4667 1693 4733 1727
rect 4767 1693 4833 1727
rect 4867 1693 4933 1727
rect 4967 1693 5033 1727
rect 5067 1693 5133 1727
rect 5167 1693 5233 1727
rect 5267 1693 5333 1727
rect 5367 1693 5433 1727
rect 5467 1693 5533 1727
rect 5567 1693 5633 1727
rect 5667 1693 5733 1727
rect 5767 1693 5833 1727
rect 5867 1693 5933 1727
rect 5967 1693 6033 1727
rect 6067 1693 6133 1727
rect 6167 1693 6233 1727
rect 6267 1693 6333 1727
rect 6367 1693 6433 1727
rect 6467 1693 6533 1727
rect 6567 1693 6633 1727
rect 6667 1693 6700 1727
rect 1500 1607 6700 1693
rect 1500 1573 1533 1607
rect 1567 1573 1633 1607
rect 1667 1573 1733 1607
rect 1767 1573 1833 1607
rect 1867 1573 1933 1607
rect 1967 1573 2033 1607
rect 2067 1573 2133 1607
rect 2167 1573 2233 1607
rect 2267 1573 2333 1607
rect 2367 1573 2433 1607
rect 2467 1573 2533 1607
rect 2567 1573 2633 1607
rect 2667 1573 2733 1607
rect 2767 1573 2833 1607
rect 2867 1573 2933 1607
rect 2967 1573 3033 1607
rect 3067 1573 3133 1607
rect 3167 1573 3233 1607
rect 3267 1573 3333 1607
rect 3367 1573 3433 1607
rect 3467 1573 3533 1607
rect 3567 1573 3633 1607
rect 3667 1573 3733 1607
rect 3767 1573 3833 1607
rect 3867 1573 3933 1607
rect 3967 1573 4033 1607
rect 4067 1573 4133 1607
rect 4167 1573 4233 1607
rect 4267 1573 4333 1607
rect 4367 1573 4433 1607
rect 4467 1573 4533 1607
rect 4567 1573 4633 1607
rect 4667 1573 4733 1607
rect 4767 1573 4833 1607
rect 4867 1573 4933 1607
rect 4967 1573 5033 1607
rect 5067 1573 5133 1607
rect 5167 1573 5233 1607
rect 5267 1573 5333 1607
rect 5367 1573 5433 1607
rect 5467 1573 5533 1607
rect 5567 1573 5633 1607
rect 5667 1573 5733 1607
rect 5767 1573 5833 1607
rect 5867 1573 5933 1607
rect 5967 1573 6033 1607
rect 6067 1573 6133 1607
rect 6167 1573 6233 1607
rect 6267 1573 6333 1607
rect 6367 1573 6433 1607
rect 6467 1573 6533 1607
rect 6567 1573 6633 1607
rect 6667 1573 6700 1607
rect 1500 1500 6700 1573
rect 6800 1798 6833 1832
rect 6867 1798 6900 1832
rect 6800 1764 6900 1798
rect 6800 1730 6833 1764
rect 6867 1730 6900 1764
rect 6800 1696 6900 1730
rect 6800 1662 6833 1696
rect 6867 1662 6900 1696
rect 6800 1628 6900 1662
rect 6800 1594 6833 1628
rect 6867 1594 6900 1628
rect 6800 1560 6900 1594
rect 6800 1526 6833 1560
rect 6867 1526 6900 1560
rect 1300 1463 1333 1497
rect 1367 1463 1400 1497
rect 1300 1429 1400 1463
rect 1300 1395 1333 1429
rect 1367 1395 1400 1429
rect 1300 1361 1400 1395
rect 1300 1327 1333 1361
rect 1367 1327 1400 1361
rect 1300 1293 1400 1327
rect 1300 1259 1333 1293
rect 1367 1259 1400 1293
rect 1300 1225 1400 1259
rect 1300 1191 1333 1225
rect 1367 1191 1400 1225
rect 1300 1157 1400 1191
rect 1300 1123 1333 1157
rect 1367 1123 1400 1157
rect 1300 1089 1400 1123
rect 1300 1055 1333 1089
rect 1367 1055 1400 1089
rect 1300 1021 1400 1055
rect 1300 987 1333 1021
rect 1367 987 1400 1021
rect 1300 953 1400 987
rect 1300 919 1333 953
rect 1367 919 1400 953
rect 1300 885 1400 919
rect 1300 851 1333 885
rect 1367 851 1400 885
rect 1300 817 1400 851
rect 1300 783 1333 817
rect 1367 783 1400 817
rect 1300 749 1400 783
rect 1300 715 1333 749
rect 1367 715 1400 749
rect 1300 681 1400 715
rect 1300 647 1333 681
rect 1367 647 1400 681
rect 1300 613 1400 647
rect 1300 579 1333 613
rect 1367 579 1400 613
rect 1300 545 1400 579
rect 1300 511 1333 545
rect 1367 511 1400 545
rect 1300 477 1400 511
rect 1300 443 1333 477
rect 1367 443 1400 477
rect 1300 409 1400 443
rect 1300 375 1333 409
rect 1367 375 1400 409
rect 1300 341 1400 375
rect 1300 307 1333 341
rect 1367 307 1400 341
rect 1300 273 1400 307
rect 2080 300 2200 1500
rect 3900 1187 4300 1500
rect 3900 1153 4033 1187
rect 4067 1153 4133 1187
rect 4167 1153 4300 1187
rect 1300 239 1333 273
rect 1367 239 1400 273
rect 1300 205 1400 239
rect 1300 171 1333 205
rect 1367 171 1400 205
rect 1300 137 1400 171
rect 3280 140 3400 1120
rect 3900 1087 4300 1153
rect 3900 1053 4033 1087
rect 4067 1053 4133 1087
rect 4167 1053 4300 1087
rect 3900 987 4300 1053
rect 3900 953 4033 987
rect 4067 953 4133 987
rect 4167 953 4300 987
rect 3900 887 4300 953
rect 3900 853 4033 887
rect 4067 853 4133 887
rect 4167 853 4300 887
rect 3900 787 4300 853
rect 3900 753 4033 787
rect 4067 753 4133 787
rect 4167 753 4300 787
rect 3900 687 4300 753
rect 3900 653 4033 687
rect 4067 653 4133 687
rect 4167 653 4300 687
rect 3900 587 4300 653
rect 3900 553 4033 587
rect 4067 553 4133 587
rect 4167 553 4300 587
rect 3900 487 4300 553
rect 3900 453 4033 487
rect 4067 453 4133 487
rect 4167 453 4300 487
rect 3900 387 4300 453
rect 3900 353 4033 387
rect 4067 353 4133 387
rect 4167 353 4300 387
rect 3900 287 4300 353
rect 3900 253 4033 287
rect 4067 253 4133 287
rect 4167 253 4300 287
rect 3900 187 4300 253
rect 3900 153 4033 187
rect 4067 153 4133 187
rect 4167 153 4300 187
rect 3900 140 4300 153
rect 4800 140 4920 1120
rect 5980 300 6100 1500
rect 6800 1492 6900 1526
rect 6800 1458 6833 1492
rect 6867 1458 6900 1492
rect 6800 1424 6900 1458
rect 6800 1390 6833 1424
rect 6867 1390 6900 1424
rect 6800 1356 6900 1390
rect 6800 1322 6833 1356
rect 6867 1322 6900 1356
rect 6800 1288 6900 1322
rect 6800 1254 6833 1288
rect 6867 1254 6900 1288
rect 6800 1220 6900 1254
rect 6800 1186 6833 1220
rect 6867 1186 6900 1220
rect 6800 1152 6900 1186
rect 6800 1118 6833 1152
rect 6867 1118 6900 1152
rect 6800 1084 6900 1118
rect 6800 1050 6833 1084
rect 6867 1050 6900 1084
rect 6800 1016 6900 1050
rect 6800 982 6833 1016
rect 6867 982 6900 1016
rect 6800 948 6900 982
rect 6800 914 6833 948
rect 6867 914 6900 948
rect 6800 880 6900 914
rect 6800 846 6833 880
rect 6867 846 6900 880
rect 6800 812 6900 846
rect 6800 778 6833 812
rect 6867 778 6900 812
rect 6800 744 6900 778
rect 6800 710 6833 744
rect 6867 710 6900 744
rect 6800 676 6900 710
rect 6800 642 6833 676
rect 6867 642 6900 676
rect 6800 608 6900 642
rect 6800 574 6833 608
rect 6867 574 6900 608
rect 6800 540 6900 574
rect 6800 506 6833 540
rect 6867 506 6900 540
rect 6800 472 6900 506
rect 6800 438 6833 472
rect 6867 438 6900 472
rect 6800 404 6900 438
rect 6800 370 6833 404
rect 6867 370 6900 404
rect 6800 336 6900 370
rect 6800 302 6833 336
rect 6867 302 6900 336
rect 6800 268 6900 302
rect 6800 234 6833 268
rect 6867 234 6900 268
rect 6800 200 6900 234
rect 6800 166 6833 200
rect 6867 166 6900 200
rect 1300 103 1333 137
rect 1367 103 1400 137
rect 1300 69 1400 103
rect 1300 35 1333 69
rect 1367 35 1400 69
rect 3000 87 5200 140
rect 3000 53 4033 87
rect 4067 53 4133 87
rect 4167 53 5200 87
rect 3000 40 5200 53
rect 6800 132 6900 166
rect 6800 98 6833 132
rect 6867 98 6900 132
rect 6800 64 6900 98
rect 1300 1 1400 35
rect 1300 -33 1333 1
rect 1367 0 1400 1
rect 1367 -33 3900 0
rect 1300 -67 1623 -33
rect 1657 -67 1691 -33
rect 1725 -67 1759 -33
rect 1793 -67 1827 -33
rect 1861 -67 1895 -33
rect 1929 -67 1963 -33
rect 1997 -67 2031 -33
rect 2065 -67 2099 -33
rect 2133 -67 2167 -33
rect 2201 -67 2235 -33
rect 2269 -67 2303 -33
rect 2337 -67 2371 -33
rect 2405 -67 2439 -33
rect 2473 -67 2507 -33
rect 2541 -67 2575 -33
rect 2609 -67 2643 -33
rect 2677 -67 2823 -33
rect 2857 -67 2891 -33
rect 2925 -67 2959 -33
rect 2993 -67 3027 -33
rect 3061 -67 3095 -33
rect 3129 -67 3163 -33
rect 3197 -67 3231 -33
rect 3265 -67 3299 -33
rect 3333 -67 3367 -33
rect 3401 -67 3435 -33
rect 3469 -67 3503 -33
rect 3537 -67 3571 -33
rect 3605 -67 3639 -33
rect 3673 -67 3707 -33
rect 3741 -67 3775 -33
rect 3809 -67 3843 -33
rect 3877 -67 3900 -33
rect 1300 -101 1333 -67
rect 1367 -100 3900 -67
rect 3960 -13 4240 40
rect 6800 30 6833 64
rect 6867 30 6900 64
rect 6800 2 6900 30
rect 6480 0 6900 2
rect 3960 -47 4033 -13
rect 4067 -47 4133 -13
rect 4167 -47 4240 -13
rect 3960 -100 4240 -47
rect 4300 -4 6900 0
rect 4300 -33 6833 -4
rect 4300 -67 4323 -33
rect 4357 -67 4391 -33
rect 4425 -67 4459 -33
rect 4493 -67 4527 -33
rect 4561 -67 4595 -33
rect 4629 -67 4663 -33
rect 4697 -67 4731 -33
rect 4765 -67 4799 -33
rect 4833 -67 4867 -33
rect 4901 -67 4935 -33
rect 4969 -67 5003 -33
rect 5037 -67 5071 -33
rect 5105 -67 5139 -33
rect 5173 -67 5207 -33
rect 5241 -67 5275 -33
rect 5309 -67 5343 -33
rect 5377 -67 5523 -33
rect 5557 -67 5591 -33
rect 5625 -67 5659 -33
rect 5693 -67 5727 -33
rect 5761 -67 5795 -33
rect 5829 -67 5863 -33
rect 5897 -67 5931 -33
rect 5965 -67 5999 -33
rect 6033 -67 6067 -33
rect 6101 -67 6135 -33
rect 6169 -67 6203 -33
rect 6237 -67 6271 -33
rect 6305 -67 6339 -33
rect 6373 -67 6407 -33
rect 6441 -67 6475 -33
rect 6509 -67 6543 -33
rect 6577 -38 6833 -33
rect 6867 -38 6900 -4
rect 6577 -67 6900 -38
rect 4300 -72 6900 -67
rect 4300 -100 6833 -72
rect 1367 -101 1720 -100
rect 1300 -102 1720 -101
rect 1300 -135 1400 -102
rect 1300 -169 1333 -135
rect 1367 -169 1400 -135
rect 1300 -200 1400 -169
rect 6800 -106 6833 -100
rect 6867 -106 6900 -72
rect 6800 -140 6900 -106
rect 6800 -174 6833 -140
rect 6867 -174 6900 -140
rect 6800 -200 6900 -174
rect 1300 -233 6900 -200
rect 1300 -267 1333 -233
rect 1367 -267 1431 -233
rect 1465 -267 1499 -233
rect 1533 -267 1567 -233
rect 1601 -267 1635 -233
rect 1669 -267 1703 -233
rect 1737 -267 1771 -233
rect 1805 -267 1839 -233
rect 1873 -267 1907 -233
rect 1941 -267 1975 -233
rect 2009 -267 2043 -233
rect 2077 -267 2111 -233
rect 2145 -267 2179 -233
rect 2213 -267 2247 -233
rect 2281 -267 2315 -233
rect 2349 -267 2383 -233
rect 2417 -267 2451 -233
rect 2485 -267 2519 -233
rect 2553 -267 2587 -233
rect 2621 -267 2655 -233
rect 2689 -267 2723 -233
rect 2757 -267 2791 -233
rect 2825 -267 2859 -233
rect 2893 -267 2927 -233
rect 2961 -267 2995 -233
rect 3029 -267 3063 -233
rect 3097 -267 3131 -233
rect 3165 -267 3199 -233
rect 3233 -267 3267 -233
rect 3301 -267 3335 -233
rect 3369 -267 3403 -233
rect 3437 -267 3471 -233
rect 3505 -267 3539 -233
rect 3573 -267 3607 -233
rect 3641 -267 3675 -233
rect 3709 -267 3743 -233
rect 3777 -267 3811 -233
rect 3845 -267 3879 -233
rect 3913 -267 3947 -233
rect 3981 -267 4015 -233
rect 4049 -267 4083 -233
rect 4117 -267 4151 -233
rect 4185 -267 4219 -233
rect 4253 -267 4287 -233
rect 4321 -267 4355 -233
rect 4389 -267 4423 -233
rect 4457 -267 4491 -233
rect 4525 -267 4559 -233
rect 4593 -267 4627 -233
rect 4661 -267 4695 -233
rect 4729 -267 4763 -233
rect 4797 -267 4831 -233
rect 4865 -267 4899 -233
rect 4933 -267 4967 -233
rect 5001 -267 5035 -233
rect 5069 -267 5103 -233
rect 5137 -267 5171 -233
rect 5205 -267 5239 -233
rect 5273 -267 5307 -233
rect 5341 -267 5375 -233
rect 5409 -267 5443 -233
rect 5477 -267 5511 -233
rect 5545 -267 5579 -233
rect 5613 -267 5647 -233
rect 5681 -267 5715 -233
rect 5749 -267 5783 -233
rect 5817 -267 5851 -233
rect 5885 -267 5919 -233
rect 5953 -267 5987 -233
rect 6021 -267 6055 -233
rect 6089 -267 6123 -233
rect 6157 -267 6191 -233
rect 6225 -267 6259 -233
rect 6293 -267 6327 -233
rect 6361 -267 6395 -233
rect 6429 -267 6463 -233
rect 6497 -267 6531 -233
rect 6565 -267 6599 -233
rect 6633 -267 6667 -233
rect 6701 -267 6735 -233
rect 6769 -267 6900 -233
rect 1300 -300 6900 -267
<< viali >>
rect 4033 3313 4067 3347
rect 4133 3313 4167 3347
rect 4033 3213 4067 3247
rect 4133 3213 4167 3247
rect 4033 3113 4067 3147
rect 4133 3113 4167 3147
rect 4033 3013 4067 3047
rect 4133 3013 4167 3047
rect 4033 2913 4067 2947
rect 4133 2913 4167 2947
rect 4033 2813 4067 2847
rect 4133 2813 4167 2847
rect 4033 2713 4067 2747
rect 4133 2713 4167 2747
rect 4033 2613 4067 2647
rect 4133 2613 4167 2647
rect 4033 2513 4067 2547
rect 4133 2513 4167 2547
rect 4033 2413 4067 2447
rect 4133 2413 4167 2447
rect 4033 2313 4067 2347
rect 4133 2313 4167 2347
rect 4033 2213 4067 2247
rect 4133 2213 4167 2247
rect 4033 2113 4067 2147
rect 4133 2113 4167 2147
rect 1533 1693 1567 1727
rect 1633 1693 1667 1727
rect 1733 1693 1767 1727
rect 1833 1693 1867 1727
rect 1933 1693 1967 1727
rect 2033 1693 2067 1727
rect 2133 1693 2167 1727
rect 2233 1693 2267 1727
rect 2333 1693 2367 1727
rect 2433 1693 2467 1727
rect 2533 1693 2567 1727
rect 2633 1693 2667 1727
rect 2733 1693 2767 1727
rect 2833 1693 2867 1727
rect 2933 1693 2967 1727
rect 3033 1693 3067 1727
rect 3133 1693 3167 1727
rect 3233 1693 3267 1727
rect 3333 1693 3367 1727
rect 3433 1693 3467 1727
rect 3533 1693 3567 1727
rect 3633 1693 3667 1727
rect 3733 1693 3767 1727
rect 3833 1693 3867 1727
rect 3933 1693 3967 1727
rect 4033 1693 4067 1727
rect 4133 1693 4167 1727
rect 4233 1693 4267 1727
rect 4333 1693 4367 1727
rect 4433 1693 4467 1727
rect 4533 1693 4567 1727
rect 4633 1693 4667 1727
rect 4733 1693 4767 1727
rect 4833 1693 4867 1727
rect 4933 1693 4967 1727
rect 5033 1693 5067 1727
rect 5133 1693 5167 1727
rect 5233 1693 5267 1727
rect 5333 1693 5367 1727
rect 5433 1693 5467 1727
rect 5533 1693 5567 1727
rect 5633 1693 5667 1727
rect 5733 1693 5767 1727
rect 5833 1693 5867 1727
rect 5933 1693 5967 1727
rect 6033 1693 6067 1727
rect 6133 1693 6167 1727
rect 6233 1693 6267 1727
rect 6333 1693 6367 1727
rect 6433 1693 6467 1727
rect 6533 1693 6567 1727
rect 6633 1693 6667 1727
rect 1533 1573 1567 1607
rect 1633 1573 1667 1607
rect 1733 1573 1767 1607
rect 1833 1573 1867 1607
rect 1933 1573 1967 1607
rect 2033 1573 2067 1607
rect 2133 1573 2167 1607
rect 2233 1573 2267 1607
rect 2333 1573 2367 1607
rect 2433 1573 2467 1607
rect 2533 1573 2567 1607
rect 2633 1573 2667 1607
rect 2733 1573 2767 1607
rect 2833 1573 2867 1607
rect 2933 1573 2967 1607
rect 3033 1573 3067 1607
rect 3133 1573 3167 1607
rect 3233 1573 3267 1607
rect 3333 1573 3367 1607
rect 3433 1573 3467 1607
rect 3533 1573 3567 1607
rect 3633 1573 3667 1607
rect 3733 1573 3767 1607
rect 3833 1573 3867 1607
rect 3933 1573 3967 1607
rect 4033 1573 4067 1607
rect 4133 1573 4167 1607
rect 4233 1573 4267 1607
rect 4333 1573 4367 1607
rect 4433 1573 4467 1607
rect 4533 1573 4567 1607
rect 4633 1573 4667 1607
rect 4733 1573 4767 1607
rect 4833 1573 4867 1607
rect 4933 1573 4967 1607
rect 5033 1573 5067 1607
rect 5133 1573 5167 1607
rect 5233 1573 5267 1607
rect 5333 1573 5367 1607
rect 5433 1573 5467 1607
rect 5533 1573 5567 1607
rect 5633 1573 5667 1607
rect 5733 1573 5767 1607
rect 5833 1573 5867 1607
rect 5933 1573 5967 1607
rect 6033 1573 6067 1607
rect 6133 1573 6167 1607
rect 6233 1573 6267 1607
rect 6333 1573 6367 1607
rect 6433 1573 6467 1607
rect 6533 1573 6567 1607
rect 6633 1573 6667 1607
rect 4033 1153 4067 1187
rect 4133 1153 4167 1187
rect 4033 1053 4067 1087
rect 4133 1053 4167 1087
rect 4033 953 4067 987
rect 4133 953 4167 987
rect 4033 853 4067 887
rect 4133 853 4167 887
rect 4033 753 4067 787
rect 4133 753 4167 787
rect 4033 653 4067 687
rect 4133 653 4167 687
rect 4033 553 4067 587
rect 4133 553 4167 587
rect 4033 453 4067 487
rect 4133 453 4167 487
rect 4033 353 4067 387
rect 4133 353 4167 387
rect 4033 253 4067 287
rect 4133 253 4167 287
rect 4033 153 4067 187
rect 4133 153 4167 187
rect 4033 53 4067 87
rect 4133 53 4167 87
rect 4033 -47 4067 -13
rect 4133 -47 4167 -13
rect 1333 -267 1367 -233
<< metal1 >>
rect 2020 3356 2280 3380
rect 2020 3304 2044 3356
rect 2096 3304 2204 3356
rect 2256 3304 2280 3356
rect 2020 3256 2280 3304
rect 2020 3204 2044 3256
rect 2096 3204 2204 3256
rect 2256 3204 2280 3256
rect 1800 2876 1980 3140
rect 2020 3060 2280 3204
rect 4000 3376 4200 3400
rect 4000 3324 4024 3376
rect 4076 3324 4124 3376
rect 4176 3324 4200 3376
rect 4000 3313 4033 3324
rect 4067 3313 4133 3324
rect 4167 3313 4200 3324
rect 4000 3296 4200 3313
rect 4000 3244 4024 3296
rect 4076 3244 4124 3296
rect 4176 3244 4200 3296
rect 4000 3216 4033 3244
rect 4067 3216 4133 3244
rect 4167 3216 4200 3244
rect 4000 3164 4024 3216
rect 4076 3164 4124 3216
rect 4176 3164 4200 3216
rect 4000 3147 4200 3164
rect 5920 3356 6180 3380
rect 5920 3304 5944 3356
rect 5996 3304 6104 3356
rect 6156 3304 6180 3356
rect 5920 3256 6180 3304
rect 5920 3204 5944 3256
rect 5996 3204 6104 3256
rect 6156 3204 6180 3256
rect 1800 2824 1824 2876
rect 1876 2824 1980 2876
rect 1800 2776 1980 2824
rect 1800 2724 1824 2776
rect 1876 2724 1980 2776
rect 1800 2100 1980 2724
rect 2320 2876 2500 3140
rect 3000 2900 3180 3140
rect 2320 2824 2424 2876
rect 2476 2824 2500 2876
rect 2320 2776 2500 2824
rect 2320 2724 2424 2776
rect 2476 2724 2500 2776
rect 2320 2100 2500 2724
rect 2980 2700 3180 2900
rect 3000 2500 3180 2700
rect 2980 2476 3180 2500
rect 2980 2424 3004 2476
rect 3056 2424 3180 2476
rect 2980 2376 3180 2424
rect 2980 2324 3004 2376
rect 3056 2324 3180 2376
rect 2980 2300 3180 2324
rect 3000 2100 3180 2300
rect 3520 2476 3700 3140
rect 3520 2424 3624 2476
rect 3676 2424 3700 2476
rect 3520 2376 3700 2424
rect 3520 2324 3624 2376
rect 3676 2324 3700 2376
rect 3240 2140 3460 2160
rect 3220 2000 3480 2140
rect 3520 2100 3700 2324
rect 4000 3136 4033 3147
rect 4067 3136 4133 3147
rect 4167 3136 4200 3147
rect 4000 3084 4024 3136
rect 4076 3084 4124 3136
rect 4176 3084 4200 3136
rect 4000 3056 4200 3084
rect 4000 3004 4024 3056
rect 4076 3004 4124 3056
rect 4176 3004 4200 3056
rect 4000 2976 4200 3004
rect 4000 2924 4024 2976
rect 4076 2924 4124 2976
rect 4176 2924 4200 2976
rect 4000 2913 4033 2924
rect 4067 2913 4133 2924
rect 4167 2913 4200 2924
rect 4000 2896 4200 2913
rect 4000 2844 4024 2896
rect 4076 2844 4124 2896
rect 4176 2844 4200 2896
rect 4000 2816 4033 2844
rect 4067 2816 4133 2844
rect 4167 2816 4200 2844
rect 4000 2764 4024 2816
rect 4076 2764 4124 2816
rect 4176 2764 4200 2816
rect 4000 2747 4200 2764
rect 4000 2736 4033 2747
rect 4067 2736 4133 2747
rect 4167 2736 4200 2747
rect 4000 2684 4024 2736
rect 4076 2684 4124 2736
rect 4176 2684 4200 2736
rect 4000 2656 4200 2684
rect 4000 2604 4024 2656
rect 4076 2604 4124 2656
rect 4176 2604 4200 2656
rect 4000 2576 4200 2604
rect 4000 2524 4024 2576
rect 4076 2524 4124 2576
rect 4176 2524 4200 2576
rect 4000 2513 4033 2524
rect 4067 2513 4133 2524
rect 4167 2513 4200 2524
rect 4000 2496 4200 2513
rect 4500 2500 4680 3140
rect 4000 2444 4024 2496
rect 4076 2444 4124 2496
rect 4176 2444 4200 2496
rect 4000 2416 4033 2444
rect 4067 2416 4133 2444
rect 4167 2416 4200 2444
rect 4000 2364 4024 2416
rect 4076 2364 4124 2416
rect 4176 2364 4200 2416
rect 4000 2347 4200 2364
rect 4000 2336 4033 2347
rect 4067 2336 4133 2347
rect 4167 2336 4200 2347
rect 4000 2284 4024 2336
rect 4076 2284 4124 2336
rect 4176 2284 4200 2336
rect 4480 2476 4680 2500
rect 4480 2424 4504 2476
rect 4556 2424 4680 2476
rect 4480 2376 4680 2424
rect 4480 2324 4504 2376
rect 4556 2324 4680 2376
rect 4480 2300 4680 2324
rect 4000 2256 4200 2284
rect 4000 2204 4024 2256
rect 4076 2204 4124 2256
rect 4176 2204 4200 2256
rect 4000 2176 4200 2204
rect 4000 2124 4024 2176
rect 4076 2124 4124 2176
rect 4176 2124 4200 2176
rect 4000 2113 4033 2124
rect 4067 2113 4133 2124
rect 4167 2113 4200 2124
rect 4000 2080 4200 2113
rect 4500 2100 4680 2300
rect 5020 2500 5180 3140
rect 5700 2900 5880 3160
rect 5920 3060 6180 3204
rect 5680 2876 5880 2900
rect 5680 2824 5704 2876
rect 5756 2824 5880 2876
rect 5680 2776 5880 2824
rect 5680 2724 5704 2776
rect 5756 2724 5880 2776
rect 5680 2700 5880 2724
rect 5020 2476 5200 2500
rect 5020 2424 5124 2476
rect 5176 2424 5200 2476
rect 5020 2376 5200 2424
rect 5020 2324 5124 2376
rect 5176 2324 5200 2376
rect 5020 2300 5200 2324
rect 4720 2000 4980 2160
rect 5020 2100 5180 2300
rect 5700 2100 5880 2700
rect 6220 2876 6400 3160
rect 6220 2824 6324 2876
rect 6376 2824 6400 2876
rect 6220 2776 6400 2824
rect 6220 2724 6324 2776
rect 6376 2724 6400 2776
rect 6220 2100 6400 2724
rect 900 1976 7300 2000
rect 900 1924 1524 1976
rect 1576 1924 1624 1976
rect 1676 1924 6524 1976
rect 6576 1924 6624 1976
rect 6676 1924 7300 1976
rect 900 1876 7300 1924
rect 900 1824 1524 1876
rect 1576 1824 1624 1876
rect 1676 1824 6524 1876
rect 6576 1824 6624 1876
rect 6676 1824 7300 1876
rect 900 1800 7300 1824
rect 1500 1736 6700 1760
rect 1500 1727 4024 1736
rect 1500 1693 1533 1727
rect 1567 1693 1633 1727
rect 1667 1693 1733 1727
rect 1767 1693 1833 1727
rect 1867 1693 1933 1727
rect 1967 1693 2033 1727
rect 2067 1693 2133 1727
rect 2167 1693 2233 1727
rect 2267 1693 2333 1727
rect 2367 1693 2433 1727
rect 2467 1693 2533 1727
rect 2567 1693 2633 1727
rect 2667 1693 2733 1727
rect 2767 1693 2833 1727
rect 2867 1693 2933 1727
rect 2967 1693 3033 1727
rect 3067 1693 3133 1727
rect 3167 1693 3233 1727
rect 3267 1693 3333 1727
rect 3367 1693 3433 1727
rect 3467 1693 3533 1727
rect 3567 1693 3633 1727
rect 3667 1693 3733 1727
rect 3767 1693 3833 1727
rect 3867 1693 3933 1727
rect 3967 1693 4024 1727
rect 1500 1684 4024 1693
rect 4076 1684 4124 1736
rect 4176 1727 6700 1736
rect 4176 1693 4233 1727
rect 4267 1693 4333 1727
rect 4367 1693 4433 1727
rect 4467 1693 4533 1727
rect 4567 1693 4633 1727
rect 4667 1693 4733 1727
rect 4767 1693 4833 1727
rect 4867 1693 4933 1727
rect 4967 1693 5033 1727
rect 5067 1693 5133 1727
rect 5167 1693 5233 1727
rect 5267 1693 5333 1727
rect 5367 1693 5433 1727
rect 5467 1693 5533 1727
rect 5567 1693 5633 1727
rect 5667 1693 5733 1727
rect 5767 1693 5833 1727
rect 5867 1693 5933 1727
rect 5967 1693 6033 1727
rect 6067 1693 6133 1727
rect 6167 1693 6233 1727
rect 6267 1693 6333 1727
rect 6367 1693 6433 1727
rect 6467 1693 6533 1727
rect 6567 1693 6633 1727
rect 6667 1693 6700 1727
rect 4176 1684 6700 1693
rect 1500 1616 6700 1684
rect 1500 1607 4024 1616
rect 1500 1573 1533 1607
rect 1567 1573 1633 1607
rect 1667 1573 1733 1607
rect 1767 1573 1833 1607
rect 1867 1573 1933 1607
rect 1967 1573 2033 1607
rect 2067 1573 2133 1607
rect 2167 1573 2233 1607
rect 2267 1573 2333 1607
rect 2367 1573 2433 1607
rect 2467 1573 2533 1607
rect 2567 1573 2633 1607
rect 2667 1573 2733 1607
rect 2767 1573 2833 1607
rect 2867 1573 2933 1607
rect 2967 1573 3033 1607
rect 3067 1573 3133 1607
rect 3167 1573 3233 1607
rect 3267 1573 3333 1607
rect 3367 1573 3433 1607
rect 3467 1573 3533 1607
rect 3567 1573 3633 1607
rect 3667 1573 3733 1607
rect 3767 1573 3833 1607
rect 3867 1573 3933 1607
rect 3967 1573 4024 1607
rect 1500 1564 4024 1573
rect 4076 1564 4124 1616
rect 4176 1607 6700 1616
rect 4176 1573 4233 1607
rect 4267 1573 4333 1607
rect 4367 1573 4433 1607
rect 4467 1573 4533 1607
rect 4567 1573 4633 1607
rect 4667 1573 4733 1607
rect 4767 1573 4833 1607
rect 4867 1573 4933 1607
rect 4967 1573 5033 1607
rect 5067 1573 5133 1607
rect 5167 1573 5233 1607
rect 5267 1573 5333 1607
rect 5367 1573 5433 1607
rect 5467 1573 5533 1607
rect 5567 1573 5633 1607
rect 5667 1573 5733 1607
rect 5767 1573 5833 1607
rect 5867 1573 5933 1607
rect 5967 1573 6033 1607
rect 6067 1573 6133 1607
rect 6167 1573 6233 1607
rect 6267 1573 6333 1607
rect 6367 1573 6433 1607
rect 6467 1573 6533 1607
rect 6567 1573 6633 1607
rect 6667 1573 6700 1607
rect 4176 1564 6700 1573
rect 1500 1540 6700 1564
rect 900 1476 7300 1500
rect 900 1424 2624 1476
rect 2676 1424 2724 1476
rect 2776 1424 5424 1476
rect 5476 1424 5524 1476
rect 5576 1424 7300 1476
rect 900 1376 7300 1424
rect 900 1324 2624 1376
rect 2676 1324 2724 1376
rect 2776 1324 5424 1376
rect 5476 1324 5524 1376
rect 5576 1324 7300 1376
rect 900 1300 7300 1324
rect 1800 976 1980 1260
rect 1800 924 1824 976
rect 1876 924 1980 976
rect 1800 876 1980 924
rect 1800 824 1824 876
rect 1876 824 1980 876
rect 1800 200 1980 824
rect 2320 976 2500 1260
rect 2320 924 2404 976
rect 2456 924 2500 976
rect 2320 876 2500 924
rect 2320 824 2404 876
rect 2456 824 2500 876
rect 2020 96 2280 240
rect 2320 200 2500 824
rect 3000 576 3180 1260
rect 3220 1160 3480 1300
rect 3000 524 3024 576
rect 3076 524 3180 576
rect 3000 476 3180 524
rect 3000 424 3024 476
rect 3076 424 3180 476
rect 3000 200 3180 424
rect 3520 576 3700 1260
rect 3520 524 3604 576
rect 3656 524 3700 576
rect 3520 476 3700 524
rect 3520 424 3604 476
rect 3656 424 3700 476
rect 3520 200 3700 424
rect 4000 1187 4200 1220
rect 4000 1176 4033 1187
rect 4067 1176 4133 1187
rect 4167 1176 4200 1187
rect 4000 1124 4024 1176
rect 4076 1124 4124 1176
rect 4176 1124 4200 1176
rect 4000 1096 4200 1124
rect 4000 1044 4024 1096
rect 4076 1044 4124 1096
rect 4176 1044 4200 1096
rect 4000 1016 4200 1044
rect 4000 964 4024 1016
rect 4076 964 4124 1016
rect 4176 964 4200 1016
rect 4000 953 4033 964
rect 4067 953 4133 964
rect 4167 953 4200 964
rect 4000 936 4200 953
rect 4000 884 4024 936
rect 4076 884 4124 936
rect 4176 884 4200 936
rect 4000 856 4033 884
rect 4067 856 4133 884
rect 4167 856 4200 884
rect 4000 804 4024 856
rect 4076 804 4124 856
rect 4176 804 4200 856
rect 4000 787 4200 804
rect 4000 776 4033 787
rect 4067 776 4133 787
rect 4167 776 4200 787
rect 4000 724 4024 776
rect 4076 724 4124 776
rect 4176 724 4200 776
rect 4000 696 4200 724
rect 4000 644 4024 696
rect 4076 644 4124 696
rect 4176 644 4200 696
rect 4000 616 4200 644
rect 4000 564 4024 616
rect 4076 564 4124 616
rect 4176 564 4200 616
rect 4000 553 4033 564
rect 4067 553 4133 564
rect 4167 553 4200 564
rect 4000 536 4200 553
rect 4000 484 4024 536
rect 4076 484 4124 536
rect 4176 484 4200 536
rect 4000 456 4033 484
rect 4067 456 4133 484
rect 4167 456 4200 484
rect 4000 404 4024 456
rect 4076 404 4124 456
rect 4176 404 4200 456
rect 4000 387 4200 404
rect 4000 376 4033 387
rect 4067 376 4133 387
rect 4167 376 4200 387
rect 4000 324 4024 376
rect 4076 324 4124 376
rect 4176 324 4200 376
rect 4000 296 4200 324
rect 4000 244 4024 296
rect 4076 244 4124 296
rect 4176 244 4200 296
rect 4000 216 4200 244
rect 2020 44 2044 96
rect 2096 44 2204 96
rect 2256 44 2280 96
rect 2020 -4 2280 44
rect 2020 -56 2044 -4
rect 2096 -56 2204 -4
rect 2256 -56 2280 -4
rect 2020 -80 2280 -56
rect 4000 164 4024 216
rect 4076 164 4124 216
rect 4176 164 4200 216
rect 4500 576 4680 1260
rect 4720 1160 4980 1300
rect 4500 524 4524 576
rect 4576 524 4680 576
rect 4500 476 4680 524
rect 4500 424 4524 476
rect 4576 424 4680 476
rect 4500 200 4680 424
rect 5020 576 5200 1260
rect 5020 524 5104 576
rect 5156 524 5200 576
rect 5020 476 5200 524
rect 5020 424 5104 476
rect 5156 424 5200 476
rect 5020 200 5200 424
rect 5700 976 5880 1260
rect 5700 924 5724 976
rect 5776 924 5880 976
rect 5700 876 5880 924
rect 5700 824 5724 876
rect 5776 824 5880 876
rect 5700 200 5880 824
rect 6220 976 6400 1260
rect 6220 924 6304 976
rect 6356 924 6400 976
rect 6220 876 6400 924
rect 6220 824 6304 876
rect 6356 824 6400 876
rect 4000 153 4033 164
rect 4067 153 4133 164
rect 4167 153 4200 164
rect 4000 136 4200 153
rect 4000 84 4024 136
rect 4076 84 4124 136
rect 4176 84 4200 136
rect 4000 56 4033 84
rect 4067 56 4133 84
rect 4167 56 4200 84
rect 4000 4 4024 56
rect 4076 4 4124 56
rect 4176 4 4200 56
rect 4000 -13 4200 4
rect 4000 -24 4033 -13
rect 4067 -24 4133 -13
rect 4167 -24 4200 -13
rect 4000 -76 4024 -24
rect 4076 -76 4124 -24
rect 4176 -76 4200 -24
rect 4000 -100 4200 -76
rect 5920 96 6180 260
rect 6220 200 6400 824
rect 5920 44 5944 96
rect 5996 44 6104 96
rect 6156 44 6180 96
rect 5920 -4 6180 44
rect 5920 -56 5944 -4
rect 5996 -56 6104 -4
rect 6156 -56 6180 -4
rect 5920 -80 6180 -56
rect 300 -124 500 -100
rect 300 -176 324 -124
rect 376 -176 424 -124
rect 476 -176 500 -124
rect 300 -224 500 -176
rect 300 -276 324 -224
rect 376 -276 424 -224
rect 476 -276 500 -224
rect 300 -300 500 -276
rect 600 -124 800 -100
rect 600 -176 624 -124
rect 676 -176 724 -124
rect 776 -176 800 -124
rect 600 -224 800 -176
rect 7400 -124 7600 -100
rect 7400 -176 7424 -124
rect 7476 -176 7524 -124
rect 7576 -176 7600 -124
rect 600 -276 624 -224
rect 676 -276 724 -224
rect 776 -276 800 -224
rect 600 -300 800 -276
rect 1300 -233 1400 -200
rect 1300 -267 1333 -233
rect 1367 -267 1400 -233
rect 1300 -300 1400 -267
rect 7400 -224 7600 -176
rect 7400 -276 7424 -224
rect 7476 -276 7524 -224
rect 7576 -276 7600 -224
rect 7400 -300 7600 -276
rect 7700 -124 7900 -100
rect 7700 -176 7724 -124
rect 7776 -176 7824 -124
rect 7876 -176 7900 -124
rect 7700 -224 7900 -176
rect 7700 -276 7724 -224
rect 7776 -276 7824 -224
rect 7876 -276 7900 -224
rect 7700 -300 7900 -276
rect 4000 -324 4200 -300
rect 4000 -376 4024 -324
rect 4076 -376 4124 -324
rect 4176 -376 4200 -324
rect 4000 -424 4200 -376
rect 4000 -476 4024 -424
rect 4076 -476 4124 -424
rect 4176 -476 4200 -424
rect 4000 -500 4200 -476
<< via1 >>
rect 2044 3304 2096 3356
rect 2204 3304 2256 3356
rect 2044 3204 2096 3256
rect 2204 3204 2256 3256
rect 4024 3347 4076 3376
rect 4024 3324 4033 3347
rect 4033 3324 4067 3347
rect 4067 3324 4076 3347
rect 4124 3347 4176 3376
rect 4124 3324 4133 3347
rect 4133 3324 4167 3347
rect 4167 3324 4176 3347
rect 4024 3247 4076 3296
rect 4024 3244 4033 3247
rect 4033 3244 4067 3247
rect 4067 3244 4076 3247
rect 4124 3247 4176 3296
rect 4124 3244 4133 3247
rect 4133 3244 4167 3247
rect 4167 3244 4176 3247
rect 4024 3213 4033 3216
rect 4033 3213 4067 3216
rect 4067 3213 4076 3216
rect 4024 3164 4076 3213
rect 4124 3213 4133 3216
rect 4133 3213 4167 3216
rect 4167 3213 4176 3216
rect 4124 3164 4176 3213
rect 5944 3304 5996 3356
rect 6104 3304 6156 3356
rect 5944 3204 5996 3256
rect 6104 3204 6156 3256
rect 1824 2824 1876 2876
rect 1824 2724 1876 2776
rect 2424 2824 2476 2876
rect 2424 2724 2476 2776
rect 3004 2424 3056 2476
rect 3004 2324 3056 2376
rect 3624 2424 3676 2476
rect 3624 2324 3676 2376
rect 4024 3113 4033 3136
rect 4033 3113 4067 3136
rect 4067 3113 4076 3136
rect 4024 3084 4076 3113
rect 4124 3113 4133 3136
rect 4133 3113 4167 3136
rect 4167 3113 4176 3136
rect 4124 3084 4176 3113
rect 4024 3047 4076 3056
rect 4024 3013 4033 3047
rect 4033 3013 4067 3047
rect 4067 3013 4076 3047
rect 4024 3004 4076 3013
rect 4124 3047 4176 3056
rect 4124 3013 4133 3047
rect 4133 3013 4167 3047
rect 4167 3013 4176 3047
rect 4124 3004 4176 3013
rect 4024 2947 4076 2976
rect 4024 2924 4033 2947
rect 4033 2924 4067 2947
rect 4067 2924 4076 2947
rect 4124 2947 4176 2976
rect 4124 2924 4133 2947
rect 4133 2924 4167 2947
rect 4167 2924 4176 2947
rect 4024 2847 4076 2896
rect 4024 2844 4033 2847
rect 4033 2844 4067 2847
rect 4067 2844 4076 2847
rect 4124 2847 4176 2896
rect 4124 2844 4133 2847
rect 4133 2844 4167 2847
rect 4167 2844 4176 2847
rect 4024 2813 4033 2816
rect 4033 2813 4067 2816
rect 4067 2813 4076 2816
rect 4024 2764 4076 2813
rect 4124 2813 4133 2816
rect 4133 2813 4167 2816
rect 4167 2813 4176 2816
rect 4124 2764 4176 2813
rect 4024 2713 4033 2736
rect 4033 2713 4067 2736
rect 4067 2713 4076 2736
rect 4024 2684 4076 2713
rect 4124 2713 4133 2736
rect 4133 2713 4167 2736
rect 4167 2713 4176 2736
rect 4124 2684 4176 2713
rect 4024 2647 4076 2656
rect 4024 2613 4033 2647
rect 4033 2613 4067 2647
rect 4067 2613 4076 2647
rect 4024 2604 4076 2613
rect 4124 2647 4176 2656
rect 4124 2613 4133 2647
rect 4133 2613 4167 2647
rect 4167 2613 4176 2647
rect 4124 2604 4176 2613
rect 4024 2547 4076 2576
rect 4024 2524 4033 2547
rect 4033 2524 4067 2547
rect 4067 2524 4076 2547
rect 4124 2547 4176 2576
rect 4124 2524 4133 2547
rect 4133 2524 4167 2547
rect 4167 2524 4176 2547
rect 4024 2447 4076 2496
rect 4024 2444 4033 2447
rect 4033 2444 4067 2447
rect 4067 2444 4076 2447
rect 4124 2447 4176 2496
rect 4124 2444 4133 2447
rect 4133 2444 4167 2447
rect 4167 2444 4176 2447
rect 4024 2413 4033 2416
rect 4033 2413 4067 2416
rect 4067 2413 4076 2416
rect 4024 2364 4076 2413
rect 4124 2413 4133 2416
rect 4133 2413 4167 2416
rect 4167 2413 4176 2416
rect 4124 2364 4176 2413
rect 4024 2313 4033 2336
rect 4033 2313 4067 2336
rect 4067 2313 4076 2336
rect 4024 2284 4076 2313
rect 4124 2313 4133 2336
rect 4133 2313 4167 2336
rect 4167 2313 4176 2336
rect 4124 2284 4176 2313
rect 4504 2424 4556 2476
rect 4504 2324 4556 2376
rect 4024 2247 4076 2256
rect 4024 2213 4033 2247
rect 4033 2213 4067 2247
rect 4067 2213 4076 2247
rect 4024 2204 4076 2213
rect 4124 2247 4176 2256
rect 4124 2213 4133 2247
rect 4133 2213 4167 2247
rect 4167 2213 4176 2247
rect 4124 2204 4176 2213
rect 4024 2147 4076 2176
rect 4024 2124 4033 2147
rect 4033 2124 4067 2147
rect 4067 2124 4076 2147
rect 4124 2147 4176 2176
rect 4124 2124 4133 2147
rect 4133 2124 4167 2147
rect 4167 2124 4176 2147
rect 5704 2824 5756 2876
rect 5704 2724 5756 2776
rect 5124 2424 5176 2476
rect 5124 2324 5176 2376
rect 6324 2824 6376 2876
rect 6324 2724 6376 2776
rect 1524 1924 1576 1976
rect 1624 1924 1676 1976
rect 6524 1924 6576 1976
rect 6624 1924 6676 1976
rect 1524 1824 1576 1876
rect 1624 1824 1676 1876
rect 6524 1824 6576 1876
rect 6624 1824 6676 1876
rect 4024 1727 4076 1736
rect 4024 1693 4033 1727
rect 4033 1693 4067 1727
rect 4067 1693 4076 1727
rect 4024 1684 4076 1693
rect 4124 1727 4176 1736
rect 4124 1693 4133 1727
rect 4133 1693 4167 1727
rect 4167 1693 4176 1727
rect 4124 1684 4176 1693
rect 4024 1607 4076 1616
rect 4024 1573 4033 1607
rect 4033 1573 4067 1607
rect 4067 1573 4076 1607
rect 4024 1564 4076 1573
rect 4124 1607 4176 1616
rect 4124 1573 4133 1607
rect 4133 1573 4167 1607
rect 4167 1573 4176 1607
rect 4124 1564 4176 1573
rect 2624 1424 2676 1476
rect 2724 1424 2776 1476
rect 5424 1424 5476 1476
rect 5524 1424 5576 1476
rect 2624 1324 2676 1376
rect 2724 1324 2776 1376
rect 5424 1324 5476 1376
rect 5524 1324 5576 1376
rect 1824 924 1876 976
rect 1824 824 1876 876
rect 2404 924 2456 976
rect 2404 824 2456 876
rect 3024 524 3076 576
rect 3024 424 3076 476
rect 3604 524 3656 576
rect 3604 424 3656 476
rect 4024 1153 4033 1176
rect 4033 1153 4067 1176
rect 4067 1153 4076 1176
rect 4024 1124 4076 1153
rect 4124 1153 4133 1176
rect 4133 1153 4167 1176
rect 4167 1153 4176 1176
rect 4124 1124 4176 1153
rect 4024 1087 4076 1096
rect 4024 1053 4033 1087
rect 4033 1053 4067 1087
rect 4067 1053 4076 1087
rect 4024 1044 4076 1053
rect 4124 1087 4176 1096
rect 4124 1053 4133 1087
rect 4133 1053 4167 1087
rect 4167 1053 4176 1087
rect 4124 1044 4176 1053
rect 4024 987 4076 1016
rect 4024 964 4033 987
rect 4033 964 4067 987
rect 4067 964 4076 987
rect 4124 987 4176 1016
rect 4124 964 4133 987
rect 4133 964 4167 987
rect 4167 964 4176 987
rect 4024 887 4076 936
rect 4024 884 4033 887
rect 4033 884 4067 887
rect 4067 884 4076 887
rect 4124 887 4176 936
rect 4124 884 4133 887
rect 4133 884 4167 887
rect 4167 884 4176 887
rect 4024 853 4033 856
rect 4033 853 4067 856
rect 4067 853 4076 856
rect 4024 804 4076 853
rect 4124 853 4133 856
rect 4133 853 4167 856
rect 4167 853 4176 856
rect 4124 804 4176 853
rect 4024 753 4033 776
rect 4033 753 4067 776
rect 4067 753 4076 776
rect 4024 724 4076 753
rect 4124 753 4133 776
rect 4133 753 4167 776
rect 4167 753 4176 776
rect 4124 724 4176 753
rect 4024 687 4076 696
rect 4024 653 4033 687
rect 4033 653 4067 687
rect 4067 653 4076 687
rect 4024 644 4076 653
rect 4124 687 4176 696
rect 4124 653 4133 687
rect 4133 653 4167 687
rect 4167 653 4176 687
rect 4124 644 4176 653
rect 4024 587 4076 616
rect 4024 564 4033 587
rect 4033 564 4067 587
rect 4067 564 4076 587
rect 4124 587 4176 616
rect 4124 564 4133 587
rect 4133 564 4167 587
rect 4167 564 4176 587
rect 4024 487 4076 536
rect 4024 484 4033 487
rect 4033 484 4067 487
rect 4067 484 4076 487
rect 4124 487 4176 536
rect 4124 484 4133 487
rect 4133 484 4167 487
rect 4167 484 4176 487
rect 4024 453 4033 456
rect 4033 453 4067 456
rect 4067 453 4076 456
rect 4024 404 4076 453
rect 4124 453 4133 456
rect 4133 453 4167 456
rect 4167 453 4176 456
rect 4124 404 4176 453
rect 4024 353 4033 376
rect 4033 353 4067 376
rect 4067 353 4076 376
rect 4024 324 4076 353
rect 4124 353 4133 376
rect 4133 353 4167 376
rect 4167 353 4176 376
rect 4124 324 4176 353
rect 4024 287 4076 296
rect 4024 253 4033 287
rect 4033 253 4067 287
rect 4067 253 4076 287
rect 4024 244 4076 253
rect 4124 287 4176 296
rect 4124 253 4133 287
rect 4133 253 4167 287
rect 4167 253 4176 287
rect 4124 244 4176 253
rect 2044 44 2096 96
rect 2204 44 2256 96
rect 2044 -56 2096 -4
rect 2204 -56 2256 -4
rect 4024 187 4076 216
rect 4024 164 4033 187
rect 4033 164 4067 187
rect 4067 164 4076 187
rect 4124 187 4176 216
rect 4124 164 4133 187
rect 4133 164 4167 187
rect 4167 164 4176 187
rect 4524 524 4576 576
rect 4524 424 4576 476
rect 5104 524 5156 576
rect 5104 424 5156 476
rect 5724 924 5776 976
rect 5724 824 5776 876
rect 6304 924 6356 976
rect 6304 824 6356 876
rect 4024 87 4076 136
rect 4024 84 4033 87
rect 4033 84 4067 87
rect 4067 84 4076 87
rect 4124 87 4176 136
rect 4124 84 4133 87
rect 4133 84 4167 87
rect 4167 84 4176 87
rect 4024 53 4033 56
rect 4033 53 4067 56
rect 4067 53 4076 56
rect 4024 4 4076 53
rect 4124 53 4133 56
rect 4133 53 4167 56
rect 4167 53 4176 56
rect 4124 4 4176 53
rect 4024 -47 4033 -24
rect 4033 -47 4067 -24
rect 4067 -47 4076 -24
rect 4024 -76 4076 -47
rect 4124 -47 4133 -24
rect 4133 -47 4167 -24
rect 4167 -47 4176 -24
rect 4124 -76 4176 -47
rect 5944 44 5996 96
rect 6104 44 6156 96
rect 5944 -56 5996 -4
rect 6104 -56 6156 -4
rect 324 -176 376 -124
rect 424 -176 476 -124
rect 324 -276 376 -224
rect 424 -276 476 -224
rect 624 -176 676 -124
rect 724 -176 776 -124
rect 7424 -176 7476 -124
rect 7524 -176 7576 -124
rect 624 -276 676 -224
rect 724 -276 776 -224
rect 7424 -276 7476 -224
rect 7524 -276 7576 -224
rect 7724 -176 7776 -124
rect 7824 -176 7876 -124
rect 7724 -276 7776 -224
rect 7824 -276 7876 -224
rect 4024 -376 4076 -324
rect 4124 -376 4176 -324
rect 4024 -476 4076 -424
rect 4124 -476 4176 -424
<< metal2 >>
rect 300 2478 500 3600
rect 300 2422 322 2478
rect 378 2422 422 2478
rect 478 2422 500 2478
rect 300 2378 500 2422
rect 300 2322 322 2378
rect 378 2322 422 2378
rect 478 2322 500 2378
rect 300 978 500 2322
rect 300 922 322 978
rect 378 922 422 978
rect 478 922 500 978
rect 300 878 500 922
rect 300 822 322 878
rect 378 822 422 878
rect 478 822 500 878
rect 300 -124 500 822
rect 300 -176 324 -124
rect 376 -176 424 -124
rect 476 -176 500 -124
rect 300 -224 500 -176
rect 300 -276 324 -224
rect 376 -276 424 -224
rect 476 -276 500 -224
rect 300 -300 500 -276
rect 600 2878 800 3600
rect 2000 3356 2800 3380
rect 2000 3304 2044 3356
rect 2096 3304 2204 3356
rect 2256 3304 2800 3356
rect 2000 3256 2800 3304
rect 2000 3204 2044 3256
rect 2096 3204 2204 3256
rect 2256 3204 2800 3256
rect 2000 3180 2800 3204
rect 600 2822 622 2878
rect 678 2822 722 2878
rect 778 2822 800 2878
rect 600 2778 800 2822
rect 600 2722 622 2778
rect 678 2722 722 2778
rect 778 2722 800 2778
rect 600 578 800 2722
rect 1800 2878 1900 2900
rect 1800 2822 1822 2878
rect 1878 2822 1900 2878
rect 1800 2778 1900 2822
rect 1800 2722 1822 2778
rect 1878 2722 1900 2778
rect 1800 2700 1900 2722
rect 2400 2878 2500 2900
rect 2400 2822 2422 2878
rect 2478 2822 2500 2878
rect 2400 2778 2500 2822
rect 2400 2722 2422 2778
rect 2478 2722 2500 2778
rect 2400 2700 2500 2722
rect 600 522 622 578
rect 678 522 722 578
rect 778 522 800 578
rect 600 478 800 522
rect 600 422 622 478
rect 678 422 722 478
rect 778 422 800 478
rect 600 -124 800 422
rect 1500 1976 1700 2000
rect 1500 1924 1524 1976
rect 1576 1924 1624 1976
rect 1676 1924 1700 1976
rect 1500 1876 1700 1924
rect 1500 1824 1524 1876
rect 1576 1824 1624 1876
rect 1676 1824 1700 1876
rect 1500 120 1700 1824
rect 2600 1476 2800 3180
rect 4000 3376 4200 3400
rect 4000 3324 4024 3376
rect 4076 3324 4124 3376
rect 4176 3324 4200 3376
rect 4000 3296 4200 3324
rect 4000 3244 4024 3296
rect 4076 3244 4124 3296
rect 4176 3244 4200 3296
rect 4000 3216 4200 3244
rect 4000 3164 4024 3216
rect 4076 3164 4124 3216
rect 4176 3164 4200 3216
rect 4000 3136 4200 3164
rect 4000 3084 4024 3136
rect 4076 3084 4124 3136
rect 4176 3084 4200 3136
rect 4000 3056 4200 3084
rect 4000 3004 4024 3056
rect 4076 3004 4124 3056
rect 4176 3004 4200 3056
rect 4000 2976 4200 3004
rect 4000 2924 4024 2976
rect 4076 2924 4124 2976
rect 4176 2924 4200 2976
rect 4000 2896 4200 2924
rect 4000 2844 4024 2896
rect 4076 2844 4124 2896
rect 4176 2844 4200 2896
rect 4000 2816 4200 2844
rect 4000 2764 4024 2816
rect 4076 2764 4124 2816
rect 4176 2764 4200 2816
rect 4000 2736 4200 2764
rect 4000 2684 4024 2736
rect 4076 2684 4124 2736
rect 4176 2684 4200 2736
rect 4000 2656 4200 2684
rect 4000 2604 4024 2656
rect 4076 2604 4124 2656
rect 4176 2604 4200 2656
rect 4000 2576 4200 2604
rect 4000 2524 4024 2576
rect 4076 2524 4124 2576
rect 4176 2524 4200 2576
rect 2980 2478 3080 2500
rect 2980 2422 3002 2478
rect 3058 2422 3080 2478
rect 2980 2378 3080 2422
rect 2980 2322 3002 2378
rect 3058 2322 3080 2378
rect 2980 2300 3080 2322
rect 3600 2478 3700 2500
rect 3600 2422 3622 2478
rect 3678 2422 3700 2478
rect 3600 2378 3700 2422
rect 3600 2322 3622 2378
rect 3678 2322 3700 2378
rect 3600 2300 3700 2322
rect 4000 2496 4200 2524
rect 5400 3356 6200 3380
rect 5400 3304 5944 3356
rect 5996 3304 6104 3356
rect 6156 3304 6200 3356
rect 5400 3256 6200 3304
rect 5400 3204 5944 3256
rect 5996 3204 6104 3256
rect 6156 3204 6200 3256
rect 5400 3180 6200 3204
rect 4000 2444 4024 2496
rect 4076 2444 4124 2496
rect 4176 2444 4200 2496
rect 4000 2416 4200 2444
rect 4000 2364 4024 2416
rect 4076 2364 4124 2416
rect 4176 2364 4200 2416
rect 4000 2336 4200 2364
rect 2600 1424 2624 1476
rect 2676 1424 2724 1476
rect 2776 1424 2800 1476
rect 2600 1376 2800 1424
rect 2600 1324 2624 1376
rect 2676 1324 2724 1376
rect 2776 1324 2800 1376
rect 2600 1300 2800 1324
rect 4000 2284 4024 2336
rect 4076 2284 4124 2336
rect 4176 2284 4200 2336
rect 4480 2478 4580 2500
rect 4480 2422 4502 2478
rect 4558 2422 4580 2478
rect 4480 2378 4580 2422
rect 4480 2322 4502 2378
rect 4558 2322 4580 2378
rect 4480 2300 4580 2322
rect 5100 2478 5200 2500
rect 5100 2422 5122 2478
rect 5178 2422 5200 2478
rect 5100 2378 5200 2422
rect 5100 2322 5122 2378
rect 5178 2322 5200 2378
rect 5100 2300 5200 2322
rect 4000 2256 4200 2284
rect 4000 2204 4024 2256
rect 4076 2204 4124 2256
rect 4176 2204 4200 2256
rect 4000 2176 4200 2204
rect 4000 2124 4024 2176
rect 4076 2124 4124 2176
rect 4176 2124 4200 2176
rect 4000 1736 4200 2124
rect 4000 1684 4024 1736
rect 4076 1684 4124 1736
rect 4176 1684 4200 1736
rect 4000 1616 4200 1684
rect 4000 1564 4024 1616
rect 4076 1564 4124 1616
rect 4176 1564 4200 1616
rect 4000 1176 4200 1564
rect 5400 1476 5600 3180
rect 5680 2878 5780 2900
rect 5680 2822 5702 2878
rect 5758 2822 5780 2878
rect 5680 2778 5780 2822
rect 5680 2722 5702 2778
rect 5758 2722 5780 2778
rect 5680 2700 5780 2722
rect 6300 2878 6400 2900
rect 6300 2822 6322 2878
rect 6378 2822 6400 2878
rect 6300 2778 6400 2822
rect 6300 2722 6322 2778
rect 6378 2722 6400 2778
rect 6300 2700 6400 2722
rect 7400 2878 7600 3600
rect 7400 2822 7422 2878
rect 7478 2822 7522 2878
rect 7578 2822 7600 2878
rect 7400 2778 7600 2822
rect 7400 2722 7422 2778
rect 7478 2722 7522 2778
rect 7578 2722 7600 2778
rect 5400 1424 5424 1476
rect 5476 1424 5524 1476
rect 5576 1424 5600 1476
rect 5400 1376 5600 1424
rect 5400 1324 5424 1376
rect 5476 1324 5524 1376
rect 5576 1324 5600 1376
rect 5400 1300 5600 1324
rect 6500 1976 6700 2000
rect 6500 1924 6524 1976
rect 6576 1924 6624 1976
rect 6676 1924 6700 1976
rect 6500 1876 6700 1924
rect 6500 1824 6524 1876
rect 6576 1824 6624 1876
rect 6676 1824 6700 1876
rect 4000 1124 4024 1176
rect 4076 1124 4124 1176
rect 4176 1124 4200 1176
rect 4000 1096 4200 1124
rect 4000 1044 4024 1096
rect 4076 1044 4124 1096
rect 4176 1044 4200 1096
rect 4000 1016 4200 1044
rect 1800 978 1900 1000
rect 1800 922 1822 978
rect 1878 922 1900 978
rect 1800 878 1900 922
rect 1800 822 1822 878
rect 1878 822 1900 878
rect 1800 800 1900 822
rect 2380 978 2480 1000
rect 2380 922 2402 978
rect 2458 922 2480 978
rect 2380 878 2480 922
rect 2380 822 2402 878
rect 2458 822 2480 878
rect 2380 800 2480 822
rect 4000 964 4024 1016
rect 4076 964 4124 1016
rect 4176 964 4200 1016
rect 4000 936 4200 964
rect 4000 884 4024 936
rect 4076 884 4124 936
rect 4176 884 4200 936
rect 4000 856 4200 884
rect 4000 804 4024 856
rect 4076 804 4124 856
rect 4176 804 4200 856
rect 4000 776 4200 804
rect 5700 978 5800 1000
rect 5700 922 5722 978
rect 5778 922 5800 978
rect 5700 878 5800 922
rect 5700 822 5722 878
rect 5778 822 5800 878
rect 5700 800 5800 822
rect 6280 978 6380 1000
rect 6280 922 6302 978
rect 6358 922 6380 978
rect 6280 878 6380 922
rect 6280 822 6302 878
rect 6358 822 6380 878
rect 6280 800 6380 822
rect 4000 724 4024 776
rect 4076 724 4124 776
rect 4176 724 4200 776
rect 4000 696 4200 724
rect 4000 644 4024 696
rect 4076 644 4124 696
rect 4176 644 4200 696
rect 4000 616 4200 644
rect 3000 578 3100 600
rect 3000 522 3022 578
rect 3078 522 3100 578
rect 3000 478 3100 522
rect 3000 422 3022 478
rect 3078 422 3100 478
rect 3000 400 3100 422
rect 3580 578 3680 600
rect 3580 522 3602 578
rect 3658 522 3680 578
rect 3580 478 3680 522
rect 3580 422 3602 478
rect 3658 422 3680 478
rect 3580 400 3680 422
rect 4000 564 4024 616
rect 4076 564 4124 616
rect 4176 564 4200 616
rect 4000 536 4200 564
rect 4000 484 4024 536
rect 4076 484 4124 536
rect 4176 484 4200 536
rect 4000 456 4200 484
rect 4000 404 4024 456
rect 4076 404 4124 456
rect 4176 404 4200 456
rect 4000 376 4200 404
rect 4500 578 4600 600
rect 4500 522 4522 578
rect 4578 522 4600 578
rect 4500 478 4600 522
rect 4500 422 4522 478
rect 4578 422 4600 478
rect 4500 400 4600 422
rect 5080 578 5180 600
rect 5080 522 5102 578
rect 5158 522 5180 578
rect 5080 478 5180 522
rect 5080 422 5102 478
rect 5158 422 5180 478
rect 5080 400 5180 422
rect 4000 324 4024 376
rect 4076 324 4124 376
rect 4176 324 4200 376
rect 4000 296 4200 324
rect 4000 244 4024 296
rect 4076 244 4124 296
rect 4176 244 4200 296
rect 4000 216 4200 244
rect 4000 164 4024 216
rect 4076 164 4124 216
rect 4176 164 4200 216
rect 4000 136 4200 164
rect 1500 96 2300 120
rect 1500 44 2044 96
rect 2096 44 2204 96
rect 2256 44 2300 96
rect 1500 -4 2300 44
rect 1500 -56 2044 -4
rect 2096 -56 2204 -4
rect 2256 -56 2300 -4
rect 1500 -80 2300 -56
rect 4000 84 4024 136
rect 4076 84 4124 136
rect 4176 84 4200 136
rect 6500 120 6700 1824
rect 4000 56 4200 84
rect 4000 4 4024 56
rect 4076 4 4124 56
rect 4176 4 4200 56
rect 4000 -24 4200 4
rect 4000 -76 4024 -24
rect 4076 -76 4124 -24
rect 4176 -76 4200 -24
rect 600 -176 624 -124
rect 676 -176 724 -124
rect 776 -176 800 -124
rect 600 -224 800 -176
rect 600 -276 624 -224
rect 676 -276 724 -224
rect 776 -276 800 -224
rect 600 -300 800 -276
rect 4000 -324 4200 -76
rect 5900 96 6700 120
rect 5900 44 5944 96
rect 5996 44 6104 96
rect 6156 44 6700 96
rect 5900 -4 6700 44
rect 5900 -56 5944 -4
rect 5996 -56 6104 -4
rect 6156 -56 6700 -4
rect 5900 -80 6700 -56
rect 7400 578 7600 2722
rect 7400 522 7422 578
rect 7478 522 7522 578
rect 7578 522 7600 578
rect 7400 478 7600 522
rect 7400 422 7422 478
rect 7478 422 7522 478
rect 7578 422 7600 478
rect 7400 -124 7600 422
rect 7400 -176 7424 -124
rect 7476 -176 7524 -124
rect 7576 -176 7600 -124
rect 7400 -224 7600 -176
rect 7400 -276 7424 -224
rect 7476 -276 7524 -224
rect 7576 -276 7600 -224
rect 7400 -300 7600 -276
rect 7700 2478 7900 3600
rect 7700 2422 7722 2478
rect 7778 2422 7822 2478
rect 7878 2422 7900 2478
rect 7700 2378 7900 2422
rect 7700 2322 7722 2378
rect 7778 2322 7822 2378
rect 7878 2322 7900 2378
rect 7700 978 7900 2322
rect 7700 922 7722 978
rect 7778 922 7822 978
rect 7878 922 7900 978
rect 7700 878 7900 922
rect 7700 822 7722 878
rect 7778 822 7822 878
rect 7878 822 7900 878
rect 7700 -124 7900 822
rect 7700 -176 7724 -124
rect 7776 -176 7824 -124
rect 7876 -176 7900 -124
rect 7700 -224 7900 -176
rect 7700 -276 7724 -224
rect 7776 -276 7824 -224
rect 7876 -276 7900 -224
rect 7700 -300 7900 -276
rect 4000 -376 4024 -324
rect 4076 -376 4124 -324
rect 4176 -376 4200 -324
rect 4000 -424 4200 -376
rect 4000 -476 4024 -424
rect 4076 -476 4124 -424
rect 4176 -476 4200 -424
rect 4000 -500 4200 -476
<< via2 >>
rect 322 2422 378 2478
rect 422 2422 478 2478
rect 322 2322 378 2378
rect 422 2322 478 2378
rect 322 922 378 978
rect 422 922 478 978
rect 322 822 378 878
rect 422 822 478 878
rect 622 2822 678 2878
rect 722 2822 778 2878
rect 622 2722 678 2778
rect 722 2722 778 2778
rect 1822 2876 1878 2878
rect 1822 2824 1824 2876
rect 1824 2824 1876 2876
rect 1876 2824 1878 2876
rect 1822 2822 1878 2824
rect 1822 2776 1878 2778
rect 1822 2724 1824 2776
rect 1824 2724 1876 2776
rect 1876 2724 1878 2776
rect 1822 2722 1878 2724
rect 2422 2876 2478 2878
rect 2422 2824 2424 2876
rect 2424 2824 2476 2876
rect 2476 2824 2478 2876
rect 2422 2822 2478 2824
rect 2422 2776 2478 2778
rect 2422 2724 2424 2776
rect 2424 2724 2476 2776
rect 2476 2724 2478 2776
rect 2422 2722 2478 2724
rect 622 522 678 578
rect 722 522 778 578
rect 622 422 678 478
rect 722 422 778 478
rect 3002 2476 3058 2478
rect 3002 2424 3004 2476
rect 3004 2424 3056 2476
rect 3056 2424 3058 2476
rect 3002 2422 3058 2424
rect 3002 2376 3058 2378
rect 3002 2324 3004 2376
rect 3004 2324 3056 2376
rect 3056 2324 3058 2376
rect 3002 2322 3058 2324
rect 3622 2476 3678 2478
rect 3622 2424 3624 2476
rect 3624 2424 3676 2476
rect 3676 2424 3678 2476
rect 3622 2422 3678 2424
rect 3622 2376 3678 2378
rect 3622 2324 3624 2376
rect 3624 2324 3676 2376
rect 3676 2324 3678 2376
rect 3622 2322 3678 2324
rect 4502 2476 4558 2478
rect 4502 2424 4504 2476
rect 4504 2424 4556 2476
rect 4556 2424 4558 2476
rect 4502 2422 4558 2424
rect 4502 2376 4558 2378
rect 4502 2324 4504 2376
rect 4504 2324 4556 2376
rect 4556 2324 4558 2376
rect 4502 2322 4558 2324
rect 5122 2476 5178 2478
rect 5122 2424 5124 2476
rect 5124 2424 5176 2476
rect 5176 2424 5178 2476
rect 5122 2422 5178 2424
rect 5122 2376 5178 2378
rect 5122 2324 5124 2376
rect 5124 2324 5176 2376
rect 5176 2324 5178 2376
rect 5122 2322 5178 2324
rect 5702 2876 5758 2878
rect 5702 2824 5704 2876
rect 5704 2824 5756 2876
rect 5756 2824 5758 2876
rect 5702 2822 5758 2824
rect 5702 2776 5758 2778
rect 5702 2724 5704 2776
rect 5704 2724 5756 2776
rect 5756 2724 5758 2776
rect 5702 2722 5758 2724
rect 6322 2876 6378 2878
rect 6322 2824 6324 2876
rect 6324 2824 6376 2876
rect 6376 2824 6378 2876
rect 6322 2822 6378 2824
rect 6322 2776 6378 2778
rect 6322 2724 6324 2776
rect 6324 2724 6376 2776
rect 6376 2724 6378 2776
rect 6322 2722 6378 2724
rect 7422 2822 7478 2878
rect 7522 2822 7578 2878
rect 7422 2722 7478 2778
rect 7522 2722 7578 2778
rect 1822 976 1878 978
rect 1822 924 1824 976
rect 1824 924 1876 976
rect 1876 924 1878 976
rect 1822 922 1878 924
rect 1822 876 1878 878
rect 1822 824 1824 876
rect 1824 824 1876 876
rect 1876 824 1878 876
rect 1822 822 1878 824
rect 2402 976 2458 978
rect 2402 924 2404 976
rect 2404 924 2456 976
rect 2456 924 2458 976
rect 2402 922 2458 924
rect 2402 876 2458 878
rect 2402 824 2404 876
rect 2404 824 2456 876
rect 2456 824 2458 876
rect 2402 822 2458 824
rect 5722 976 5778 978
rect 5722 924 5724 976
rect 5724 924 5776 976
rect 5776 924 5778 976
rect 5722 922 5778 924
rect 5722 876 5778 878
rect 5722 824 5724 876
rect 5724 824 5776 876
rect 5776 824 5778 876
rect 5722 822 5778 824
rect 6302 976 6358 978
rect 6302 924 6304 976
rect 6304 924 6356 976
rect 6356 924 6358 976
rect 6302 922 6358 924
rect 6302 876 6358 878
rect 6302 824 6304 876
rect 6304 824 6356 876
rect 6356 824 6358 876
rect 6302 822 6358 824
rect 3022 576 3078 578
rect 3022 524 3024 576
rect 3024 524 3076 576
rect 3076 524 3078 576
rect 3022 522 3078 524
rect 3022 476 3078 478
rect 3022 424 3024 476
rect 3024 424 3076 476
rect 3076 424 3078 476
rect 3022 422 3078 424
rect 3602 576 3658 578
rect 3602 524 3604 576
rect 3604 524 3656 576
rect 3656 524 3658 576
rect 3602 522 3658 524
rect 3602 476 3658 478
rect 3602 424 3604 476
rect 3604 424 3656 476
rect 3656 424 3658 476
rect 3602 422 3658 424
rect 4522 576 4578 578
rect 4522 524 4524 576
rect 4524 524 4576 576
rect 4576 524 4578 576
rect 4522 522 4578 524
rect 4522 476 4578 478
rect 4522 424 4524 476
rect 4524 424 4576 476
rect 4576 424 4578 476
rect 4522 422 4578 424
rect 5102 576 5158 578
rect 5102 524 5104 576
rect 5104 524 5156 576
rect 5156 524 5158 576
rect 5102 522 5158 524
rect 5102 476 5158 478
rect 5102 424 5104 476
rect 5104 424 5156 476
rect 5156 424 5158 476
rect 5102 422 5158 424
rect 7422 522 7478 578
rect 7522 522 7578 578
rect 7422 422 7478 478
rect 7522 422 7578 478
rect 7722 2422 7778 2478
rect 7822 2422 7878 2478
rect 7722 2322 7778 2378
rect 7822 2322 7878 2378
rect 7722 922 7778 978
rect 7822 922 7878 978
rect 7722 822 7778 878
rect 7822 822 7878 878
<< metal3 >>
rect 300 2878 7900 2900
rect 300 2822 622 2878
rect 678 2822 722 2878
rect 778 2822 1822 2878
rect 1878 2822 2422 2878
rect 2478 2822 5702 2878
rect 5758 2822 6322 2878
rect 6378 2822 7422 2878
rect 7478 2822 7522 2878
rect 7578 2822 7900 2878
rect 300 2778 7900 2822
rect 300 2722 622 2778
rect 678 2722 722 2778
rect 778 2722 1822 2778
rect 1878 2722 2422 2778
rect 2478 2722 5702 2778
rect 5758 2722 6322 2778
rect 6378 2722 7422 2778
rect 7478 2722 7522 2778
rect 7578 2722 7900 2778
rect 300 2700 7900 2722
rect 300 2478 7900 2500
rect 300 2422 322 2478
rect 378 2422 422 2478
rect 478 2422 3002 2478
rect 3058 2422 3622 2478
rect 3678 2422 4502 2478
rect 4558 2422 5122 2478
rect 5178 2422 7722 2478
rect 7778 2422 7822 2478
rect 7878 2422 7900 2478
rect 300 2378 7900 2422
rect 300 2322 322 2378
rect 378 2322 422 2378
rect 478 2322 3002 2378
rect 3058 2322 3622 2378
rect 3678 2322 4502 2378
rect 4558 2322 5122 2378
rect 5178 2322 7722 2378
rect 7778 2322 7822 2378
rect 7878 2322 7900 2378
rect 300 2300 7900 2322
rect 300 978 7900 1000
rect 300 922 322 978
rect 378 922 422 978
rect 478 922 1822 978
rect 1878 922 2402 978
rect 2458 922 5722 978
rect 5778 922 6302 978
rect 6358 922 7722 978
rect 7778 922 7822 978
rect 7878 922 7900 978
rect 300 878 7900 922
rect 300 822 322 878
rect 378 822 422 878
rect 478 822 1822 878
rect 1878 822 2402 878
rect 2458 822 5722 878
rect 5778 822 6302 878
rect 6358 822 7722 878
rect 7778 822 7822 878
rect 7878 822 7900 878
rect 300 800 7900 822
rect 300 578 7900 600
rect 300 522 622 578
rect 678 522 722 578
rect 778 522 3022 578
rect 3078 522 3602 578
rect 3658 522 4522 578
rect 4578 522 5102 578
rect 5158 522 7422 578
rect 7478 522 7522 578
rect 7578 522 7900 578
rect 300 478 7900 522
rect 300 422 622 478
rect 678 422 722 478
rect 778 422 3022 478
rect 3078 422 3602 478
rect 3658 422 4522 478
rect 4578 422 5102 478
rect 5158 422 7422 478
rect 7478 422 7522 478
rect 7578 422 7900 478
rect 300 400 7900 422
use sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH  sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_0
timestamp 1770083657
transform 1 0 3345 0 1 2632
box -371 -532 371 532
use sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH  sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_1
timestamp 1770083657
transform 1 0 6045 0 1 732
box -371 -532 371 532
use sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH  sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_2
timestamp 1770083657
transform 1 0 2145 0 1 732
box -371 -532 371 532
use sky130_fd_pr__nfet_g5v0d10v5_SNDLS5  sky130_fd_pr__nfet_g5v0d10v5_SNDLS5_0
timestamp 1770083657
transform 1 0 4845 0 1 2632
box -371 -532 371 532
use sky130_fd_pr__nfet_g5v0d10v5_X57ESK  sky130_fd_pr__nfet_g5v0d10v5_X57ESK_0
timestamp 1770083657
transform 1 0 2145 0 1 2632
box -371 -532 371 532
use sky130_fd_pr__nfet_g5v0d10v5_X57ESK  sky130_fd_pr__nfet_g5v0d10v5_X57ESK_1
timestamp 1770083657
transform 1 0 6045 0 1 2632
box -371 -532 371 532
use sky130_fd_pr__nfet_g5v0d10v5_X57ESK  sky130_fd_pr__nfet_g5v0d10v5_X57ESK_2
timestamp 1770083657
transform 1 0 4845 0 1 732
box -371 -532 371 532
use sky130_fd_pr__nfet_g5v0d10v5_X57ESK  sky130_fd_pr__nfet_g5v0d10v5_X57ESK_3
timestamp 1770083657
transform 1 0 3345 0 1 732
box -371 -532 371 532
<< labels >>
flabel metal1 s 900 1300 1100 1500 0 FreeSans 320 0 0 0 VP
port 1 nsew
flabel metal1 s 900 1800 1100 2000 0 FreeSans 320 0 0 0 VN
port 2 nsew
flabel metal1 s 4060 -460 4160 -360 0 FreeSans 320 0 0 0 S
port 3 nsew
flabel metal1 s 320 -300 420 -200 0 FreeSans 320 0 0 0 D2
port 4 nsew
flabel metal1 s 640 -300 740 -200 0 FreeSans 320 0 0 0 D1
port 5 nsew
flabel metal1 s 1300 -300 1400 -200 0 FreeSans 320 0 0 0 VSS
port 6 nsew
<< end >>
