magic
tech sky130A
magscale 1 2
timestamp 1769150038
<< nwell >>
rect 760 -800 5140 240
<< pwell >>
rect 800 -2440 5100 -800
<< psubdiff >>
rect 2200 -920 3600 -900
rect 2200 -980 2340 -920
rect 3440 -980 3600 -920
rect 2200 -1000 3600 -980
rect 2200 -1700 2220 -1000
rect 1700 -1720 2220 -1700
rect 2280 -1700 2300 -1000
rect 3500 -1700 3520 -1000
rect 2280 -1720 3520 -1700
rect 3580 -1700 3600 -1000
rect 3580 -1720 4200 -1700
rect 1700 -1780 1800 -1720
rect 4100 -1780 4200 -1720
rect 1700 -1800 4200 -1780
rect 1700 -1820 1800 -1800
rect 1700 -2260 1720 -1820
rect 1780 -2260 1800 -1820
rect 1700 -2300 1800 -2260
rect 4100 -1820 4200 -1800
rect 4100 -2260 4120 -1820
rect 4180 -2260 4200 -1820
rect 4100 -2300 4200 -2260
rect 1700 -2320 4200 -2300
rect 1700 -2380 1800 -2320
rect 4100 -2380 4200 -2320
rect 1700 -2400 4200 -2380
<< nsubdiff >>
rect 800 180 5100 200
rect 800 120 900 180
rect 5000 120 5100 180
rect 800 100 5100 120
rect 800 80 900 100
rect 800 -580 820 80
rect 880 -580 900 80
rect 800 -600 900 -580
rect 5000 80 5100 100
rect 5000 -580 5020 80
rect 5080 -580 5100 80
rect 5000 -600 5100 -580
rect 800 -620 5100 -600
rect 800 -680 900 -620
rect 5000 -680 5100 -620
rect 800 -700 5100 -680
<< psubdiffcont >>
rect 2340 -980 3440 -920
rect 2220 -1720 2280 -1000
rect 3520 -1720 3580 -1000
rect 1800 -1780 4100 -1720
rect 1720 -2260 1780 -1820
rect 4120 -2260 4180 -1820
rect 1800 -2380 4100 -2320
<< nsubdiffcont >>
rect 900 120 5000 180
rect 820 -580 880 80
rect 5020 -580 5080 80
rect 900 -680 5000 -620
<< locali >>
rect 760 180 5140 360
rect 760 160 820 180
rect 800 120 820 160
rect 880 120 900 180
rect 5000 120 5020 180
rect 5080 160 5140 180
rect 5080 120 5100 160
rect 800 100 5100 120
rect 800 80 900 100
rect 800 -580 820 80
rect 880 -580 900 80
rect 960 -400 1080 0
rect 1280 -400 1380 100
rect 1920 -400 2040 100
rect 2240 -440 2340 0
rect 2560 -400 2680 100
rect 3200 -400 3320 100
rect 3540 -440 3640 0
rect 3840 -400 3960 100
rect 4260 -400 4380 0
rect 4500 -400 4600 100
rect 5000 80 5100 100
rect 1080 -500 2860 -440
rect 3020 -500 4800 -440
rect 800 -600 900 -580
rect 5000 -580 5020 80
rect 5080 -580 5100 80
rect 5000 -600 5100 -580
rect 800 -620 5100 -600
rect 800 -680 820 -620
rect 880 -680 900 -620
rect 5000 -680 5020 -620
rect 5080 -680 5100 -620
rect 800 -700 5100 -680
rect 2200 -920 3600 -900
rect 2200 -980 2220 -920
rect 2280 -980 2340 -920
rect 3440 -980 3520 -920
rect 3580 -980 3600 -920
rect 2200 -1000 3600 -980
rect 2200 -1700 2220 -1000
rect 1700 -1720 2220 -1700
rect 2280 -1700 2300 -1000
rect 3114 -1078 3150 -1069
rect 3230 -1077 3254 -1069
rect 2680 -1400 2720 -1080
rect 2680 -1416 2718 -1400
rect 3134 -1416 3150 -1078
rect 3500 -1700 3520 -1000
rect 2280 -1720 3520 -1700
rect 3580 -1700 3600 -1000
rect 3580 -1720 4200 -1700
rect 1700 -1780 1720 -1720
rect 1780 -1780 1800 -1720
rect 4100 -1780 4120 -1720
rect 4180 -1780 4200 -1720
rect 1700 -1800 4200 -1780
rect 1700 -1820 1800 -1800
rect 1700 -2260 1720 -1820
rect 1780 -2260 1800 -1820
rect 4100 -1820 4200 -1800
rect 1700 -2300 1800 -2260
rect 2240 -2300 2360 -1980
rect 2860 -2300 3020 -1980
rect 3520 -2300 3640 -1980
rect 4100 -2260 4120 -1820
rect 4180 -2260 4200 -1820
rect 4100 -2300 4200 -2260
rect 800 -2320 5140 -2300
rect 800 -2380 1720 -2320
rect 1780 -2380 1800 -2320
rect 4100 -2380 4120 -2320
rect 4180 -2380 5140 -2320
rect 800 -2500 5140 -2380
<< viali >>
rect 820 120 880 180
rect 5020 120 5080 180
rect 820 -680 880 -620
rect 5020 -680 5080 -620
rect 2220 -980 2280 -920
rect 3520 -980 3580 -920
rect 1720 -1780 1780 -1720
rect 4120 -1780 4180 -1720
rect 1720 -2380 1780 -2320
rect 4120 -2380 4180 -2320
<< metal1 >>
rect 760 180 5140 360
rect 760 160 820 180
rect 800 120 820 160
rect 880 120 5020 180
rect 5080 160 5140 180
rect 5080 120 5100 160
rect 800 100 5100 120
rect 800 -600 900 100
rect 960 -60 1080 0
rect 960 -140 980 -60
rect 1060 -140 1080 -60
rect 960 -180 1080 -140
rect 960 -260 980 -180
rect 1060 -260 1080 -180
rect 960 -400 1080 -260
rect 1500 -60 1620 0
rect 1500 -140 1520 -60
rect 1600 -140 1620 -60
rect 1500 -180 1620 -140
rect 1500 -260 1520 -180
rect 1600 -260 1620 -180
rect 1500 -400 1620 -260
rect 1680 -60 1800 0
rect 1680 -140 1700 -60
rect 1780 -140 1800 -60
rect 1680 -180 1800 -140
rect 1680 -260 1700 -180
rect 1780 -260 1800 -180
rect 1680 -300 1800 -260
rect 1680 -380 1700 -300
rect 1780 -380 1800 -300
rect 1680 -400 1800 -380
rect 2220 -80 2260 0
rect 2340 -80 2380 0
rect 2220 -100 2380 -80
rect 2220 -180 2260 -100
rect 2340 -180 2380 -100
rect 2220 -200 2380 -180
rect 2220 -280 2260 -200
rect 2340 -280 2380 -200
rect 2220 -300 2380 -280
rect 2220 -380 2260 -300
rect 2340 -380 2380 -300
rect 2220 -400 2380 -380
rect 3500 -80 3540 0
rect 3620 -80 3700 0
rect 3500 -100 3700 -80
rect 3500 -180 3540 -100
rect 3620 -180 3700 -100
rect 3500 -200 3700 -180
rect 3500 -280 3540 -200
rect 3620 -280 3700 -200
rect 3500 -300 3700 -280
rect 3500 -380 3540 -300
rect 3620 -380 3700 -300
rect 3500 -400 3700 -380
rect 4080 -60 4200 0
rect 4080 -140 4100 -60
rect 4180 -140 4200 -60
rect 4080 -180 4200 -140
rect 4080 -260 4100 -180
rect 4180 -260 4200 -180
rect 4080 -300 4200 -260
rect 4080 -380 4100 -300
rect 4180 -380 4200 -300
rect 4080 -400 4200 -380
rect 4260 -60 4380 0
rect 4260 -140 4280 -60
rect 4360 -140 4380 -60
rect 4260 -180 4380 -140
rect 4260 -260 4280 -180
rect 4360 -260 4380 -180
rect 4260 -300 4380 -260
rect 4260 -380 4280 -300
rect 4360 -380 4380 -300
rect 4260 -400 4380 -380
rect 4800 -60 4920 0
rect 4800 -140 4820 -60
rect 4900 -140 4920 -60
rect 4800 -180 4920 -140
rect 4800 -260 4820 -180
rect 4900 -260 4920 -180
rect 4800 -300 4920 -260
rect 4800 -380 4820 -300
rect 4900 -380 4920 -300
rect 4800 -400 4920 -380
rect 5000 -600 5100 100
rect 800 -620 5100 -600
rect 800 -680 820 -620
rect 880 -680 5020 -620
rect 5080 -680 5100 -620
rect 800 -700 5100 -680
rect 2200 -920 3600 -900
rect 2200 -980 2220 -920
rect 2280 -980 3520 -920
rect 3580 -980 3600 -920
rect 2200 -1000 3600 -980
rect 2200 -1700 2300 -1000
rect 2360 -1120 2440 -1060
rect 2420 -1180 2440 -1120
rect 2360 -1220 2440 -1180
rect 2420 -1280 2440 -1220
rect 2360 -1320 2440 -1280
rect 2420 -1380 2440 -1320
rect 2360 -1400 2440 -1380
rect 2560 -1080 2740 -1060
rect 2560 -1180 2600 -1080
rect 2700 -1180 2740 -1080
rect 2560 -1260 2740 -1180
rect 2560 -1360 2600 -1260
rect 2700 -1360 2740 -1260
rect 2560 -1400 2740 -1360
rect 2860 -1100 2980 -1060
rect 2860 -1180 2880 -1100
rect 2960 -1180 2980 -1100
rect 2860 -1200 2980 -1180
rect 2860 -1280 2880 -1200
rect 2960 -1280 2980 -1200
rect 2860 -1300 2980 -1280
rect 2860 -1380 2880 -1300
rect 2960 -1380 2980 -1300
rect 2860 -1400 2980 -1380
rect 3100 -1080 3280 -1060
rect 3100 -1180 3140 -1080
rect 3240 -1180 3280 -1080
rect 3100 -1260 3280 -1180
rect 3100 -1360 3140 -1260
rect 3240 -1360 3280 -1260
rect 3100 -1400 3280 -1360
rect 3380 -1120 3460 -1060
rect 3380 -1180 3400 -1120
rect 3380 -1220 3460 -1180
rect 3380 -1280 3400 -1220
rect 3380 -1320 3460 -1280
rect 3380 -1380 3400 -1320
rect 3380 -1400 3460 -1380
rect 2460 -1480 2560 -1440
rect 3280 -1480 3380 -1440
rect 2420 -1500 2600 -1480
rect 2420 -1560 2440 -1500
rect 2500 -1560 2540 -1500
rect 2420 -1580 2600 -1560
rect 2420 -1640 2440 -1580
rect 2500 -1640 2540 -1580
rect 2420 -1660 2600 -1640
rect 3240 -1500 3420 -1480
rect 3300 -1560 3320 -1500
rect 3380 -1560 3420 -1500
rect 3240 -1580 3420 -1560
rect 3300 -1640 3320 -1580
rect 3380 -1640 3420 -1580
rect 3240 -1660 3420 -1640
rect 3500 -1700 3600 -1000
rect 1700 -1720 4200 -1700
rect 1700 -1780 1720 -1720
rect 1780 -1780 4120 -1720
rect 4180 -1780 4200 -1720
rect 1700 -1800 4200 -1780
rect 1700 -2300 1800 -1800
rect 2060 -1900 2080 -1840
rect 2140 -1900 2180 -1840
rect 2240 -1900 2360 -1840
rect 2420 -1900 2460 -1840
rect 2520 -1900 2540 -1840
rect 2060 -1920 2540 -1900
rect 2700 -1900 2720 -1840
rect 2780 -1900 2800 -1840
rect 2860 -1900 2880 -1840
rect 3000 -1900 3020 -1840
rect 3080 -1900 3100 -1840
rect 3160 -1900 3180 -1840
rect 2700 -1920 3180 -1900
rect 3340 -1900 3360 -1840
rect 3420 -1900 3460 -1840
rect 3520 -1900 3640 -1840
rect 3700 -1900 3740 -1840
rect 3800 -1900 3820 -1840
rect 3340 -1920 3820 -1900
rect 1940 -2020 2100 -2000
rect 1940 -2140 1960 -2020
rect 2080 -2140 2100 -2020
rect 1940 -2160 2100 -2140
rect 2420 -2020 2580 -2000
rect 2420 -2140 2440 -2020
rect 2560 -2140 2580 -2020
rect 2420 -2160 2580 -2140
rect 2640 -2040 2800 -1960
rect 2640 -2160 2660 -2040
rect 2780 -2160 2800 -2040
rect 2640 -2180 2800 -2160
rect 3080 -2040 3240 -1980
rect 3080 -2160 3100 -2040
rect 3220 -2160 3240 -2040
rect 3300 -2020 3460 -2000
rect 3300 -2140 3320 -2020
rect 3440 -2140 3460 -2020
rect 3300 -2160 3460 -2140
rect 3780 -2020 3940 -2000
rect 3780 -2140 3800 -2020
rect 3920 -2140 3940 -2020
rect 3780 -2160 3940 -2140
rect 3080 -2180 3240 -2160
rect 4100 -2300 4200 -1800
rect 800 -2320 5140 -2300
rect 800 -2380 1720 -2320
rect 1780 -2380 4120 -2320
rect 4180 -2380 5140 -2320
rect 800 -2500 5140 -2380
rect 1100 -2800 1300 -2600
rect 1600 -2800 1800 -2600
rect 2840 -2820 3040 -2620
rect 4100 -2800 4300 -2600
rect 4600 -2800 4800 -2600
<< via1 >>
rect 980 -140 1060 -60
rect 980 -260 1060 -180
rect 1520 -140 1600 -60
rect 1520 -260 1600 -180
rect 1700 -140 1780 -60
rect 1700 -260 1780 -180
rect 1700 -380 1780 -300
rect 2260 -80 2340 0
rect 2260 -180 2340 -100
rect 2260 -280 2340 -200
rect 2260 -380 2340 -300
rect 3540 -80 3620 0
rect 3540 -180 3620 -100
rect 3540 -280 3620 -200
rect 3540 -380 3620 -300
rect 4100 -140 4180 -60
rect 4100 -260 4180 -180
rect 4100 -380 4180 -300
rect 4280 -140 4360 -60
rect 4280 -260 4360 -180
rect 4280 -380 4360 -300
rect 4820 -140 4900 -60
rect 4820 -260 4900 -180
rect 4820 -380 4900 -300
rect 2360 -1180 2420 -1120
rect 2360 -1280 2420 -1220
rect 2360 -1380 2420 -1320
rect 2600 -1180 2700 -1080
rect 2600 -1360 2700 -1260
rect 2880 -1180 2960 -1100
rect 2880 -1280 2960 -1200
rect 2880 -1380 2960 -1300
rect 3140 -1180 3240 -1080
rect 3140 -1360 3240 -1260
rect 3400 -1180 3460 -1120
rect 3400 -1280 3460 -1220
rect 3400 -1380 3460 -1320
rect 2440 -1560 2500 -1500
rect 2540 -1560 2600 -1500
rect 2440 -1640 2500 -1580
rect 2540 -1640 2600 -1580
rect 3240 -1560 3300 -1500
rect 3320 -1560 3380 -1500
rect 3240 -1640 3300 -1580
rect 3320 -1640 3380 -1580
rect 2080 -1900 2140 -1840
rect 2180 -1900 2240 -1840
rect 2360 -1900 2420 -1840
rect 2460 -1900 2520 -1840
rect 2720 -1900 2780 -1840
rect 2800 -1900 2860 -1840
rect 2880 -1900 3000 -1840
rect 3020 -1900 3080 -1840
rect 3100 -1900 3160 -1840
rect 3360 -1900 3420 -1840
rect 3460 -1900 3520 -1840
rect 3640 -1900 3700 -1840
rect 3740 -1900 3800 -1840
rect 1960 -2140 2080 -2020
rect 2440 -2140 2560 -2020
rect 2660 -2160 2780 -2040
rect 3100 -2160 3220 -2040
rect 3320 -2140 3440 -2020
rect 3800 -2140 3920 -2020
<< metal2 >>
rect 960 -60 1080 0
rect 960 -140 980 -60
rect 1060 -140 1080 -60
rect 960 -180 1080 -140
rect 960 -260 980 -180
rect 1060 -260 1080 -180
rect 960 -300 1080 -260
rect 960 -380 980 -300
rect 1060 -380 1080 -300
rect 960 -400 1080 -380
rect 1500 -60 1620 0
rect 1500 -140 1520 -60
rect 1600 -140 1620 -60
rect 1500 -180 1620 -140
rect 1500 -260 1520 -180
rect 1600 -260 1620 -180
rect 1500 -300 1620 -260
rect 1500 -380 1520 -300
rect 1600 -380 1620 -300
rect 1500 -400 1620 -380
rect 1680 -60 1800 0
rect 1680 -140 1700 -60
rect 1780 -140 1800 -60
rect 1680 -180 1800 -140
rect 1680 -260 1700 -180
rect 1780 -260 1800 -180
rect 1680 -300 1800 -260
rect 1680 -380 1700 -300
rect 1780 -380 1800 -300
rect 1680 -400 1800 -380
rect 2200 -20 2260 0
rect 2340 -20 2400 0
rect 2200 -80 2220 -20
rect 2380 -80 2400 -20
rect 2200 -100 2400 -80
rect 2200 -120 2260 -100
rect 2340 -120 2400 -100
rect 2200 -180 2220 -120
rect 2380 -180 2400 -120
rect 2200 -200 2400 -180
rect 2200 -220 2260 -200
rect 2340 -220 2400 -200
rect 2200 -280 2220 -220
rect 2380 -280 2400 -220
rect 2200 -300 2400 -280
rect 2200 -320 2260 -300
rect 2340 -320 2400 -300
rect 2200 -380 2220 -320
rect 2380 -380 2400 -320
rect 2200 -400 2400 -380
rect 3500 -20 3540 0
rect 3620 -20 3700 0
rect 3500 -80 3520 -20
rect 3680 -80 3700 -20
rect 3500 -100 3700 -80
rect 3500 -120 3540 -100
rect 3620 -120 3700 -100
rect 3500 -180 3520 -120
rect 3680 -180 3700 -120
rect 3500 -200 3700 -180
rect 3500 -220 3540 -200
rect 3620 -220 3700 -200
rect 3500 -280 3520 -220
rect 3680 -280 3700 -220
rect 3500 -300 3700 -280
rect 3500 -320 3540 -300
rect 3620 -320 3700 -300
rect 3500 -380 3520 -320
rect 3680 -380 3700 -320
rect 3500 -400 3700 -380
rect 4080 -60 4200 0
rect 4080 -140 4100 -60
rect 4180 -140 4200 -60
rect 4080 -180 4200 -140
rect 4080 -260 4100 -180
rect 4180 -260 4200 -180
rect 4080 -300 4200 -260
rect 4080 -380 4100 -300
rect 4180 -380 4200 -300
rect 4080 -400 4200 -380
rect 4260 -60 4380 0
rect 4260 -140 4280 -60
rect 4360 -140 4380 -60
rect 4260 -180 4380 -140
rect 4260 -260 4280 -180
rect 4360 -260 4380 -180
rect 4260 -300 4380 -260
rect 4260 -380 4280 -300
rect 4360 -380 4380 -300
rect 4260 -400 4380 -380
rect 4800 -60 4920 0
rect 4800 -140 4820 -60
rect 4900 -140 4920 -60
rect 4800 -180 4920 -140
rect 4800 -260 4820 -180
rect 4900 -260 4920 -180
rect 4800 -300 4920 -260
rect 4800 -380 4820 -300
rect 4900 -380 4920 -300
rect 4800 -400 4920 -380
rect 2240 -580 2360 -400
rect 2240 -660 2260 -580
rect 2340 -660 2360 -580
rect 2240 -700 2360 -660
rect 2240 -780 2260 -700
rect 2340 -780 2360 -700
rect 2240 -820 2360 -780
rect 2240 -900 2260 -820
rect 2340 -900 2360 -820
rect 2240 -920 2360 -900
rect 2860 -660 2980 -620
rect 3520 -660 3640 -400
rect 2860 -780 3640 -660
rect 2360 -1120 2440 -1060
rect 2420 -1180 2440 -1120
rect 2360 -1220 2440 -1180
rect 2420 -1280 2440 -1220
rect 2360 -1320 2440 -1280
rect 2420 -1380 2440 -1320
rect 2360 -1400 2440 -1380
rect 2560 -1080 2740 -1060
rect 2560 -1180 2600 -1080
rect 2700 -1180 2740 -1080
rect 2560 -1260 2740 -1180
rect 2560 -1360 2600 -1260
rect 2700 -1360 2740 -1260
rect 2560 -1400 2740 -1360
rect 2860 -1100 2980 -780
rect 3520 -800 3640 -780
rect 2860 -1180 2880 -1100
rect 2960 -1180 2980 -1100
rect 2860 -1200 2980 -1180
rect 2860 -1280 2880 -1200
rect 2960 -1280 2980 -1200
rect 2860 -1300 2980 -1280
rect 2860 -1380 2880 -1300
rect 2960 -1380 2980 -1300
rect 2860 -1400 2980 -1380
rect 3100 -1080 3280 -1060
rect 3100 -1180 3140 -1080
rect 3240 -1180 3280 -1080
rect 3100 -1260 3280 -1180
rect 3100 -1360 3140 -1260
rect 3240 -1360 3280 -1260
rect 3100 -1400 3280 -1360
rect 3380 -1120 3460 -1060
rect 3380 -1180 3400 -1120
rect 3380 -1220 3460 -1180
rect 3380 -1280 3400 -1220
rect 3380 -1320 3460 -1280
rect 3380 -1380 3400 -1320
rect 3380 -1400 3460 -1380
rect 1600 -1560 2440 -1500
rect 2500 -1560 2540 -1500
rect 2600 -1560 3240 -1500
rect 3300 -1560 3320 -1500
rect 3380 -1560 3420 -1500
rect 1600 -1580 3420 -1560
rect 1600 -1640 2440 -1580
rect 2500 -1640 2540 -1580
rect 2600 -1640 3240 -1580
rect 3300 -1640 3320 -1580
rect 3380 -1640 3420 -1580
rect 1600 -1680 3420 -1640
rect 1100 -1840 1300 -1820
rect 1100 -1900 1120 -1840
rect 1180 -1900 1220 -1840
rect 1280 -1900 1300 -1840
rect 1100 -1940 1300 -1900
rect 1100 -2000 1120 -1940
rect 1180 -2000 1220 -1940
rect 1280 -2000 1300 -1940
rect 1100 -2800 1300 -2000
rect 1600 -2800 1800 -1680
rect 2060 -1840 2540 -1820
rect 2060 -1900 2080 -1840
rect 2140 -1900 2180 -1840
rect 2240 -1900 2360 -1840
rect 2420 -1900 2460 -1840
rect 2520 -1900 2540 -1840
rect 2060 -1940 2540 -1900
rect 2700 -1840 3180 -1820
rect 2700 -1900 2720 -1840
rect 2780 -1900 2800 -1840
rect 2860 -1900 2880 -1840
rect 3000 -1900 3020 -1840
rect 3080 -1900 3100 -1840
rect 3160 -1900 3180 -1840
rect 2700 -1940 3180 -1900
rect 3340 -1840 3820 -1820
rect 3340 -1900 3360 -1840
rect 3420 -1900 3460 -1840
rect 3520 -1900 3640 -1840
rect 3700 -1900 3740 -1840
rect 3800 -1900 3820 -1840
rect 3340 -1940 3820 -1900
rect 1940 -2020 2100 -2000
rect 1940 -2140 1960 -2020
rect 2080 -2140 2100 -2020
rect 1940 -2160 2100 -2140
rect 2420 -2020 2580 -2000
rect 2420 -2140 2440 -2020
rect 2560 -2140 2580 -2020
rect 2420 -2160 2580 -2140
rect 2640 -2040 2800 -1980
rect 2640 -2160 2660 -2040
rect 2780 -2160 2800 -2040
rect 2640 -2180 2800 -2160
rect 2840 -2820 3040 -1940
rect 3080 -2040 3240 -1980
rect 3080 -2160 3100 -2040
rect 3220 -2160 3240 -2040
rect 3300 -2020 3460 -2000
rect 3300 -2140 3320 -2020
rect 3440 -2140 3460 -2020
rect 3300 -2160 3460 -2140
rect 3780 -2020 3940 -2000
rect 3780 -2140 3800 -2020
rect 3920 -2140 3940 -2020
rect 3780 -2160 3940 -2140
rect 3080 -2180 3240 -2160
rect 4100 -2800 4300 -1500
<< via2 >>
rect 980 -140 1060 -60
rect 980 -260 1060 -180
rect 980 -380 1060 -300
rect 1520 -140 1600 -60
rect 1520 -260 1600 -180
rect 1520 -380 1600 -300
rect 1700 -140 1780 -60
rect 1700 -260 1780 -180
rect 1700 -380 1780 -300
rect 2220 -80 2260 -20
rect 2260 -80 2280 -20
rect 2320 -80 2340 -20
rect 2340 -80 2380 -20
rect 2220 -180 2260 -120
rect 2260 -180 2280 -120
rect 2320 -180 2340 -120
rect 2340 -180 2380 -120
rect 2220 -280 2260 -220
rect 2260 -280 2280 -220
rect 2320 -280 2340 -220
rect 2340 -280 2380 -220
rect 2220 -380 2260 -320
rect 2260 -380 2280 -320
rect 2320 -380 2340 -320
rect 2340 -380 2380 -320
rect 3520 -80 3540 -20
rect 3540 -80 3580 -20
rect 3620 -80 3680 -20
rect 3520 -180 3540 -120
rect 3540 -180 3580 -120
rect 3620 -180 3680 -120
rect 3520 -280 3540 -220
rect 3540 -280 3580 -220
rect 3620 -280 3680 -220
rect 3520 -380 3540 -320
rect 3540 -380 3580 -320
rect 3620 -380 3680 -320
rect 4100 -140 4180 -60
rect 4100 -380 4180 -300
rect 4280 -140 4360 -60
rect 4280 -260 4360 -180
rect 4280 -380 4360 -300
rect 4820 -140 4900 -60
rect 4820 -260 4900 -180
rect 4820 -380 4900 -300
rect 2260 -660 2340 -580
rect 2260 -780 2340 -700
rect 2260 -900 2340 -820
rect 2360 -1180 2420 -1120
rect 2360 -1280 2420 -1220
rect 2360 -1380 2420 -1320
rect 2600 -1180 2700 -1080
rect 2600 -1360 2700 -1260
rect 3140 -1180 3240 -1080
rect 3140 -1360 3240 -1260
rect 3400 -1180 3460 -1120
rect 3400 -1280 3460 -1220
rect 3400 -1380 3460 -1320
rect 1120 -1900 1180 -1840
rect 1220 -1900 1280 -1840
rect 1120 -2000 1180 -1940
rect 1220 -2000 1280 -1940
rect 2080 -1900 2140 -1840
rect 2180 -1900 2240 -1840
rect 2360 -1900 2420 -1840
rect 2460 -1900 2520 -1840
rect 3360 -1900 3420 -1840
rect 3460 -1900 3520 -1840
rect 3640 -1900 3700 -1840
rect 3740 -1900 3800 -1840
rect 1960 -2140 2080 -2020
rect 2440 -2140 2560 -2020
rect 2660 -2160 2780 -2040
rect 3100 -2160 3220 -2040
rect 3320 -2140 3440 -2020
rect 3800 -2140 3920 -2020
<< metal3 >>
rect 960 -60 1080 0
rect 960 -140 980 -60
rect 1060 -140 1080 -60
rect 960 -180 1080 -140
rect 960 -260 980 -180
rect 1060 -260 1080 -180
rect 960 -300 1080 -260
rect 960 -380 980 -300
rect 1060 -380 1080 -300
rect 960 -400 1080 -380
rect 1500 -60 1620 0
rect 1500 -140 1520 -60
rect 1600 -140 1620 -60
rect 1500 -180 1620 -140
rect 1500 -260 1520 -180
rect 1600 -260 1620 -180
rect 1500 -300 1620 -260
rect 1500 -380 1520 -300
rect 1600 -380 1620 -300
rect 1500 -400 1620 -380
rect 1680 -60 1800 0
rect 1680 -140 1700 -60
rect 1780 -140 1800 -60
rect 1680 -180 1800 -140
rect 1680 -260 1700 -180
rect 1780 -260 1800 -180
rect 1680 -300 1800 -260
rect 1680 -380 1700 -300
rect 1780 -380 1800 -300
rect 1680 -400 1800 -380
rect 2200 -20 3100 0
rect 2200 -80 2220 -20
rect 2280 -80 2320 -20
rect 2380 -80 3000 -20
rect 2200 -100 3000 -80
rect 3080 -100 3100 -20
rect 2200 -120 3100 -100
rect 2200 -180 2220 -120
rect 2280 -180 2320 -120
rect 2380 -180 2400 -120
rect 2200 -220 2400 -180
rect 2200 -280 2220 -220
rect 2280 -280 2320 -220
rect 2380 -280 2400 -220
rect 2200 -320 2400 -280
rect 2200 -380 2220 -320
rect 2280 -380 2320 -320
rect 2380 -380 2400 -320
rect 2200 -400 2400 -380
rect 2800 -200 2920 -180
rect 2800 -280 2820 -200
rect 2900 -280 2920 -200
rect 2980 -200 3000 -120
rect 3080 -200 3100 -120
rect 2980 -220 3100 -200
rect 3500 -20 3700 0
rect 3500 -80 3520 -20
rect 3580 -80 3620 -20
rect 3680 -80 3700 -20
rect 3500 -120 3700 -80
rect 3500 -180 3520 -120
rect 3580 -180 3620 -120
rect 3680 -180 3700 -120
rect 3500 -220 3700 -180
rect 3500 -280 3520 -220
rect 3580 -280 3620 -220
rect 3680 -280 3700 -220
rect 2800 -300 3700 -280
rect 2800 -380 2820 -300
rect 2900 -320 3700 -300
rect 2900 -380 3520 -320
rect 3580 -380 3620 -320
rect 3680 -380 3700 -320
rect 2800 -400 3700 -380
rect 4080 -60 4200 0
rect 4080 -140 4100 -60
rect 4180 -140 4200 -60
rect 4080 -180 4200 -140
rect 4080 -260 4100 -180
rect 4180 -260 4200 -180
rect 4080 -300 4200 -260
rect 4080 -380 4100 -300
rect 4180 -380 4200 -300
rect 4080 -400 4200 -380
rect 4260 -60 4380 0
rect 4260 -140 4280 -60
rect 4360 -140 4380 -60
rect 4260 -180 4380 -140
rect 4260 -260 4280 -180
rect 4360 -260 4380 -180
rect 4260 -300 4380 -260
rect 4260 -380 4280 -300
rect 4360 -380 4380 -300
rect 4260 -400 4380 -380
rect 4800 -60 4920 0
rect 4800 -140 4820 -60
rect 4900 -140 4920 -60
rect 4800 -180 4920 -140
rect 4800 -260 4820 -180
rect 4900 -260 4920 -180
rect 4800 -300 4920 -260
rect 4800 -380 4820 -300
rect 4900 -380 4920 -300
rect 4800 -400 4920 -380
rect 2240 -580 2360 -560
rect 2240 -660 2260 -580
rect 2340 -660 2360 -580
rect 2240 -700 2360 -660
rect 2240 -780 2260 -700
rect 2340 -780 2360 -700
rect 2240 -800 2360 -780
rect 2240 -820 3500 -800
rect 2240 -900 2260 -820
rect 2340 -900 3500 -820
rect 2240 -920 3500 -900
rect 2320 -1120 2440 -920
rect 2320 -1180 2360 -1120
rect 2420 -1180 2440 -1120
rect 2320 -1220 2440 -1180
rect 2320 -1280 2360 -1220
rect 2420 -1280 2440 -1220
rect 2320 -1320 2440 -1280
rect 2320 -1380 2360 -1320
rect 2420 -1380 2440 -1320
rect 2320 -1420 2440 -1380
rect 2560 -1080 2740 -1060
rect 2560 -1180 2600 -1080
rect 2700 -1180 2740 -1080
rect 2560 -1260 2740 -1180
rect 2560 -1360 2600 -1260
rect 2700 -1360 2740 -1260
rect 2560 -1400 2740 -1360
rect 3100 -1080 3280 -1060
rect 3100 -1180 3140 -1080
rect 3240 -1180 3280 -1080
rect 3100 -1260 3280 -1180
rect 3100 -1360 3140 -1260
rect 3240 -1360 3280 -1260
rect 3100 -1400 3280 -1360
rect 3380 -1120 3500 -920
rect 3380 -1180 3400 -1120
rect 3460 -1180 3500 -1120
rect 3380 -1220 3500 -1180
rect 3380 -1280 3400 -1220
rect 3460 -1280 3500 -1220
rect 3380 -1320 3500 -1280
rect 3380 -1380 3400 -1320
rect 3460 -1380 3500 -1320
rect 3380 -1420 3500 -1380
rect 1100 -1840 3880 -1820
rect 1100 -1900 1120 -1840
rect 1180 -1900 1220 -1840
rect 1280 -1900 2080 -1840
rect 2140 -1900 2180 -1840
rect 2240 -1900 2360 -1840
rect 2420 -1900 2460 -1840
rect 2520 -1900 3360 -1840
rect 3420 -1900 3460 -1840
rect 3520 -1900 3640 -1840
rect 3700 -1900 3740 -1840
rect 3800 -1900 3880 -1840
rect 1100 -1940 3880 -1900
rect 1100 -2000 1120 -1940
rect 1180 -2000 1220 -1940
rect 1280 -2000 1300 -1940
rect 1100 -2020 1300 -2000
rect 1940 -2020 2100 -2000
rect 1940 -2140 1960 -2020
rect 2080 -2140 2100 -2020
rect 1940 -2160 2100 -2140
rect 2420 -2020 2580 -2000
rect 2420 -2140 2440 -2020
rect 2560 -2140 2580 -2020
rect 2420 -2160 2580 -2140
rect 2640 -2040 2800 -2000
rect 2640 -2160 2660 -2040
rect 2780 -2160 2800 -2040
rect 2640 -2180 2800 -2160
rect 3080 -2040 3240 -2000
rect 3080 -2160 3100 -2040
rect 3220 -2160 3240 -2040
rect 3300 -2020 3460 -2000
rect 3300 -2140 3320 -2020
rect 3440 -2140 3460 -2020
rect 3300 -2160 3460 -2140
rect 3780 -2020 3940 -2000
rect 3780 -2140 3800 -2020
rect 3920 -2140 3940 -2020
rect 3780 -2160 3940 -2140
rect 3080 -2180 3240 -2160
<< via3 >>
rect 980 -140 1060 -60
rect 980 -260 1060 -180
rect 980 -380 1060 -300
rect 1520 -140 1600 -60
rect 1520 -260 1600 -180
rect 1520 -380 1600 -300
rect 1700 -140 1780 -60
rect 1700 -260 1780 -180
rect 1700 -380 1780 -300
rect 3000 -100 3080 -20
rect 2820 -280 2900 -200
rect 3000 -200 3080 -120
rect 2820 -380 2900 -300
rect 4100 -140 4180 -60
rect 4100 -260 4180 -180
rect 4100 -380 4180 -300
rect 4280 -140 4360 -60
rect 4280 -260 4360 -180
rect 4280 -380 4360 -300
rect 4820 -140 4900 -60
rect 4820 -260 4900 -180
rect 4820 -380 4900 -300
rect 2600 -1180 2700 -1080
rect 2600 -1360 2700 -1260
rect 3140 -1180 3240 -1080
rect 3140 -1360 3240 -1260
rect 1960 -2140 2080 -2020
rect 2440 -2140 2560 -2020
rect 2660 -2160 2780 -2040
rect 3100 -2160 3220 -2040
rect 3320 -2140 3440 -2020
rect 3800 -2140 3920 -2020
<< metal4 >>
rect 960 -60 1080 0
rect 960 -140 980 -60
rect 1060 -140 1080 -60
rect 960 -180 1080 -140
rect 960 -260 980 -180
rect 1060 -260 1080 -180
rect 960 -300 1080 -260
rect 960 -380 980 -300
rect 1060 -380 1080 -300
rect 960 -760 1080 -380
rect 1500 -60 1620 0
rect 1500 -140 1520 -60
rect 1600 -140 1620 -60
rect 1500 -180 1620 -140
rect 1500 -260 1520 -180
rect 1600 -260 1620 -180
rect 1500 -300 1620 -260
rect 1500 -380 1520 -300
rect 1600 -380 1620 -300
rect 1500 -760 1620 -380
rect 1680 -60 1800 0
rect 1680 -140 1700 -60
rect 1780 -140 1800 -60
rect 1680 -180 1800 -140
rect 1680 -260 1700 -180
rect 1780 -260 1800 -180
rect 1680 -300 1800 -260
rect 1680 -380 1700 -300
rect 1780 -380 1800 -300
rect 1680 -580 1800 -380
rect 2800 -200 2920 0
rect 2800 -280 2820 -200
rect 2900 -280 2920 -200
rect 2800 -300 2920 -280
rect 2800 -380 2820 -300
rect 2900 -380 2920 -300
rect 2800 -580 2920 -380
rect 1680 -700 2920 -580
rect 2980 -20 3100 0
rect 2980 -100 3000 -20
rect 3080 -100 3100 -20
rect 2980 -120 3100 -100
rect 2980 -200 3000 -120
rect 3080 -200 3100 -120
rect 2980 -600 3100 -200
rect 4080 -60 4200 0
rect 4080 -140 4100 -60
rect 4180 -140 4200 -60
rect 4080 -180 4200 -140
rect 4080 -260 4100 -180
rect 4180 -260 4200 -180
rect 4080 -300 4200 -260
rect 4080 -380 4100 -300
rect 4180 -380 4200 -300
rect 4080 -600 4200 -380
rect 2980 -700 4200 -600
rect 4260 -60 4380 0
rect 4260 -140 4280 -60
rect 4360 -140 4380 -60
rect 4260 -180 4380 -140
rect 4260 -260 4280 -180
rect 4360 -260 4380 -180
rect 4260 -300 4380 -260
rect 4260 -380 4280 -300
rect 4360 -380 4380 -300
rect 960 -940 1620 -760
rect 4260 -780 4380 -380
rect 4800 -60 4920 0
rect 4800 -140 4820 -60
rect 4900 -140 4920 -60
rect 4800 -180 4920 -140
rect 4800 -260 4820 -180
rect 4900 -260 4920 -180
rect 4800 -300 4920 -260
rect 4800 -380 4820 -300
rect 4900 -380 4920 -300
rect 4800 -780 4920 -380
rect 4260 -940 4920 -780
rect 1100 -1960 1300 -940
rect 2560 -1080 2740 -1060
rect 2560 -1180 2600 -1080
rect 2700 -1180 2740 -1080
rect 2560 -1260 2740 -1180
rect 2560 -1360 2600 -1260
rect 2700 -1360 2740 -1260
rect 2560 -1400 2740 -1360
rect 3100 -1080 3280 -1060
rect 3100 -1180 3140 -1080
rect 3240 -1180 3280 -1080
rect 3100 -1260 3280 -1180
rect 3100 -1360 3140 -1260
rect 3240 -1360 3280 -1260
rect 3100 -1400 3280 -1360
rect 2580 -1800 2720 -1400
rect 2640 -1960 2720 -1800
rect 3140 -1800 3260 -1400
rect 3140 -1960 3240 -1800
rect 4580 -1960 4780 -940
rect 1100 -2020 2580 -1960
rect 1100 -2140 1960 -2020
rect 2080 -2140 2440 -2020
rect 2560 -2140 2580 -2020
rect 1100 -2180 2580 -2140
rect 2640 -2040 2800 -1960
rect 2640 -2160 2660 -2040
rect 2780 -2160 2800 -2040
rect 2640 -2180 2800 -2160
rect 3080 -2040 3240 -1960
rect 3080 -2160 3100 -2040
rect 3220 -2160 3240 -2040
rect 3080 -2180 3240 -2160
rect 3300 -2020 4780 -1960
rect 3300 -2140 3320 -2020
rect 3440 -2140 3800 -2020
rect 3920 -2140 4780 -2020
rect 3300 -2180 4780 -2140
use sky130_fd_pr__pfet_01v8_N6P669  XM5
timestamp 1769135993
transform 1 0 2940 0 1 -241
box -1940 -259 1940 293
use sky130_fd_pr__nfet_01v8_9PCEP7  XM8
timestamp 1769135993
transform 1 0 2916 0 1 -1273
box -516 -227 516 227
use sky130_fd_pr__nfet_01v8_VU2R7C  XM9
timestamp 1769135993
transform 1 0 2938 0 1 -2038
box -938 -162 938 162
<< labels >>
flabel metal1 800 -2500 1000 -2300 0 FreeSans 256 0 0 0 VSS
port 6 nsew
flabel metal1 760 160 960 360 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1600 -2800 1800 -2600 0 FreeSans 256 0 0 0 REF
port 1 nsew
flabel metal1 4100 -2800 4300 -2600 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal1 1100 -2800 1300 -2600 0 FreeSans 256 0 0 0 B2
port 5 nsew
flabel metal1 4600 -2800 4800 -2600 0 FreeSans 256 0 0 0 OUT
port 3 nsew
flabel metal1 2840 -2820 3040 -2620 0 FreeSans 256 0 0 0 B1
port 4 nsew
<< end >>
