magic
tech sky130A
magscale 1 2
timestamp 1770196220
<< error_p >>
rect -2559 1038 2559 1042
rect -2559 -970 -2529 1038
rect -2493 972 2493 976
rect -2493 -904 -2463 972
rect 2463 -904 2493 972
rect 2529 -970 2559 1038
<< nwell >>
rect -2529 -1004 2529 1038
<< mvpmos >>
rect -2435 -904 -2185 976
rect -2127 -904 -1877 976
rect -1819 -904 -1569 976
rect -1511 -904 -1261 976
rect -1203 -904 -953 976
rect -895 -904 -645 976
rect -587 -904 -337 976
rect -279 -904 -29 976
rect 29 -904 279 976
rect 337 -904 587 976
rect 645 -904 895 976
rect 953 -904 1203 976
rect 1261 -904 1511 976
rect 1569 -904 1819 976
rect 1877 -904 2127 976
rect 2185 -904 2435 976
<< mvpdiff >>
rect -2493 778 -2435 976
rect -2493 -706 -2481 778
rect -2447 -706 -2435 778
rect -2493 -904 -2435 -706
rect -2185 778 -2127 976
rect -2185 -706 -2173 778
rect -2139 -706 -2127 778
rect -2185 -904 -2127 -706
rect -1877 778 -1819 976
rect -1877 -706 -1865 778
rect -1831 -706 -1819 778
rect -1877 -904 -1819 -706
rect -1569 778 -1511 976
rect -1569 -706 -1557 778
rect -1523 -706 -1511 778
rect -1569 -904 -1511 -706
rect -1261 778 -1203 976
rect -1261 -706 -1249 778
rect -1215 -706 -1203 778
rect -1261 -904 -1203 -706
rect -953 778 -895 976
rect -953 -706 -941 778
rect -907 -706 -895 778
rect -953 -904 -895 -706
rect -645 778 -587 976
rect -645 -706 -633 778
rect -599 -706 -587 778
rect -645 -904 -587 -706
rect -337 778 -279 976
rect -337 -706 -325 778
rect -291 -706 -279 778
rect -337 -904 -279 -706
rect -29 778 29 976
rect -29 -706 -17 778
rect 17 -706 29 778
rect -29 -904 29 -706
rect 279 778 337 976
rect 279 -706 291 778
rect 325 -706 337 778
rect 279 -904 337 -706
rect 587 778 645 976
rect 587 -706 599 778
rect 633 -706 645 778
rect 587 -904 645 -706
rect 895 778 953 976
rect 895 -706 907 778
rect 941 -706 953 778
rect 895 -904 953 -706
rect 1203 778 1261 976
rect 1203 -706 1215 778
rect 1249 -706 1261 778
rect 1203 -904 1261 -706
rect 1511 778 1569 976
rect 1511 -706 1523 778
rect 1557 -706 1569 778
rect 1511 -904 1569 -706
rect 1819 778 1877 976
rect 1819 -706 1831 778
rect 1865 -706 1877 778
rect 1819 -904 1877 -706
rect 2127 778 2185 976
rect 2127 -706 2139 778
rect 2173 -706 2185 778
rect 2127 -904 2185 -706
rect 2435 778 2493 976
rect 2435 -706 2447 778
rect 2481 -706 2493 778
rect 2435 -904 2493 -706
<< mvpdiffc >>
rect -2481 -706 -2447 778
rect -2173 -706 -2139 778
rect -1865 -706 -1831 778
rect -1557 -706 -1523 778
rect -1249 -706 -1215 778
rect -941 -706 -907 778
rect -633 -706 -599 778
rect -325 -706 -291 778
rect -17 -706 17 778
rect 291 -706 325 778
rect 599 -706 633 778
rect 907 -706 941 778
rect 1215 -706 1249 778
rect 1523 -706 1557 778
rect 1831 -706 1865 778
rect 2139 -706 2173 778
rect 2447 -706 2481 778
<< poly >>
rect -2435 976 -2185 1002
rect -2127 976 -1877 1002
rect -1819 976 -1569 1002
rect -1511 976 -1261 1002
rect -1203 976 -953 1002
rect -895 976 -645 1002
rect -587 976 -337 1002
rect -279 976 -29 1002
rect 29 976 279 1002
rect 337 976 587 1002
rect 645 976 895 1002
rect 953 976 1203 1002
rect 1261 976 1511 1002
rect 1569 976 1819 1002
rect 1877 976 2127 1002
rect 2185 976 2435 1002
rect -2435 -951 -2185 -904
rect -2435 -985 -2419 -951
rect -2201 -985 -2185 -951
rect -2435 -1001 -2185 -985
rect -2127 -951 -1877 -904
rect -2127 -985 -2111 -951
rect -1893 -985 -1877 -951
rect -2127 -1001 -1877 -985
rect -1819 -951 -1569 -904
rect -1819 -985 -1803 -951
rect -1585 -985 -1569 -951
rect -1819 -1001 -1569 -985
rect -1511 -951 -1261 -904
rect -1511 -985 -1495 -951
rect -1277 -985 -1261 -951
rect -1511 -1001 -1261 -985
rect -1203 -951 -953 -904
rect -1203 -985 -1187 -951
rect -969 -985 -953 -951
rect -1203 -1001 -953 -985
rect -895 -951 -645 -904
rect -895 -985 -879 -951
rect -661 -985 -645 -951
rect -895 -1001 -645 -985
rect -587 -951 -337 -904
rect -587 -985 -571 -951
rect -353 -985 -337 -951
rect -587 -1001 -337 -985
rect -279 -951 -29 -904
rect -279 -985 -263 -951
rect -45 -985 -29 -951
rect -279 -1001 -29 -985
rect 29 -951 279 -904
rect 29 -985 45 -951
rect 263 -985 279 -951
rect 29 -1001 279 -985
rect 337 -951 587 -904
rect 337 -985 353 -951
rect 571 -985 587 -951
rect 337 -1001 587 -985
rect 645 -951 895 -904
rect 645 -985 661 -951
rect 879 -985 895 -951
rect 645 -1001 895 -985
rect 953 -951 1203 -904
rect 953 -985 969 -951
rect 1187 -985 1203 -951
rect 953 -1001 1203 -985
rect 1261 -951 1511 -904
rect 1261 -985 1277 -951
rect 1495 -985 1511 -951
rect 1261 -1001 1511 -985
rect 1569 -951 1819 -904
rect 1569 -985 1585 -951
rect 1803 -985 1819 -951
rect 1569 -1001 1819 -985
rect 1877 -951 2127 -904
rect 1877 -985 1893 -951
rect 2111 -985 2127 -951
rect 1877 -1001 2127 -985
rect 2185 -951 2435 -904
rect 2185 -985 2201 -951
rect 2419 -985 2435 -951
rect 2185 -1001 2435 -985
<< polycont >>
rect -2419 -985 -2201 -951
rect -2111 -985 -1893 -951
rect -1803 -985 -1585 -951
rect -1495 -985 -1277 -951
rect -1187 -985 -969 -951
rect -879 -985 -661 -951
rect -571 -985 -353 -951
rect -263 -985 -45 -951
rect 45 -985 263 -951
rect 353 -985 571 -951
rect 661 -985 879 -951
rect 969 -985 1187 -951
rect 1277 -985 1495 -951
rect 1585 -985 1803 -951
rect 1893 -985 2111 -951
rect 2201 -985 2419 -951
<< locali >>
rect -2481 778 -2447 794
rect -2481 -722 -2447 -706
rect -2173 778 -2139 794
rect -2173 -722 -2139 -706
rect -1865 778 -1831 794
rect -1865 -722 -1831 -706
rect -1557 778 -1523 794
rect -1557 -722 -1523 -706
rect -1249 778 -1215 794
rect -1249 -722 -1215 -706
rect -941 778 -907 794
rect -941 -722 -907 -706
rect -633 778 -599 794
rect -633 -722 -599 -706
rect -325 778 -291 794
rect -325 -722 -291 -706
rect -17 778 17 794
rect -17 -722 17 -706
rect 291 778 325 794
rect 291 -722 325 -706
rect 599 778 633 794
rect 599 -722 633 -706
rect 907 778 941 794
rect 907 -722 941 -706
rect 1215 778 1249 794
rect 1215 -722 1249 -706
rect 1523 778 1557 794
rect 1523 -722 1557 -706
rect 1831 778 1865 794
rect 1831 -722 1865 -706
rect 2139 778 2173 794
rect 2139 -722 2173 -706
rect 2447 778 2481 794
rect 2447 -722 2481 -706
rect -2435 -985 -2419 -951
rect -2201 -985 -2185 -951
rect -2127 -985 -2111 -951
rect -1893 -985 -1877 -951
rect -1819 -985 -1803 -951
rect -1585 -985 -1569 -951
rect -1511 -985 -1495 -951
rect -1277 -985 -1261 -951
rect -1203 -985 -1187 -951
rect -969 -985 -953 -951
rect -895 -985 -879 -951
rect -661 -985 -645 -951
rect -587 -985 -571 -951
rect -353 -985 -337 -951
rect -279 -985 -263 -951
rect -45 -985 -29 -951
rect 29 -985 45 -951
rect 263 -985 279 -951
rect 337 -985 353 -951
rect 571 -985 587 -951
rect 645 -985 661 -951
rect 879 -985 895 -951
rect 953 -985 969 -951
rect 1187 -985 1203 -951
rect 1261 -985 1277 -951
rect 1495 -985 1511 -951
rect 1569 -985 1585 -951
rect 1803 -985 1819 -951
rect 1877 -985 1893 -951
rect 2111 -985 2127 -951
rect 2185 -985 2201 -951
rect 2419 -985 2435 -951
<< viali >>
rect -2481 -706 -2447 778
rect -2173 -706 -2139 778
rect -1865 -706 -1831 778
rect -1557 -706 -1523 778
rect -1249 -706 -1215 778
rect -941 -706 -907 778
rect -633 -706 -599 778
rect -325 -706 -291 778
rect -17 -706 17 778
rect 291 -706 325 778
rect 599 -706 633 778
rect 907 -706 941 778
rect 1215 -706 1249 778
rect 1523 -706 1557 778
rect 1831 -706 1865 778
rect 2139 -706 2173 778
rect 2447 -706 2481 778
rect -2419 -985 -2201 -951
rect -2111 -985 -1893 -951
rect -1803 -985 -1585 -951
rect -1495 -985 -1277 -951
rect -1187 -985 -969 -951
rect -879 -985 -661 -951
rect -571 -985 -353 -951
rect -263 -985 -45 -951
rect 45 -985 263 -951
rect 353 -985 571 -951
rect 661 -985 879 -951
rect 969 -985 1187 -951
rect 1277 -985 1495 -951
rect 1585 -985 1803 -951
rect 1893 -985 2111 -951
rect 2201 -985 2419 -951
<< metal1 >>
rect -2487 778 -2441 790
rect -2487 -706 -2481 778
rect -2447 -706 -2441 778
rect -2487 -718 -2441 -706
rect -2179 778 -2133 790
rect -2179 -706 -2173 778
rect -2139 -706 -2133 778
rect -2179 -718 -2133 -706
rect -1871 778 -1825 790
rect -1871 -706 -1865 778
rect -1831 -706 -1825 778
rect -1871 -718 -1825 -706
rect -1563 778 -1517 790
rect -1563 -706 -1557 778
rect -1523 -706 -1517 778
rect -1563 -718 -1517 -706
rect -1255 778 -1209 790
rect -1255 -706 -1249 778
rect -1215 -706 -1209 778
rect -1255 -718 -1209 -706
rect -947 778 -901 790
rect -947 -706 -941 778
rect -907 -706 -901 778
rect -947 -718 -901 -706
rect -639 778 -593 790
rect -639 -706 -633 778
rect -599 -706 -593 778
rect -639 -718 -593 -706
rect -331 778 -285 790
rect -331 -706 -325 778
rect -291 -706 -285 778
rect -331 -718 -285 -706
rect -23 778 23 790
rect -23 -706 -17 778
rect 17 -706 23 778
rect -23 -718 23 -706
rect 285 778 331 790
rect 285 -706 291 778
rect 325 -706 331 778
rect 285 -718 331 -706
rect 593 778 639 790
rect 593 -706 599 778
rect 633 -706 639 778
rect 593 -718 639 -706
rect 901 778 947 790
rect 901 -706 907 778
rect 941 -706 947 778
rect 901 -718 947 -706
rect 1209 778 1255 790
rect 1209 -706 1215 778
rect 1249 -706 1255 778
rect 1209 -718 1255 -706
rect 1517 778 1563 790
rect 1517 -706 1523 778
rect 1557 -706 1563 778
rect 1517 -718 1563 -706
rect 1825 778 1871 790
rect 1825 -706 1831 778
rect 1865 -706 1871 778
rect 1825 -718 1871 -706
rect 2133 778 2179 790
rect 2133 -706 2139 778
rect 2173 -706 2179 778
rect 2133 -718 2179 -706
rect 2441 778 2487 790
rect 2441 -706 2447 778
rect 2481 -706 2487 778
rect 2441 -718 2487 -706
rect -2431 -951 -2189 -945
rect -2431 -985 -2419 -951
rect -2201 -985 -2189 -951
rect -2431 -991 -2189 -985
rect -2123 -951 -1881 -945
rect -2123 -985 -2111 -951
rect -1893 -985 -1881 -951
rect -2123 -991 -1881 -985
rect -1815 -951 -1573 -945
rect -1815 -985 -1803 -951
rect -1585 -985 -1573 -951
rect -1815 -991 -1573 -985
rect -1507 -951 -1265 -945
rect -1507 -985 -1495 -951
rect -1277 -985 -1265 -951
rect -1507 -991 -1265 -985
rect -1199 -951 -957 -945
rect -1199 -985 -1187 -951
rect -969 -985 -957 -951
rect -1199 -991 -957 -985
rect -891 -951 -649 -945
rect -891 -985 -879 -951
rect -661 -985 -649 -951
rect -891 -991 -649 -985
rect -583 -951 -341 -945
rect -583 -985 -571 -951
rect -353 -985 -341 -951
rect -583 -991 -341 -985
rect -275 -951 -33 -945
rect -275 -985 -263 -951
rect -45 -985 -33 -951
rect -275 -991 -33 -985
rect 33 -951 275 -945
rect 33 -985 45 -951
rect 263 -985 275 -951
rect 33 -991 275 -985
rect 341 -951 583 -945
rect 341 -985 353 -951
rect 571 -985 583 -951
rect 341 -991 583 -985
rect 649 -951 891 -945
rect 649 -985 661 -951
rect 879 -985 891 -951
rect 649 -991 891 -985
rect 957 -951 1199 -945
rect 957 -985 969 -951
rect 1187 -985 1199 -951
rect 957 -991 1199 -985
rect 1265 -951 1507 -945
rect 1265 -985 1277 -951
rect 1495 -985 1507 -951
rect 1265 -991 1507 -985
rect 1573 -951 1815 -945
rect 1573 -985 1585 -951
rect 1803 -985 1815 -951
rect 1573 -991 1815 -985
rect 1881 -951 2123 -945
rect 1881 -985 1893 -951
rect 2111 -985 2123 -951
rect 1881 -991 2123 -985
rect 2189 -951 2431 -945
rect 2189 -985 2201 -951
rect 2419 -985 2431 -951
rect 2189 -991 2431 -985
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9.4 l 1.25 m 1 nf 16 diffcov 80 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 80 viadrn 80 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
