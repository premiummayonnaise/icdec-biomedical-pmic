magic
tech sky130A
magscale 1 2
timestamp 1769573366
<< nwell >>
rect -2600 1120 11920 3680
<< pwell >>
rect -2600 -3640 11920 1120
<< locali >>
rect -2600 3900 11920 3940
rect -2600 3834 -2560 3900
rect -2602 3620 -2560 3834
rect -2260 3620 -2220 3900
rect -1920 3620 -1880 3900
rect -1580 3620 -1540 3900
rect -1240 3620 -1200 3900
rect -900 3620 -860 3900
rect -560 3620 -520 3900
rect -220 3620 -180 3900
rect 120 3620 160 3900
rect 460 3620 500 3900
rect 800 3620 840 3900
rect 1140 3620 1180 3900
rect 1480 3620 1520 3900
rect 1820 3620 1860 3900
rect 2160 3620 2200 3900
rect 2500 3620 2540 3900
rect 2840 3620 2880 3900
rect 3180 3620 3220 3900
rect 3520 3620 3560 3900
rect 3860 3620 3900 3900
rect 4200 3620 4240 3900
rect 4540 3620 4580 3900
rect 4880 3620 4920 3900
rect 5220 3620 5260 3900
rect 5560 3620 5600 3900
rect 5900 3620 5940 3900
rect 6240 3620 6280 3900
rect 6580 3620 6620 3900
rect 6920 3620 6960 3900
rect 7260 3620 7300 3900
rect 7600 3620 7640 3900
rect 7940 3620 7980 3900
rect 8280 3620 8320 3900
rect 8620 3620 8660 3900
rect 8960 3620 9000 3900
rect 9300 3620 9340 3900
rect 9640 3620 9680 3900
rect 9980 3620 10020 3900
rect 10320 3620 10360 3900
rect 10660 3620 10700 3900
rect 11000 3620 11040 3900
rect 11340 3620 11380 3900
rect 11680 3620 11920 3900
rect -2602 3564 11920 3620
rect -2600 3560 11920 3564
rect -920 1460 -760 3560
rect -300 1460 -140 3560
rect 320 1460 480 3560
rect 920 1460 1080 3560
rect 2100 3540 7240 3560
rect 2480 1560 2560 3540
rect 3100 1560 3180 3540
rect 3700 1560 3780 3540
rect 4320 1560 4400 3540
rect 4940 1560 5020 3540
rect 5560 1560 5640 3540
rect 6180 1560 6260 3540
rect 6780 1560 6860 3540
rect 8280 1440 8440 3560
rect 8900 1440 9060 3560
rect 9500 1440 9660 3560
rect 10120 1440 10280 3560
rect 3340 -220 3380 860
rect -2380 -240 3380 -220
rect -2380 -320 -2360 -240
rect -2280 -320 -2240 -240
rect -2020 -320 -1980 -240
rect -1900 -320 3380 -240
rect -2380 -360 3380 -320
rect -2380 -460 -2360 -360
rect -2280 -460 -2240 -360
rect -2020 -460 -1980 -360
rect -1900 -460 3380 -360
rect -2380 -500 3380 -460
rect 4700 -300 5800 -200
rect 5940 -220 5980 860
rect 5940 -240 11700 -220
rect 4700 -500 4800 -300
rect -2380 -580 -2360 -500
rect -2280 -580 -2240 -500
rect -2020 -580 -1980 -500
rect -1900 -580 3380 -500
rect -2380 -600 3380 -580
rect 3520 -520 4800 -500
rect 3520 -580 3540 -520
rect 3600 -580 3640 -520
rect 3700 -580 4800 -520
rect 3520 -600 4800 -580
rect 5940 -320 11220 -240
rect 11300 -320 11380 -240
rect 11520 -320 11600 -240
rect 11680 -320 11700 -240
rect 5940 -360 11700 -320
rect 5940 -460 11220 -360
rect 11300 -460 11380 -360
rect 11520 -460 11600 -360
rect 11680 -460 11700 -360
rect 5940 -500 11700 -460
rect 5940 -580 11220 -500
rect 11300 -580 11380 -500
rect 11520 -580 11600 -500
rect 11680 -580 11700 -500
rect 5940 -600 11700 -580
rect 3340 -1660 3380 -600
rect 5940 -1660 5980 -600
rect -520 -1900 9880 -1800
rect -300 -3560 -200 -1940
rect 300 -3560 400 -1940
rect 2120 -3460 2280 -1900
rect 3300 -1920 3500 -1900
rect 4540 -1910 4740 -1900
rect 2420 -3560 2580 -1940
rect 3040 -3560 3200 -1940
rect 3340 -3460 3500 -1920
rect 3640 -3560 3800 -1940
rect 4260 -3560 4420 -1940
rect 4580 -3460 4740 -1910
rect 5820 -1910 6040 -1900
rect 7000 -1910 7200 -1900
rect 4890 -3560 5050 -1940
rect 5500 -3560 5660 -1940
rect 5820 -3460 5980 -1910
rect 6140 -3560 6300 -1940
rect 6740 -3560 6900 -1940
rect 7040 -3460 7200 -1910
rect 8940 -3560 9040 -1960
rect 9540 -3560 9640 -1960
rect -2600 -3620 11920 -3560
rect -2600 -3900 -2560 -3620
rect -2260 -3900 -2220 -3620
rect -1920 -3900 -1880 -3620
rect -1580 -3900 -1540 -3620
rect -1240 -3900 -1200 -3620
rect -900 -3900 -860 -3620
rect -560 -3900 -520 -3620
rect -220 -3900 -180 -3620
rect 120 -3900 160 -3620
rect 460 -3900 500 -3620
rect 800 -3900 840 -3620
rect 1140 -3900 1180 -3620
rect 1480 -3900 1520 -3620
rect 1820 -3900 1860 -3620
rect 2160 -3900 2200 -3620
rect 2500 -3900 2540 -3620
rect 2840 -3900 2880 -3620
rect 3180 -3900 3220 -3620
rect 3520 -3900 3560 -3620
rect 3860 -3900 3900 -3620
rect 4200 -3900 4240 -3620
rect 4540 -3900 4580 -3620
rect 4880 -3900 4920 -3620
rect 5220 -3900 5260 -3620
rect 5560 -3900 5600 -3620
rect 5900 -3900 5940 -3620
rect 6240 -3900 6280 -3620
rect 6580 -3900 6620 -3620
rect 6920 -3900 6960 -3620
rect 7260 -3900 7300 -3620
rect 7600 -3900 7640 -3620
rect 7940 -3900 7980 -3620
rect 8280 -3900 8320 -3620
rect 8620 -3900 8660 -3620
rect 8960 -3900 9020 -3620
rect 9320 -3900 9360 -3620
rect 9660 -3900 9700 -3620
rect 10000 -3900 10040 -3620
rect 10340 -3900 10380 -3620
rect 10680 -3900 10720 -3620
rect 11020 -3900 11060 -3620
rect 11360 -3900 11400 -3620
rect 11700 -3900 11920 -3620
rect -2600 -3940 11920 -3900
<< viali >>
rect -2560 3620 -2260 3900
rect -2220 3620 -1920 3900
rect -1880 3620 -1580 3900
rect -1540 3620 -1240 3900
rect -1200 3620 -900 3900
rect -860 3620 -560 3900
rect -520 3620 -220 3900
rect -180 3620 120 3900
rect 160 3620 460 3900
rect 500 3620 800 3900
rect 840 3620 1140 3900
rect 1180 3620 1480 3900
rect 1520 3620 1820 3900
rect 1860 3620 2160 3900
rect 2200 3620 2500 3900
rect 2540 3620 2840 3900
rect 2880 3620 3180 3900
rect 3220 3620 3520 3900
rect 3560 3620 3860 3900
rect 3900 3620 4200 3900
rect 4240 3620 4540 3900
rect 4580 3620 4880 3900
rect 4920 3620 5220 3900
rect 5260 3620 5560 3900
rect 5600 3620 5900 3900
rect 5940 3620 6240 3900
rect 6280 3620 6580 3900
rect 6620 3620 6920 3900
rect 6960 3620 7260 3900
rect 7300 3620 7600 3900
rect 7640 3620 7940 3900
rect 7980 3620 8280 3900
rect 8320 3620 8620 3900
rect 8660 3620 8960 3900
rect 9000 3620 9300 3900
rect 9340 3620 9640 3900
rect 9680 3620 9980 3900
rect 10020 3620 10320 3900
rect 10360 3620 10660 3900
rect 10700 3620 11000 3900
rect 11040 3620 11340 3900
rect 11380 3620 11680 3900
rect -2360 -320 -2280 -240
rect -2240 -320 -2020 -240
rect -1980 -320 -1900 -240
rect -2360 -460 -2280 -360
rect -2240 -460 -2020 -360
rect -1980 -460 -1900 -360
rect -2360 -580 -2280 -500
rect -2240 -580 -2020 -500
rect -1980 -580 -1900 -500
rect 3540 -580 3600 -520
rect 3640 -580 3700 -520
rect 11220 -320 11300 -240
rect 11380 -320 11520 -240
rect 11600 -320 11680 -240
rect 11220 -460 11300 -360
rect 11380 -460 11520 -360
rect 11600 -460 11680 -360
rect 11220 -580 11300 -500
rect 11380 -580 11520 -500
rect 11600 -580 11680 -500
rect -2560 -3900 -2260 -3620
rect -2220 -3900 -1920 -3620
rect -1880 -3900 -1580 -3620
rect -1540 -3900 -1240 -3620
rect -1200 -3900 -900 -3620
rect -860 -3900 -560 -3620
rect -520 -3900 -220 -3620
rect -180 -3900 120 -3620
rect 160 -3900 460 -3620
rect 500 -3900 800 -3620
rect 840 -3900 1140 -3620
rect 1180 -3900 1480 -3620
rect 1520 -3900 1820 -3620
rect 1860 -3900 2160 -3620
rect 2200 -3900 2500 -3620
rect 2540 -3900 2840 -3620
rect 2880 -3900 3180 -3620
rect 3220 -3900 3520 -3620
rect 3560 -3900 3860 -3620
rect 3900 -3900 4200 -3620
rect 4240 -3900 4540 -3620
rect 4580 -3900 4880 -3620
rect 4920 -3900 5220 -3620
rect 5260 -3900 5560 -3620
rect 5600 -3900 5900 -3620
rect 5940 -3900 6240 -3620
rect 6280 -3900 6580 -3620
rect 6620 -3900 6920 -3620
rect 6960 -3900 7260 -3620
rect 7300 -3900 7600 -3620
rect 7640 -3900 7940 -3620
rect 7980 -3900 8280 -3620
rect 8320 -3900 8620 -3620
rect 8660 -3900 8960 -3620
rect 9020 -3900 9320 -3620
rect 9360 -3900 9660 -3620
rect 9700 -3900 10000 -3620
rect 10040 -3900 10340 -3620
rect 10380 -3900 10680 -3620
rect 10720 -3900 11020 -3620
rect 11060 -3900 11360 -3620
rect 11400 -3900 11700 -3620
<< metal1 >>
rect -2600 3900 11920 3940
rect -2600 3834 -2560 3900
rect -2602 3620 -2560 3834
rect -2260 3620 -2220 3900
rect -1920 3620 -1880 3900
rect -1580 3620 -1540 3900
rect -1240 3620 -1200 3900
rect -900 3620 -860 3900
rect -560 3620 -520 3900
rect -220 3620 -180 3900
rect 120 3620 160 3900
rect 460 3620 500 3900
rect 800 3620 840 3900
rect 1140 3620 1180 3900
rect 1480 3620 1520 3900
rect 1820 3620 1860 3900
rect 2160 3620 2200 3900
rect 2500 3620 2540 3900
rect 2840 3620 2880 3900
rect 3180 3620 3220 3900
rect 3520 3620 3560 3900
rect 3860 3620 3900 3900
rect 4200 3620 4240 3900
rect 4540 3620 4580 3900
rect 4880 3620 4920 3900
rect 5220 3620 5260 3900
rect 5560 3620 5600 3900
rect 5900 3620 5940 3900
rect 6240 3620 6280 3900
rect 6580 3620 6620 3900
rect 6920 3620 6960 3900
rect 7260 3620 7300 3900
rect 7600 3620 7640 3900
rect 7940 3620 7980 3900
rect 8280 3620 8320 3900
rect 8620 3620 8660 3900
rect 8960 3620 9000 3900
rect 9300 3620 9340 3900
rect 9640 3620 9680 3900
rect 9980 3620 10020 3900
rect 10320 3620 10360 3900
rect 10660 3620 10700 3900
rect 11000 3620 11040 3900
rect 11340 3620 11380 3900
rect 11680 3620 11920 3900
rect -2602 3564 11920 3620
rect -2600 3560 11920 3564
rect -2200 3420 -2060 3440
rect -2200 3360 -2160 3420
rect -2100 3360 -2060 3420
rect -2200 3280 -2060 3360
rect -2200 3220 -2160 3280
rect -2100 3220 -2060 3280
rect -2200 3200 -2060 3220
rect -1220 3120 -1080 3140
rect -1220 3060 -1180 3120
rect -1120 3060 -1080 3120
rect -1220 3020 -1080 3060
rect -1220 2960 -1180 3020
rect -1120 2960 -1080 3020
rect -1220 2920 -1080 2960
rect -1220 2860 -1180 2920
rect -1120 2860 -1080 2920
rect -1220 2840 -1080 2860
rect -600 3120 -460 3140
rect -600 3060 -560 3120
rect -500 3060 -460 3120
rect -600 3020 -460 3060
rect -600 2960 -560 3020
rect -500 2960 -460 3020
rect -600 2920 -460 2960
rect -600 2860 -560 2920
rect -500 2860 -460 2920
rect -600 2840 -460 2860
rect 0 3120 140 3140
rect 0 3060 40 3120
rect 100 3060 140 3120
rect 0 3020 140 3060
rect 0 2960 40 3020
rect 100 2960 140 3020
rect 0 2920 140 2960
rect 0 2860 40 2920
rect 100 2860 140 2920
rect 0 2840 140 2860
rect 620 3120 760 3140
rect 620 3060 660 3120
rect 720 3060 760 3120
rect 620 3020 760 3060
rect 620 2960 660 3020
rect 720 2960 760 3020
rect 620 2920 760 2960
rect 620 2860 660 2920
rect 720 2860 760 2920
rect 620 2840 760 2860
rect 1240 3120 1380 3140
rect 1240 3060 1280 3120
rect 1340 3060 1380 3120
rect 1240 3020 1380 3060
rect 1240 2960 1280 3020
rect 1340 2960 1380 3020
rect 1240 2920 1380 2960
rect 1240 2860 1280 2920
rect 1340 2860 1380 2920
rect 1240 2840 1380 2860
rect -2440 2780 -2300 2800
rect -2440 2720 -2400 2780
rect -2340 2720 -2300 2780
rect -2440 2680 -2300 2720
rect -2440 2620 -2400 2680
rect -2340 2620 -2300 2680
rect -2440 2580 -2300 2620
rect -2440 2520 -2400 2580
rect -2340 2520 -2300 2580
rect -2440 2500 -2300 2520
rect -1960 2780 -1820 2800
rect -1960 2720 -1920 2780
rect -1860 2720 -1820 2780
rect -1960 2680 -1820 2720
rect -1960 2620 -1920 2680
rect -1860 2620 -1820 2680
rect -1960 2580 -1820 2620
rect -1960 2520 -1920 2580
rect -1860 2520 -1820 2580
rect -1960 2500 -1820 2520
rect -2380 -240 -1880 2420
rect 2160 1520 2240 3460
rect 2760 2600 2880 2620
rect 2760 2520 2780 2600
rect 2860 2520 2880 2600
rect 2760 2380 2880 2520
rect 2760 2300 2780 2380
rect 2860 2300 2880 2380
rect 2760 2280 2880 2300
rect 3400 1520 3480 3460
rect 4000 2600 4120 2620
rect 4000 2520 4020 2600
rect 4100 2520 4120 2600
rect 4000 2380 4120 2520
rect 4000 2300 4020 2380
rect 4100 2300 4120 2380
rect 4000 2280 4120 2300
rect 4640 1520 4720 3460
rect 5220 2600 5340 2620
rect 5220 2520 5240 2600
rect 5320 2520 5340 2600
rect 5220 2380 5340 2520
rect 5220 2300 5240 2380
rect 5320 2300 5340 2380
rect 5220 2280 5340 2300
rect 5860 1520 5940 3460
rect 6460 2600 6580 2620
rect 6460 2520 6480 2600
rect 6560 2520 6580 2600
rect 6460 2380 6580 2520
rect 6460 2300 6480 2380
rect 6560 2300 6580 2380
rect 6460 2280 6580 2300
rect 7100 1520 7180 3460
rect 11380 3420 11520 3440
rect 11380 3360 11420 3420
rect 11480 3360 11520 3420
rect 11380 3280 11520 3360
rect 11380 3220 11420 3280
rect 11480 3220 11520 3280
rect 11380 3200 11520 3220
rect 7980 3120 8120 3140
rect 7980 3060 8020 3120
rect 8080 3060 8120 3120
rect 7980 3020 8120 3060
rect 7980 2960 8020 3020
rect 8080 2960 8120 3020
rect 7980 2920 8120 2960
rect 7980 2860 8020 2920
rect 8080 2860 8120 2920
rect 7980 2840 8120 2860
rect 8600 3120 8740 3140
rect 8600 3060 8640 3120
rect 8700 3060 8740 3120
rect 8600 3020 8740 3060
rect 8600 2960 8640 3020
rect 8700 2960 8740 3020
rect 8600 2920 8740 2960
rect 8600 2860 8640 2920
rect 8700 2860 8740 2920
rect 8600 2840 8740 2860
rect 9200 3120 9340 3140
rect 9200 3060 9240 3120
rect 9300 3060 9340 3120
rect 9200 3020 9340 3060
rect 9200 2960 9240 3020
rect 9300 2960 9340 3020
rect 9200 2920 9340 2960
rect 9200 2860 9240 2920
rect 9300 2860 9340 2920
rect 9200 2840 9340 2860
rect 9840 3120 9980 3140
rect 9840 3060 9880 3120
rect 9940 3060 9980 3120
rect 9840 3020 9980 3060
rect 9840 2960 9880 3020
rect 9940 2960 9980 3020
rect 9840 2920 9980 2960
rect 9840 2860 9880 2920
rect 9940 2860 9980 2920
rect 9840 2840 9980 2860
rect 10440 3120 10580 3140
rect 10440 3060 10480 3120
rect 10540 3060 10580 3120
rect 10440 3020 10580 3060
rect 10440 2960 10480 3020
rect 10540 2960 10580 3020
rect 10440 2920 10580 2960
rect 10440 2860 10480 2920
rect 10540 2860 10580 2920
rect 10440 2840 10580 2860
rect 11140 2760 11280 2780
rect 11140 2700 11180 2760
rect 11240 2700 11280 2760
rect 11140 2660 11280 2700
rect 11140 2600 11180 2660
rect 11240 2600 11280 2660
rect 11140 2560 11280 2600
rect 11140 2500 11180 2560
rect 11240 2500 11280 2560
rect 11140 2480 11280 2500
rect 11620 2760 11760 2780
rect 11620 2700 11660 2760
rect 11720 2700 11760 2760
rect 11620 2660 11760 2700
rect 11620 2600 11660 2660
rect 11720 2600 11760 2660
rect 11620 2560 11760 2600
rect 11620 2500 11660 2560
rect 11720 2500 11760 2560
rect 11620 2480 11760 2500
rect 2160 1440 7180 1520
rect -1120 1380 -880 1420
rect -1120 1280 -1100 1380
rect -900 1280 -880 1380
rect -1120 1240 -880 1280
rect -1120 1140 -1100 1240
rect -900 1140 -880 1240
rect -1120 1120 -880 1140
rect -820 1380 -580 1420
rect -820 1280 -800 1380
rect -600 1280 -580 1380
rect -820 1240 -580 1280
rect -820 1140 -800 1240
rect -600 1140 -580 1240
rect -820 1120 -580 1140
rect -500 1380 -260 1420
rect -500 1280 -480 1380
rect -280 1280 -260 1380
rect -500 1240 -260 1280
rect -500 1140 -480 1240
rect -280 1140 -260 1240
rect -500 1120 -260 1140
rect -200 1380 40 1420
rect -200 1280 -180 1380
rect 20 1280 40 1380
rect -200 1240 40 1280
rect -200 1140 -180 1240
rect 20 1140 40 1240
rect -200 1120 40 1140
rect 120 1380 360 1420
rect 120 1280 140 1380
rect 340 1280 360 1380
rect 120 1240 360 1280
rect 120 1140 140 1240
rect 340 1140 360 1240
rect 120 1120 360 1140
rect 420 1380 660 1420
rect 420 1280 440 1380
rect 640 1280 660 1380
rect 420 1240 660 1280
rect 420 1140 440 1240
rect 640 1140 660 1240
rect 420 1120 660 1140
rect 720 1380 960 1420
rect 720 1280 740 1380
rect 940 1280 960 1380
rect 720 1240 960 1280
rect 720 1140 740 1240
rect 940 1140 960 1240
rect 720 1120 960 1140
rect 1040 1380 1280 1420
rect 1040 1280 1060 1380
rect 1260 1280 1280 1380
rect 1040 1240 1280 1280
rect 1040 1140 1060 1240
rect 1260 1140 1280 1240
rect 1040 1120 1280 1140
rect -2380 -320 -2360 -240
rect -2280 -320 -2240 -240
rect -2020 -320 -1980 -240
rect -1900 -320 -1880 -240
rect -2380 -360 -1880 -320
rect -2380 -460 -2360 -360
rect -2280 -460 -2240 -360
rect -2020 -460 -1980 -360
rect -1900 -460 -1880 -360
rect -2380 -500 -1880 -460
rect -2380 -580 -2360 -500
rect -2280 -580 -2240 -500
rect -2020 -580 -1980 -500
rect -1900 -580 -1880 -500
rect -2380 -3560 -1880 -580
rect 2900 740 3300 1440
rect 3620 840 5700 980
rect 2900 680 2920 740
rect 3000 680 3200 740
rect 3280 680 3300 740
rect 2900 500 3300 680
rect 2900 440 2920 500
rect 3000 440 3200 500
rect 3280 440 3300 500
rect 2900 -1220 3300 440
rect 3440 740 3560 760
rect 3440 680 3460 740
rect 3540 680 3560 740
rect 3440 620 3560 680
rect 3440 560 3460 620
rect 3540 560 3560 620
rect 3440 500 3560 560
rect 3440 440 3460 500
rect 3540 440 3560 500
rect 3440 420 3560 440
rect 3620 -140 3700 840
rect 3760 740 3880 760
rect 3760 680 3780 740
rect 3860 680 3880 740
rect 3760 620 3880 680
rect 3760 560 3780 620
rect 3860 560 3880 620
rect 3760 500 3880 560
rect 3760 440 3780 500
rect 3860 440 3880 500
rect 3760 420 3880 440
rect 3920 -140 4000 840
rect 4080 740 4200 760
rect 4080 680 4100 740
rect 4180 680 4200 740
rect 4080 620 4200 680
rect 4080 560 4100 620
rect 4180 560 4200 620
rect 4080 500 4200 560
rect 4080 440 4100 500
rect 4180 440 4200 500
rect 4080 420 4200 440
rect 3500 -220 4332 -200
rect 3500 -280 4180 -220
rect 4240 -280 4260 -220
rect 4320 -280 4332 -220
rect 3500 -300 4332 -280
rect 3520 -520 3720 -500
rect 3520 -580 3540 -520
rect 3600 -580 3640 -520
rect 3700 -580 3720 -520
rect 3520 -600 3720 -580
rect 3440 -720 3560 -700
rect 3440 -780 3460 -720
rect 3540 -780 3560 -720
rect 3440 -840 3560 -780
rect 3440 -900 3460 -840
rect 3540 -900 3560 -840
rect 3440 -960 3560 -900
rect 3440 -1020 3460 -960
rect 3540 -1020 3560 -960
rect 3440 -1040 3560 -1020
rect 2900 -1280 2920 -1220
rect 3000 -1280 3200 -1220
rect 3280 -1280 3300 -1220
rect 2900 -1460 3300 -1280
rect 2900 -1520 2920 -1460
rect 3000 -1520 3200 -1460
rect 3280 -1520 3300 -1460
rect 2900 -1540 3300 -1520
rect 3640 -1640 3720 -660
rect 3760 -720 3880 -700
rect 3760 -780 3780 -720
rect 3860 -780 3880 -720
rect 3760 -840 3880 -780
rect 3760 -900 3780 -840
rect 3860 -900 3880 -840
rect 3760 -960 3880 -900
rect 3760 -1020 3780 -960
rect 3860 -1020 3880 -960
rect 3760 -1040 3880 -1020
rect 3920 -1640 4000 -660
rect 4060 -720 4180 -700
rect 4060 -780 4080 -720
rect 4160 -780 4180 -720
rect 4060 -840 4180 -780
rect 4060 -900 4080 -840
rect 4160 -900 4180 -840
rect 4060 -960 4180 -900
rect 4060 -1020 4080 -960
rect 4160 -1020 4180 -960
rect 4060 -1040 4180 -1020
rect 4580 -1640 4800 840
rect 5140 220 5260 240
rect 5140 160 5160 220
rect 5240 160 5260 220
rect 5140 100 5260 160
rect 5140 40 5160 100
rect 5240 40 5260 100
rect 5140 -20 5260 40
rect 5140 -80 5160 -20
rect 5240 -80 5260 -20
rect 5140 -100 5260 -80
rect 5340 -140 5420 840
rect 5460 220 5580 240
rect 5460 160 5480 220
rect 5560 160 5580 220
rect 5460 100 5580 160
rect 5460 40 5480 100
rect 5560 40 5580 100
rect 5460 -20 5580 40
rect 5460 -80 5480 -20
rect 5560 -80 5580 -20
rect 5460 -100 5580 -80
rect 5620 -140 5700 840
rect 6040 740 6440 1440
rect 8080 1360 8320 1400
rect 8080 1260 8100 1360
rect 8300 1260 8320 1360
rect 8080 1220 8320 1260
rect 8080 1120 8100 1220
rect 8300 1120 8320 1220
rect 8080 1100 8320 1120
rect 8380 1360 8620 1400
rect 8380 1260 8400 1360
rect 8600 1260 8620 1360
rect 8380 1220 8620 1260
rect 8380 1120 8400 1220
rect 8600 1120 8620 1220
rect 8380 1100 8620 1120
rect 8700 1360 8940 1400
rect 8700 1260 8720 1360
rect 8920 1260 8940 1360
rect 8700 1220 8940 1260
rect 8700 1120 8720 1220
rect 8920 1120 8940 1220
rect 8700 1100 8940 1120
rect 9000 1360 9240 1400
rect 9000 1260 9020 1360
rect 9220 1260 9240 1360
rect 9000 1220 9240 1260
rect 9000 1120 9020 1220
rect 9220 1120 9240 1220
rect 9000 1100 9240 1120
rect 9320 1360 9560 1400
rect 9320 1260 9340 1360
rect 9540 1260 9560 1360
rect 9320 1220 9560 1260
rect 9320 1120 9340 1220
rect 9540 1120 9560 1220
rect 9320 1100 9560 1120
rect 9620 1360 9860 1400
rect 9620 1260 9640 1360
rect 9840 1260 9860 1360
rect 9620 1220 9860 1260
rect 9620 1120 9640 1220
rect 9840 1120 9860 1220
rect 9620 1100 9860 1120
rect 9920 1360 10160 1400
rect 9920 1260 9940 1360
rect 10140 1260 10160 1360
rect 9920 1220 10160 1260
rect 9920 1120 9940 1220
rect 10140 1120 10160 1220
rect 9920 1100 10160 1120
rect 10240 1360 10480 1400
rect 10240 1260 10260 1360
rect 10460 1260 10480 1360
rect 10240 1220 10480 1260
rect 10240 1120 10260 1220
rect 10460 1120 10480 1220
rect 10240 1100 10480 1120
rect 6040 680 6060 740
rect 6140 680 6340 740
rect 6420 680 6440 740
rect 6040 500 6440 680
rect 6040 440 6060 500
rect 6140 440 6340 500
rect 6420 440 6440 500
rect 5780 220 5900 240
rect 5780 160 5800 220
rect 5880 160 5900 220
rect 5780 100 5900 160
rect 5780 40 5800 100
rect 5880 40 5900 100
rect 5780 -20 5900 40
rect 5780 -80 5800 -20
rect 5880 -80 5900 -20
rect 5780 -100 5900 -80
rect 5000 -520 5800 -500
rect 5000 -580 5020 -520
rect 5080 -580 5100 -520
rect 5160 -580 5660 -520
rect 5720 -580 5740 -520
rect 5000 -600 5800 -580
rect 5140 -1220 5260 -1200
rect 5140 -1280 5160 -1220
rect 5240 -1280 5260 -1220
rect 5140 -1340 5260 -1280
rect 5140 -1400 5160 -1340
rect 5240 -1400 5260 -1340
rect 5140 -1460 5260 -1400
rect 5140 -1520 5160 -1460
rect 5240 -1520 5260 -1460
rect 5140 -1540 5260 -1520
rect 5340 -1640 5420 -660
rect 5460 -1220 5580 -1200
rect 5460 -1280 5480 -1220
rect 5560 -1280 5580 -1220
rect 5460 -1340 5580 -1280
rect 5460 -1400 5480 -1340
rect 5560 -1400 5580 -1340
rect 5460 -1460 5580 -1400
rect 5460 -1520 5480 -1460
rect 5560 -1520 5580 -1460
rect 5460 -1540 5580 -1520
rect 5620 -1640 5700 -660
rect 5760 -1220 5880 -1200
rect 5760 -1280 5780 -1220
rect 5860 -1280 5880 -1220
rect 5760 -1340 5880 -1280
rect 5760 -1400 5780 -1340
rect 5860 -1400 5880 -1340
rect 5760 -1460 5880 -1400
rect 5760 -1520 5780 -1460
rect 5860 -1520 5880 -1460
rect 5760 -1540 5880 -1520
rect 6040 -1220 6440 440
rect 6040 -1280 6060 -1220
rect 6140 -1280 6340 -1220
rect 6420 -1280 6440 -1220
rect 6040 -1460 6440 -1280
rect 6040 -1520 6060 -1460
rect 6140 -1520 6340 -1460
rect 6420 -1520 6440 -1460
rect 6040 -1540 6440 -1520
rect 11200 -240 11700 2400
rect 11200 -320 11220 -240
rect 11300 -320 11380 -240
rect 11520 -320 11600 -240
rect 11680 -320 11700 -240
rect 11200 -360 11700 -320
rect 11200 -460 11220 -360
rect 11300 -460 11380 -360
rect 11520 -460 11600 -360
rect 11680 -460 11700 -360
rect 11200 -500 11700 -460
rect 11200 -580 11220 -500
rect 11300 -580 11380 -500
rect 11520 -580 11600 -500
rect 11680 -580 11700 -500
rect 2740 -1780 6600 -1640
rect -640 -2600 -500 -2580
rect -640 -2660 -600 -2600
rect -540 -2660 -500 -2600
rect -640 -2700 -500 -2660
rect -640 -2760 -600 -2700
rect -540 -2760 -500 -2700
rect -640 -2800 -500 -2760
rect -640 -2860 -600 -2800
rect -540 -2860 -500 -2800
rect -640 -2880 -500 -2860
rect -20 -2600 120 -2580
rect -20 -2660 20 -2600
rect 80 -2660 120 -2600
rect -20 -2700 120 -2660
rect -20 -2760 20 -2700
rect 80 -2760 120 -2700
rect -20 -2800 120 -2760
rect -20 -2860 20 -2800
rect 80 -2860 120 -2800
rect -20 -2880 120 -2860
rect 600 -2600 740 -2580
rect 600 -2660 640 -2600
rect 700 -2660 740 -2600
rect 600 -2700 740 -2660
rect 600 -2760 640 -2700
rect 700 -2760 740 -2700
rect 600 -2800 740 -2760
rect 600 -2860 640 -2800
rect 700 -2860 740 -2800
rect 600 -2880 740 -2860
rect 2740 -3440 2900 -1780
rect 3960 -3440 4120 -1780
rect 4560 -2040 4760 -1960
rect 4560 -2120 4620 -2040
rect 4700 -2120 4760 -2040
rect 4560 -2160 4760 -2120
rect 4560 -2240 4620 -2160
rect 4700 -2240 4760 -2160
rect 4560 -2280 4760 -2240
rect 4560 -2360 4620 -2280
rect 4700 -2360 4760 -2280
rect 4560 -2400 4760 -2360
rect 4560 -2480 4620 -2400
rect 4700 -2480 4760 -2400
rect 4560 -2520 4760 -2480
rect 4560 -2600 4620 -2520
rect 4700 -2600 4760 -2520
rect 4560 -2640 4760 -2600
rect 4560 -2720 4620 -2640
rect 4700 -2720 4760 -2640
rect 4560 -2760 4760 -2720
rect 4560 -2840 4620 -2760
rect 4700 -2840 4760 -2760
rect 4560 -2880 4760 -2840
rect 4560 -2960 4620 -2880
rect 4700 -2960 4760 -2880
rect 4560 -3000 4760 -2960
rect 4560 -3080 4620 -3000
rect 4700 -3080 4760 -3000
rect 4560 -3120 4760 -3080
rect 4560 -3200 4620 -3120
rect 4700 -3200 4760 -3120
rect 4560 -3240 4760 -3200
rect 4560 -3320 4620 -3240
rect 4700 -3320 4760 -3240
rect 4560 -3360 4760 -3320
rect 4560 -3440 4620 -3360
rect 4700 -3440 4760 -3360
rect 5200 -3440 5360 -1780
rect 6440 -3440 6600 -1780
rect 8600 -2580 8740 -2560
rect 8600 -2640 8640 -2580
rect 8700 -2640 8740 -2580
rect 8600 -2680 8740 -2640
rect 8600 -2740 8640 -2680
rect 8700 -2740 8740 -2680
rect 8600 -2780 8740 -2740
rect 8600 -2840 8640 -2780
rect 8700 -2840 8740 -2780
rect 8600 -2860 8740 -2840
rect 9220 -2580 9360 -2560
rect 9220 -2640 9260 -2580
rect 9320 -2640 9360 -2580
rect 9220 -2680 9360 -2640
rect 9220 -2740 9260 -2680
rect 9320 -2740 9360 -2680
rect 9220 -2780 9360 -2740
rect 9220 -2840 9260 -2780
rect 9320 -2840 9360 -2780
rect 9220 -2860 9360 -2840
rect 9840 -2580 9980 -2560
rect 9840 -2640 9880 -2580
rect 9940 -2640 9980 -2580
rect 9840 -2680 9980 -2640
rect 9840 -2740 9880 -2680
rect 9940 -2740 9980 -2680
rect 9840 -2780 9980 -2740
rect 9840 -2840 9880 -2780
rect 9940 -2840 9980 -2780
rect 9840 -2860 9980 -2840
rect 4560 -3460 4760 -3440
rect 11200 -3560 11700 -580
rect -2600 -3620 11920 -3560
rect -2600 -3900 -2560 -3620
rect -2260 -3900 -2220 -3620
rect -1920 -3900 -1880 -3620
rect -1580 -3900 -1540 -3620
rect -1240 -3900 -1200 -3620
rect -900 -3900 -860 -3620
rect -560 -3900 -520 -3620
rect -220 -3900 -180 -3620
rect 120 -3900 160 -3620
rect 460 -3900 500 -3620
rect 800 -3900 840 -3620
rect 1140 -3900 1180 -3620
rect 1480 -3900 1520 -3620
rect 1820 -3900 1860 -3620
rect 2160 -3900 2200 -3620
rect 2500 -3900 2540 -3620
rect 2840 -3900 2880 -3620
rect 3180 -3900 3220 -3620
rect 3520 -3900 3560 -3620
rect 3860 -3900 3900 -3620
rect 4200 -3900 4240 -3620
rect 4540 -3900 4580 -3620
rect 4880 -3900 4920 -3620
rect 5220 -3900 5260 -3620
rect 5560 -3900 5600 -3620
rect 5900 -3900 5940 -3620
rect 6240 -3900 6280 -3620
rect 6580 -3900 6620 -3620
rect 6920 -3900 6960 -3620
rect 7260 -3900 7300 -3620
rect 7600 -3900 7640 -3620
rect 7940 -3900 7980 -3620
rect 8280 -3900 8320 -3620
rect 8620 -3900 8660 -3620
rect 8960 -3900 9020 -3620
rect 9320 -3900 9360 -3620
rect 9660 -3900 9700 -3620
rect 10000 -3900 10040 -3620
rect 10340 -3900 10380 -3620
rect 10680 -3900 10720 -3620
rect 11020 -3900 11060 -3620
rect 11360 -3900 11400 -3620
rect 11700 -3900 11920 -3620
rect -2600 -3940 11920 -3900
rect 1200 -4160 1400 -4140
rect 8000 -4160 8200 -4140
rect 1200 -4220 1220 -4160
rect 1280 -4220 1320 -4160
rect 1380 -4220 1400 -4160
rect 1200 -4260 1400 -4220
rect 1200 -4320 1220 -4260
rect 1280 -4320 1320 -4260
rect 1380 -4320 1400 -4260
rect 1200 -4340 1400 -4320
rect 4560 -4180 4760 -4160
rect 4560 -4240 4580 -4180
rect 4640 -4240 4680 -4180
rect 4740 -4240 4760 -4180
rect 4560 -4280 4760 -4240
rect 4560 -4340 4580 -4280
rect 4640 -4340 4680 -4280
rect 4740 -4340 4760 -4280
rect 8000 -4220 8020 -4160
rect 8080 -4220 8120 -4160
rect 8180 -4220 8200 -4160
rect 8000 -4260 8200 -4220
rect 8000 -4320 8020 -4260
rect 8080 -4320 8120 -4260
rect 8180 -4320 8200 -4260
rect 8000 -4340 8200 -4320
rect 4560 -4360 4760 -4340
rect 4540 -5640 4740 -5620
rect 4540 -5700 4560 -5640
rect 4620 -5700 4660 -5640
rect 4720 -5700 4740 -5640
rect 4540 -5740 4740 -5700
rect 4540 -5800 4560 -5740
rect 4620 -5800 4660 -5740
rect 4720 -5800 4740 -5740
rect 4540 -5820 4740 -5800
<< via1 >>
rect -2160 3360 -2100 3420
rect -2160 3220 -2100 3280
rect -1180 3060 -1120 3120
rect -1180 2960 -1120 3020
rect -1180 2860 -1120 2920
rect -560 3060 -500 3120
rect -560 2960 -500 3020
rect -560 2860 -500 2920
rect 40 3060 100 3120
rect 40 2960 100 3020
rect 40 2860 100 2920
rect 660 3060 720 3120
rect 660 2960 720 3020
rect 660 2860 720 2920
rect 1280 3060 1340 3120
rect 1280 2960 1340 3020
rect 1280 2860 1340 2920
rect -2400 2720 -2340 2780
rect -2400 2620 -2340 2680
rect -2400 2520 -2340 2580
rect -1920 2720 -1860 2780
rect -1920 2620 -1860 2680
rect -1920 2520 -1860 2580
rect 2780 2520 2860 2600
rect 2780 2300 2860 2380
rect 4020 2520 4100 2600
rect 4020 2300 4100 2380
rect 5240 2520 5320 2600
rect 5240 2300 5320 2380
rect 6480 2520 6560 2600
rect 6480 2300 6560 2380
rect 11420 3360 11480 3420
rect 11420 3220 11480 3280
rect 8020 3060 8080 3120
rect 8020 2960 8080 3020
rect 8020 2860 8080 2920
rect 8640 3060 8700 3120
rect 8640 2960 8700 3020
rect 8640 2860 8700 2920
rect 9240 3060 9300 3120
rect 9240 2960 9300 3020
rect 9240 2860 9300 2920
rect 9880 3060 9940 3120
rect 9880 2960 9940 3020
rect 9880 2860 9940 2920
rect 10480 3060 10540 3120
rect 10480 2960 10540 3020
rect 10480 2860 10540 2920
rect 11180 2700 11240 2760
rect 11180 2600 11240 2660
rect 11180 2500 11240 2560
rect 11660 2700 11720 2760
rect 11660 2600 11720 2660
rect 11660 2500 11720 2560
rect -1100 1280 -900 1380
rect -1100 1140 -900 1240
rect -800 1280 -600 1380
rect -800 1140 -600 1240
rect -480 1280 -280 1380
rect -480 1140 -280 1240
rect -180 1280 20 1380
rect -180 1140 20 1240
rect 140 1280 340 1380
rect 140 1140 340 1240
rect 440 1280 640 1380
rect 440 1140 640 1240
rect 740 1280 940 1380
rect 740 1140 940 1240
rect 1060 1280 1260 1380
rect 1060 1140 1260 1240
rect 2920 680 3000 740
rect 3200 680 3280 740
rect 2920 440 3000 500
rect 3200 440 3280 500
rect 3460 680 3540 740
rect 3460 560 3540 620
rect 3460 440 3540 500
rect 3780 680 3860 740
rect 3780 560 3860 620
rect 3780 440 3860 500
rect 4100 680 4180 740
rect 4100 560 4180 620
rect 4100 440 4180 500
rect 4180 -280 4240 -220
rect 4260 -280 4320 -220
rect 3540 -580 3600 -520
rect 3640 -580 3700 -520
rect 3460 -780 3540 -720
rect 3460 -900 3540 -840
rect 3460 -1020 3540 -960
rect 2920 -1280 3000 -1220
rect 3200 -1280 3280 -1220
rect 2920 -1520 3000 -1460
rect 3200 -1520 3280 -1460
rect 3780 -780 3860 -720
rect 3780 -900 3860 -840
rect 3780 -1020 3860 -960
rect 4080 -780 4160 -720
rect 4080 -900 4160 -840
rect 4080 -1020 4160 -960
rect 5160 160 5240 220
rect 5160 40 5240 100
rect 5160 -80 5240 -20
rect 5480 160 5560 220
rect 5480 40 5560 100
rect 5480 -80 5560 -20
rect 8100 1260 8300 1360
rect 8100 1120 8300 1220
rect 8400 1260 8600 1360
rect 8400 1120 8600 1220
rect 8720 1260 8920 1360
rect 8720 1120 8920 1220
rect 9020 1260 9220 1360
rect 9020 1120 9220 1220
rect 9340 1260 9540 1360
rect 9340 1120 9540 1220
rect 9640 1260 9840 1360
rect 9640 1120 9840 1220
rect 9940 1260 10140 1360
rect 9940 1120 10140 1220
rect 10260 1260 10460 1360
rect 10260 1120 10460 1220
rect 6060 680 6140 740
rect 6340 680 6420 740
rect 6060 440 6140 500
rect 6340 440 6420 500
rect 5800 160 5880 220
rect 5800 40 5880 100
rect 5800 -80 5880 -20
rect 5020 -580 5080 -520
rect 5100 -580 5160 -520
rect 5660 -580 5720 -520
rect 5740 -580 5800 -520
rect 5160 -1280 5240 -1220
rect 5160 -1400 5240 -1340
rect 5160 -1520 5240 -1460
rect 5480 -1280 5560 -1220
rect 5480 -1400 5560 -1340
rect 5480 -1520 5560 -1460
rect 5780 -1280 5860 -1220
rect 5780 -1400 5860 -1340
rect 5780 -1520 5860 -1460
rect 6060 -1280 6140 -1220
rect 6340 -1280 6420 -1220
rect 6060 -1520 6140 -1460
rect 6340 -1520 6420 -1460
rect -600 -2660 -540 -2600
rect -600 -2760 -540 -2700
rect -600 -2860 -540 -2800
rect 20 -2660 80 -2600
rect 20 -2760 80 -2700
rect 20 -2860 80 -2800
rect 640 -2660 700 -2600
rect 640 -2760 700 -2700
rect 640 -2860 700 -2800
rect 4620 -2120 4700 -2040
rect 4620 -2240 4700 -2160
rect 4620 -2360 4700 -2280
rect 4620 -2480 4700 -2400
rect 4620 -2600 4700 -2520
rect 4620 -2720 4700 -2640
rect 4620 -2840 4700 -2760
rect 4620 -2960 4700 -2880
rect 4620 -3080 4700 -3000
rect 4620 -3200 4700 -3120
rect 4620 -3320 4700 -3240
rect 4620 -3440 4700 -3360
rect 8640 -2640 8700 -2580
rect 8640 -2740 8700 -2680
rect 8640 -2840 8700 -2780
rect 9260 -2640 9320 -2580
rect 9260 -2740 9320 -2680
rect 9260 -2840 9320 -2780
rect 9880 -2640 9940 -2580
rect 9880 -2740 9940 -2680
rect 9880 -2840 9940 -2780
rect 1220 -4220 1280 -4160
rect 1320 -4220 1380 -4160
rect 1220 -4320 1280 -4260
rect 1320 -4320 1380 -4260
rect 4580 -4240 4640 -4180
rect 4680 -4240 4740 -4180
rect 4580 -4340 4640 -4280
rect 4680 -4340 4740 -4280
rect 8020 -4220 8080 -4160
rect 8120 -4220 8180 -4160
rect 8020 -4320 8080 -4260
rect 8120 -4320 8180 -4260
rect 4560 -5700 4620 -5640
rect 4660 -5700 4720 -5640
rect 4560 -5800 4620 -5740
rect 4660 -5800 4720 -5740
<< metal2 >>
rect -2400 3420 -1260 3440
rect -2400 3360 -2160 3420
rect -2100 3360 -1640 3420
rect -1580 3360 -1540 3420
rect -1480 3360 -1440 3420
rect -1380 3360 -1340 3420
rect -1280 3360 -1260 3420
rect -2400 3280 -1260 3360
rect -2400 3220 -2160 3280
rect -2100 3220 -1640 3280
rect -1580 3220 -1540 3280
rect -1480 3220 -1440 3280
rect -1380 3220 -1340 3280
rect -1280 3220 -1260 3280
rect -2400 3200 -1260 3220
rect 10620 3420 11760 3440
rect 10620 3360 10640 3420
rect 10700 3360 10740 3420
rect 10800 3360 10840 3420
rect 10900 3360 10940 3420
rect 11000 3360 11420 3420
rect 11480 3360 11760 3420
rect 10620 3280 11760 3360
rect 10620 3220 10640 3280
rect 10700 3220 10740 3280
rect 10800 3220 10840 3280
rect 10900 3220 10940 3280
rect 11000 3220 11420 3280
rect 11480 3220 11760 3280
rect 10620 3200 11760 3220
rect -3160 3120 1460 3140
rect -3160 3060 -1180 3120
rect -1120 3060 -560 3120
rect -500 3060 40 3120
rect 100 3060 660 3120
rect 720 3060 1280 3120
rect 1340 3060 1460 3120
rect -3160 3020 1460 3060
rect -3160 2960 -1180 3020
rect -1120 2960 -560 3020
rect -500 2960 40 3020
rect 100 2960 660 3020
rect 720 2960 1280 3020
rect 1340 2960 1460 3020
rect -3160 2920 1460 2960
rect -3160 2860 -1180 2920
rect -1120 2860 -560 2920
rect -500 2860 40 2920
rect 100 2860 660 2920
rect 720 2860 1280 2920
rect 1340 2860 1460 2920
rect -3160 2840 1460 2860
rect 7860 3120 12480 3140
rect 7860 3060 8020 3120
rect 8080 3060 8640 3120
rect 8700 3060 9240 3120
rect 9300 3060 9880 3120
rect 9940 3060 10480 3120
rect 10540 3060 12480 3120
rect 7860 3020 12480 3060
rect 7860 2960 8020 3020
rect 8080 2960 8640 3020
rect 8700 2960 9240 3020
rect 9300 2960 9880 3020
rect 9940 2960 10480 3020
rect 10540 2960 12480 3020
rect 7860 2920 12480 2960
rect 7860 2860 8020 2920
rect 8080 2860 8640 2920
rect 8700 2860 9240 2920
rect 9300 2860 9880 2920
rect 9940 2860 10480 2920
rect 10540 2860 12480 2920
rect 7860 2840 12480 2860
rect -3160 2800 -2860 2840
rect -3160 2780 -1260 2800
rect 12180 2780 12480 2840
rect -3160 2720 -2400 2780
rect -2340 2720 -1920 2780
rect -1860 2720 -1260 2780
rect -3160 2680 -1260 2720
rect -3160 2620 -2400 2680
rect -2340 2620 -1920 2680
rect -1860 2620 -1260 2680
rect 10620 2760 12480 2780
rect 10620 2700 11180 2760
rect 11240 2700 11660 2760
rect 11720 2700 12480 2760
rect 10620 2660 12480 2700
rect -3160 2580 -1260 2620
rect -3160 2520 -2400 2580
rect -2340 2520 -1920 2580
rect -1860 2520 -1260 2580
rect -3160 2500 -1260 2520
rect 1600 2600 7800 2620
rect 1600 2520 2780 2600
rect 2860 2520 4020 2600
rect 4100 2520 5240 2600
rect 5320 2520 6480 2600
rect 6560 2520 7420 2600
rect 7500 2520 7560 2600
rect 7640 2520 7700 2600
rect 7780 2520 7800 2600
rect -3160 -2580 -2860 2500
rect 1600 2380 7800 2520
rect 10620 2600 11180 2660
rect 11240 2600 11660 2660
rect 11720 2600 12480 2660
rect 10620 2560 12480 2600
rect 10620 2500 11180 2560
rect 11240 2500 11660 2560
rect 11720 2500 12480 2560
rect 10620 2480 12480 2500
rect 1600 2300 2780 2380
rect 2860 2300 4020 2380
rect 4100 2300 5240 2380
rect 5320 2300 6480 2380
rect 6560 2300 7420 2380
rect 7500 2300 7560 2380
rect 7640 2300 7700 2380
rect 7780 2300 7800 2380
rect 1600 2280 7800 2300
rect -1200 1400 2000 1420
rect -1200 1380 1620 1400
rect -1200 1280 -1100 1380
rect -900 1280 -800 1380
rect -600 1280 -480 1380
rect -280 1280 -180 1380
rect 20 1280 140 1380
rect 340 1280 440 1380
rect 640 1280 740 1380
rect 940 1280 1060 1380
rect 1260 1320 1620 1380
rect 1700 1320 1760 1400
rect 1840 1320 1900 1400
rect 1980 1320 2000 1400
rect 1260 1280 2000 1320
rect -1200 1240 2000 1280
rect -1200 1140 -1100 1240
rect -900 1140 -800 1240
rect -600 1140 -480 1240
rect -280 1140 -180 1240
rect 20 1140 140 1240
rect 340 1140 440 1240
rect 640 1140 740 1240
rect 940 1140 1060 1240
rect 1260 1220 2000 1240
rect 1260 1140 1620 1220
rect 1700 1140 1760 1220
rect 1840 1140 1900 1220
rect 1980 1140 2000 1220
rect -1200 1120 2000 1140
rect 7400 1380 10540 1400
rect 7400 1300 7420 1380
rect 7500 1300 7560 1380
rect 7640 1300 7700 1380
rect 7780 1360 10540 1380
rect 7780 1300 8100 1360
rect 7400 1260 8100 1300
rect 8300 1260 8400 1360
rect 8600 1260 8720 1360
rect 8920 1260 9020 1360
rect 9220 1260 9340 1360
rect 9540 1260 9640 1360
rect 9840 1260 9940 1360
rect 10140 1260 10260 1360
rect 10460 1260 10540 1360
rect 7400 1220 10540 1260
rect 7400 1200 8100 1220
rect 7400 1120 7420 1200
rect 7500 1120 7560 1200
rect 7640 1120 7700 1200
rect 7780 1120 8100 1200
rect 8300 1120 8400 1220
rect 8600 1120 8720 1220
rect 8920 1120 9020 1220
rect 9220 1120 9340 1220
rect 9540 1120 9640 1220
rect 9840 1120 9940 1220
rect 10140 1120 10260 1220
rect 10460 1120 10540 1220
rect 7400 1100 10540 1120
rect 1600 740 7800 760
rect 1600 680 2920 740
rect 3000 680 3200 740
rect 3280 680 3460 740
rect 3540 680 3780 740
rect 3860 680 4100 740
rect 4180 680 6060 740
rect 6140 680 6340 740
rect 6420 680 7800 740
rect 1600 620 7800 680
rect 1600 560 3460 620
rect 3540 560 3780 620
rect 3860 560 4100 620
rect 4180 560 7800 620
rect 1600 500 7800 560
rect 1600 440 2920 500
rect 3000 440 3200 500
rect 3280 440 3460 500
rect 3540 440 3780 500
rect 3860 440 4100 500
rect 4180 440 6060 500
rect 6140 440 6340 500
rect 6420 440 7800 500
rect 1600 420 7800 440
rect 1600 220 7800 240
rect 1600 140 1620 220
rect 1700 140 1740 220
rect 1860 140 1900 220
rect 1980 160 5160 220
rect 5240 160 5480 220
rect 5560 160 5800 220
rect 5880 160 7420 220
rect 1980 140 7420 160
rect 7500 140 7540 220
rect 7660 140 7700 220
rect 7780 140 7800 220
rect 1600 100 7800 140
rect 1600 40 5160 100
rect 5240 40 5480 100
rect 5560 40 5800 100
rect 5880 40 7800 100
rect 1600 0 7800 40
rect 1600 -80 1620 0
rect 1700 -80 1740 0
rect 1860 -80 1900 0
rect 1980 -20 7420 0
rect 1980 -80 5160 -20
rect 5240 -80 5480 -20
rect 5560 -80 5800 -20
rect 5880 -80 7420 -20
rect 7500 -80 7540 0
rect 7660 -80 7700 0
rect 7780 -80 7800 0
rect 1600 -100 7800 -80
rect 4154 -200 4700 -198
rect 1120 -220 3300 -200
rect 1120 -300 1140 -220
rect 1220 -300 1260 -220
rect 1360 -300 1400 -220
rect 1480 -300 3300 -220
rect 4154 -220 4702 -200
rect 4154 -280 4180 -220
rect 4240 -280 4260 -220
rect 4320 -280 4702 -220
rect 4154 -300 4702 -280
rect 1120 -360 3300 -300
rect 1120 -440 1140 -360
rect 1220 -440 1260 -360
rect 1360 -440 1400 -360
rect 1480 -440 3300 -360
rect 1120 -500 3300 -440
rect 4602 -500 4702 -300
rect 6040 -220 8280 -200
rect 6040 -300 7920 -220
rect 8000 -300 8040 -220
rect 8140 -300 8180 -220
rect 8260 -300 8280 -220
rect 6040 -360 8280 -300
rect 6040 -440 7920 -360
rect 8000 -440 8040 -360
rect 8140 -440 8180 -360
rect 8260 -440 8280 -360
rect 6040 -500 8280 -440
rect 1120 -580 1140 -500
rect 1220 -580 1260 -500
rect 1360 -580 1400 -500
rect 1480 -520 3720 -500
rect 1480 -580 3540 -520
rect 3600 -580 3640 -520
rect 3700 -580 3720 -520
rect 1120 -600 3720 -580
rect 4602 -520 5170 -500
rect 4602 -580 5020 -520
rect 5080 -580 5100 -520
rect 5160 -580 5170 -520
rect 4602 -600 5170 -580
rect 5640 -520 7920 -500
rect 5640 -580 5660 -520
rect 5720 -580 5740 -520
rect 5800 -580 7920 -520
rect 8000 -580 8040 -500
rect 8140 -580 8180 -500
rect 8260 -580 8280 -500
rect 5640 -600 8280 -580
rect 1600 -720 7800 -700
rect 1600 -800 1620 -720
rect 1700 -800 1740 -720
rect 1860 -800 1900 -720
rect 1980 -780 3460 -720
rect 3540 -780 3780 -720
rect 3860 -780 4080 -720
rect 4160 -780 7420 -720
rect 1980 -800 7420 -780
rect 7500 -800 7540 -720
rect 7660 -800 7700 -720
rect 7780 -800 7800 -720
rect 1600 -840 7800 -800
rect 1600 -900 3460 -840
rect 3540 -900 3780 -840
rect 3860 -900 4080 -840
rect 4160 -900 7800 -840
rect 1600 -920 7800 -900
rect 1600 -1000 1620 -920
rect 1700 -1000 1740 -920
rect 1860 -1000 1900 -920
rect 1980 -940 7800 -920
rect 1980 -960 7420 -940
rect 1980 -1000 3460 -960
rect 1600 -1020 3460 -1000
rect 3540 -1020 3780 -960
rect 3860 -1020 4080 -960
rect 4160 -1020 7420 -960
rect 7500 -1020 7540 -940
rect 7660 -1020 7700 -940
rect 7780 -1020 7800 -940
rect 1600 -1040 7800 -1020
rect 1600 -1220 7800 -1200
rect 1600 -1280 2920 -1220
rect 3000 -1280 3200 -1220
rect 3280 -1280 5160 -1220
rect 5240 -1280 5480 -1220
rect 5560 -1280 5780 -1220
rect 5860 -1280 6060 -1220
rect 6140 -1280 6340 -1220
rect 6420 -1280 7800 -1220
rect 1600 -1340 7800 -1280
rect 1600 -1400 5160 -1340
rect 5240 -1400 5480 -1340
rect 5560 -1400 5780 -1340
rect 5860 -1400 7800 -1340
rect 1600 -1460 7800 -1400
rect 1600 -1520 2920 -1460
rect 3000 -1520 3200 -1460
rect 3280 -1520 5160 -1460
rect 5240 -1520 5480 -1460
rect 5560 -1520 5780 -1460
rect 5860 -1520 6060 -1460
rect 6140 -1520 6340 -1460
rect 6420 -1520 7800 -1460
rect 1600 -1540 7800 -1520
rect 4560 -2040 4760 -1960
rect 4560 -2120 4620 -2040
rect 4700 -2120 4760 -2040
rect 4560 -2160 4760 -2120
rect 4560 -2240 4620 -2160
rect 4700 -2240 4760 -2160
rect 4560 -2280 4760 -2240
rect 4560 -2360 4620 -2280
rect 4700 -2360 4760 -2280
rect 4560 -2400 4760 -2360
rect 4560 -2480 4620 -2400
rect 4700 -2480 4760 -2400
rect 4560 -2520 4760 -2480
rect -3160 -2600 820 -2580
rect -3160 -2660 -600 -2600
rect -540 -2660 20 -2600
rect 80 -2660 640 -2600
rect 700 -2660 820 -2600
rect -3160 -2700 820 -2660
rect -3160 -2760 -600 -2700
rect -540 -2760 20 -2700
rect 80 -2760 640 -2700
rect 700 -2760 820 -2700
rect -3160 -2800 820 -2760
rect -3160 -2860 -600 -2800
rect -540 -2860 20 -2800
rect 80 -2860 640 -2800
rect 700 -2860 820 -2800
rect -3160 -2880 820 -2860
rect 4560 -2600 4620 -2520
rect 4700 -2600 4760 -2520
rect 12180 -2560 12480 2480
rect 4560 -2640 4760 -2600
rect 4560 -2720 4620 -2640
rect 4700 -2720 4760 -2640
rect 4560 -2760 4760 -2720
rect 4560 -2840 4620 -2760
rect 4700 -2840 4760 -2760
rect 4560 -2880 4760 -2840
rect 8540 -2580 12480 -2560
rect 8540 -2640 8640 -2580
rect 8700 -2640 9260 -2580
rect 9320 -2640 9880 -2580
rect 9940 -2640 12480 -2580
rect 8540 -2680 12480 -2640
rect 8540 -2740 8640 -2680
rect 8700 -2740 9260 -2680
rect 9320 -2740 9880 -2680
rect 9940 -2740 12480 -2680
rect 8540 -2780 12480 -2740
rect 8540 -2840 8640 -2780
rect 8700 -2840 9260 -2780
rect 9320 -2840 9880 -2780
rect 9940 -2840 12480 -2780
rect 8540 -2860 12480 -2840
rect -3160 -5560 -2860 -2880
rect 4560 -2960 4620 -2880
rect 4700 -2960 4760 -2880
rect 4560 -3000 4760 -2960
rect 4560 -3080 4620 -3000
rect 4700 -3080 4760 -3000
rect 4560 -3120 4760 -3080
rect 4560 -3200 4620 -3120
rect 4700 -3200 4760 -3120
rect 4560 -3240 4760 -3200
rect 4560 -3320 4620 -3240
rect 4700 -3320 4760 -3240
rect 4560 -3360 4760 -3320
rect 4560 -3440 4620 -3360
rect 4700 -3440 4760 -3360
rect 1200 -4160 1400 -4140
rect 1200 -4220 1220 -4160
rect 1280 -4220 1320 -4160
rect 1380 -4220 1400 -4160
rect 1200 -4260 1400 -4220
rect 1200 -4320 1220 -4260
rect 1280 -4320 1320 -4260
rect 1380 -4320 1400 -4260
rect 1200 -4340 1400 -4320
rect 4560 -4180 4760 -3440
rect 4560 -4240 4580 -4180
rect 4640 -4240 4680 -4180
rect 4740 -4240 4760 -4180
rect 4560 -4280 4760 -4240
rect 4560 -4340 4580 -4280
rect 4640 -4340 4680 -4280
rect 4740 -4340 4760 -4280
rect 8000 -4160 8200 -4140
rect 8000 -4220 8020 -4160
rect 8080 -4220 8120 -4160
rect 8180 -4220 8200 -4160
rect 8000 -4260 8200 -4220
rect 8000 -4320 8020 -4260
rect 8080 -4320 8120 -4260
rect 8180 -4320 8200 -4260
rect 8000 -4340 8200 -4320
rect 4560 -4360 4760 -4340
rect 12180 -5560 12480 -2860
rect -3160 -5640 12480 -5560
rect -3160 -5700 4560 -5640
rect 4620 -5700 4660 -5640
rect 4720 -5700 12480 -5640
rect -3160 -5740 12480 -5700
rect -3160 -5800 4560 -5740
rect 4620 -5800 4660 -5740
rect 4720 -5800 12480 -5740
rect -3160 -5860 12480 -5800
<< via2 >>
rect -1640 3360 -1580 3420
rect -1540 3360 -1480 3420
rect -1440 3360 -1380 3420
rect -1340 3360 -1280 3420
rect -1640 3220 -1580 3280
rect -1540 3220 -1480 3280
rect -1440 3220 -1380 3280
rect -1340 3220 -1280 3280
rect 10640 3360 10700 3420
rect 10740 3360 10800 3420
rect 10840 3360 10900 3420
rect 10940 3360 11000 3420
rect 10640 3220 10700 3280
rect 10740 3220 10800 3280
rect 10840 3220 10900 3280
rect 10940 3220 11000 3280
rect 7420 2520 7500 2600
rect 7560 2520 7640 2600
rect 7700 2520 7780 2600
rect 7420 2300 7500 2380
rect 7560 2300 7640 2380
rect 7700 2300 7780 2380
rect 1620 1320 1700 1400
rect 1760 1320 1840 1400
rect 1900 1320 1980 1400
rect 1620 1140 1700 1220
rect 1760 1140 1840 1220
rect 1900 1140 1980 1220
rect 7420 1300 7500 1380
rect 7560 1300 7640 1380
rect 7700 1300 7780 1380
rect 7420 1120 7500 1200
rect 7560 1120 7640 1200
rect 7700 1120 7780 1200
rect 1620 140 1700 220
rect 1740 140 1860 220
rect 1900 140 1980 220
rect 7420 140 7500 220
rect 7540 140 7660 220
rect 7700 140 7780 220
rect 1620 -80 1700 0
rect 1740 -80 1860 0
rect 1900 -80 1980 0
rect 7420 -80 7500 0
rect 7540 -80 7660 0
rect 7700 -80 7780 0
rect 1140 -300 1220 -220
rect 1260 -300 1360 -220
rect 1400 -300 1480 -220
rect 1140 -440 1220 -360
rect 1260 -440 1360 -360
rect 1400 -440 1480 -360
rect 7920 -300 8000 -220
rect 8040 -300 8140 -220
rect 8180 -300 8260 -220
rect 7920 -440 8000 -360
rect 8040 -440 8140 -360
rect 8180 -440 8260 -360
rect 1140 -580 1220 -500
rect 1260 -580 1360 -500
rect 1400 -580 1480 -500
rect 7920 -580 8000 -500
rect 8040 -580 8140 -500
rect 8180 -580 8260 -500
rect 1620 -800 1700 -720
rect 1740 -800 1860 -720
rect 1900 -800 1980 -720
rect 7420 -800 7500 -720
rect 7540 -800 7660 -720
rect 7700 -800 7780 -720
rect 1620 -1000 1700 -920
rect 1740 -1000 1860 -920
rect 1900 -1000 1980 -920
rect 7420 -1020 7500 -940
rect 7540 -1020 7660 -940
rect 7700 -1020 7780 -940
rect 1220 -4220 1280 -4160
rect 1320 -4220 1380 -4160
rect 1220 -4320 1280 -4260
rect 1320 -4320 1380 -4260
rect 8020 -4220 8080 -4160
rect 8120 -4220 8180 -4160
rect 8020 -4320 8080 -4260
rect 8120 -4320 8180 -4260
<< metal3 >>
rect -1660 3420 -1260 3558
rect -1660 3360 -1640 3420
rect -1580 3360 -1540 3420
rect -1480 3360 -1440 3420
rect -1380 3360 -1340 3420
rect -1280 3360 -1260 3420
rect -1660 3280 -1260 3360
rect -1660 3220 -1640 3280
rect -1580 3220 -1540 3280
rect -1480 3220 -1440 3280
rect -1380 3220 -1340 3280
rect -1280 3220 -1260 3280
rect -1660 2160 -1260 3220
rect 10620 3420 11014 3558
rect 10620 3360 10640 3420
rect 10700 3360 10740 3420
rect 10800 3360 10840 3420
rect 10900 3360 10940 3420
rect 11000 3360 11020 3420
rect 10620 3280 11020 3360
rect 10620 3220 10640 3280
rect 10700 3220 10740 3280
rect 10800 3220 10840 3280
rect 10900 3220 10940 3280
rect 11000 3220 11020 3280
rect 1600 2600 2000 2620
rect 1600 2520 1620 2600
rect 1700 2520 1760 2600
rect 1840 2520 1900 2600
rect 1980 2520 2000 2600
rect 1600 2380 2000 2520
rect 1600 2300 1620 2380
rect 1700 2300 1760 2380
rect 1840 2300 1900 2380
rect 1980 2300 2000 2380
rect 1600 2280 2000 2300
rect 7400 2600 7800 2620
rect 7400 2520 7420 2600
rect 7500 2520 7560 2600
rect 7640 2520 7700 2600
rect 7780 2520 7800 2600
rect 7400 2380 7800 2520
rect 7400 2300 7420 2380
rect 7500 2300 7560 2380
rect 7640 2300 7700 2380
rect 7780 2300 7800 2380
rect 7400 2280 7800 2300
rect -1660 2080 -1640 2160
rect -1560 2080 -1500 2160
rect -1420 2080 -1360 2160
rect -1280 2080 -1260 2160
rect -1660 1980 -1260 2080
rect -1660 1900 -1640 1980
rect -1560 1900 -1500 1980
rect -1420 1900 -1360 1980
rect -1280 1900 -1260 1980
rect -1660 1220 -1260 1900
rect 10620 2160 11020 3220
rect 10620 2080 10640 2160
rect 10720 2080 10780 2160
rect 10860 2080 10920 2160
rect 11000 2080 11020 2160
rect 10620 1980 11020 2080
rect 10620 1900 10640 1980
rect 10720 1900 10780 1980
rect 10860 1900 10920 1980
rect 11000 1900 11020 1980
rect 1600 1400 2000 1420
rect 1600 1320 1620 1400
rect 1700 1320 1760 1400
rect 1840 1320 1900 1400
rect 1980 1320 2000 1400
rect 1600 1220 2000 1320
rect -1660 -3560 -1280 1220
rect 1600 1140 1620 1220
rect 1700 1140 1760 1220
rect 1840 1140 1900 1220
rect 1980 1140 2000 1220
rect 1600 1120 2000 1140
rect 7400 1380 7800 1400
rect 7400 1300 7420 1380
rect 7500 1300 7560 1380
rect 7640 1300 7700 1380
rect 7780 1300 7800 1380
rect 7400 1200 7800 1300
rect 10620 1200 11020 1900
rect 7400 1120 7420 1200
rect 7500 1120 7560 1200
rect 7640 1120 7700 1200
rect 7780 1120 7800 1200
rect 7400 1100 7800 1120
rect 1600 220 2000 240
rect 1600 140 1620 220
rect 1700 140 1740 220
rect 1860 140 1900 220
rect 1980 140 2000 220
rect 1600 0 2000 140
rect 1600 -80 1620 0
rect 1700 -80 1740 0
rect 1860 -80 1900 0
rect 1980 -80 2000 0
rect 1600 -100 2000 -80
rect 7400 220 7800 240
rect 7400 140 7420 220
rect 7500 140 7540 220
rect 7660 140 7700 220
rect 7780 140 7800 220
rect 7400 0 7800 140
rect 7400 -80 7420 0
rect 7500 -80 7540 0
rect 7660 -80 7700 0
rect 7780 -80 7800 0
rect 7400 -100 7800 -80
rect 1120 -220 1500 -200
rect 1120 -300 1140 -220
rect 1220 -300 1260 -220
rect 1360 -300 1400 -220
rect 1480 -300 1500 -220
rect 1120 -360 1500 -300
rect 1120 -440 1140 -360
rect 1220 -440 1260 -360
rect 1360 -440 1400 -360
rect 1480 -440 1500 -360
rect 1120 -500 1500 -440
rect 1120 -580 1140 -500
rect 1220 -580 1260 -500
rect 1360 -580 1400 -500
rect 1480 -580 1500 -500
rect 1120 -4160 1500 -580
rect 7900 -220 8280 -200
rect 7900 -300 7920 -220
rect 8000 -300 8040 -220
rect 8140 -300 8180 -220
rect 8260 -300 8280 -220
rect 7900 -360 8280 -300
rect 7900 -440 7920 -360
rect 8000 -440 8040 -360
rect 8140 -440 8180 -360
rect 8260 -440 8280 -360
rect 7900 -500 8280 -440
rect 7900 -580 7920 -500
rect 8000 -580 8040 -500
rect 8140 -580 8180 -500
rect 8260 -580 8280 -500
rect 1600 -720 2000 -700
rect 1600 -800 1620 -720
rect 1700 -800 1740 -720
rect 1860 -800 1900 -720
rect 1980 -800 2000 -720
rect 1600 -920 2000 -800
rect 1600 -1000 1620 -920
rect 1700 -1000 1740 -920
rect 1860 -1000 1900 -920
rect 1980 -1000 2000 -920
rect 1600 -1040 2000 -1000
rect 7400 -720 7800 -700
rect 7400 -800 7420 -720
rect 7500 -800 7540 -720
rect 7660 -800 7700 -720
rect 7780 -800 7800 -720
rect 7400 -940 7800 -800
rect 7400 -1020 7420 -940
rect 7500 -1020 7540 -940
rect 7660 -1020 7700 -940
rect 7780 -1020 7800 -940
rect 7400 -1040 7800 -1020
rect 1120 -4220 1220 -4160
rect 1280 -4220 1320 -4160
rect 1380 -4220 1500 -4160
rect 1120 -4260 1500 -4220
rect 1120 -4320 1220 -4260
rect 1280 -4320 1320 -4260
rect 1380 -4320 1500 -4260
rect 1120 -4340 1500 -4320
rect 7900 -4160 8280 -580
rect 10640 -3560 11020 1200
rect 7900 -4220 8020 -4160
rect 8080 -4220 8120 -4160
rect 8180 -4220 8280 -4160
rect 7900 -4260 8280 -4220
rect 7900 -4320 8020 -4260
rect 8080 -4320 8120 -4260
rect 8180 -4320 8280 -4260
rect 7900 -4340 8280 -4320
<< via3 >>
rect 1620 2520 1700 2600
rect 1760 2520 1840 2600
rect 1900 2520 1980 2600
rect 1620 2300 1700 2380
rect 1760 2300 1840 2380
rect 1900 2300 1980 2380
rect 7420 2520 7500 2600
rect 7560 2520 7640 2600
rect 7700 2520 7780 2600
rect 7420 2300 7500 2380
rect 7560 2300 7640 2380
rect 7700 2300 7780 2380
rect -1640 2080 -1560 2160
rect -1500 2080 -1420 2160
rect -1360 2080 -1280 2160
rect -1640 1900 -1560 1980
rect -1500 1900 -1420 1980
rect -1360 1900 -1280 1980
rect 10640 2080 10720 2160
rect 10780 2080 10860 2160
rect 10920 2080 11000 2160
rect 10640 1900 10720 1980
rect 10780 1900 10860 1980
rect 10920 1900 11000 1980
rect 1620 1320 1700 1400
rect 1760 1320 1840 1400
rect 1900 1320 1980 1400
rect 1620 1140 1700 1220
rect 1760 1140 1840 1220
rect 1900 1140 1980 1220
rect 7420 1300 7500 1380
rect 7560 1300 7640 1380
rect 7700 1300 7780 1380
rect 7420 1120 7500 1200
rect 7560 1120 7640 1200
rect 7700 1120 7780 1200
rect 1620 140 1700 220
rect 1740 140 1860 220
rect 1900 140 1980 220
rect 1620 -80 1700 0
rect 1740 -80 1860 0
rect 1900 -80 1980 0
rect 7420 140 7500 220
rect 7540 140 7660 220
rect 7700 140 7780 220
rect 7420 -80 7500 0
rect 7540 -80 7660 0
rect 7700 -80 7780 0
rect 1620 -800 1700 -720
rect 1740 -800 1860 -720
rect 1900 -800 1980 -720
rect 1620 -1000 1700 -920
rect 1740 -1000 1860 -920
rect 1900 -1000 1980 -920
rect 7420 -800 7500 -720
rect 7540 -800 7660 -720
rect 7700 -800 7780 -720
rect 7420 -1020 7500 -940
rect 7540 -1020 7660 -940
rect 7700 -1020 7780 -940
<< metal4 >>
rect -17200 6720 -16500 7100
rect 25980 6720 26680 7100
rect -17200 2180 -16860 6720
rect 1600 2600 2000 4140
rect 1600 2520 1620 2600
rect 1700 2520 1760 2600
rect 1840 2520 1900 2600
rect 1980 2520 2000 2600
rect 1600 2380 2000 2520
rect 1600 2300 1620 2380
rect 1700 2300 1760 2380
rect 1840 2300 1900 2380
rect 1980 2300 2000 2380
rect -17200 2160 -1200 2180
rect -17200 2080 -1640 2160
rect -1560 2080 -1500 2160
rect -1420 2080 -1360 2160
rect -1280 2080 -1200 2160
rect -17200 1980 -1200 2080
rect -17200 1900 -1640 1980
rect -1560 1900 -1500 1980
rect -1420 1900 -1360 1980
rect -1280 1900 -1200 1980
rect -17200 1880 -1200 1900
rect 1600 1400 2000 2300
rect 1600 1320 1620 1400
rect 1700 1320 1760 1400
rect 1840 1320 1900 1400
rect 1980 1320 2000 1400
rect 1600 1220 2000 1320
rect 1600 1140 1620 1220
rect 1700 1140 1760 1220
rect 1840 1140 1900 1220
rect 1980 1140 2000 1220
rect 1600 220 2000 1140
rect 1600 140 1620 220
rect 1700 140 1740 220
rect 1860 140 1900 220
rect 1980 140 2000 220
rect 1600 0 2000 140
rect 1600 -80 1620 0
rect 1700 -80 1740 0
rect 1860 -80 1900 0
rect 1980 -80 2000 0
rect 1600 -720 2000 -80
rect 1600 -800 1620 -720
rect 1700 -800 1740 -720
rect 1860 -800 1900 -720
rect 1980 -800 2000 -720
rect 1600 -920 2000 -800
rect 1600 -1000 1620 -920
rect 1700 -1000 1740 -920
rect 1860 -1000 1900 -920
rect 1980 -1000 2000 -920
rect 1600 -3560 2000 -1000
rect 7400 2600 7800 4140
rect 7400 2520 7420 2600
rect 7500 2520 7560 2600
rect 7640 2520 7700 2600
rect 7780 2520 7800 2600
rect 7400 2380 7800 2520
rect 7400 2300 7420 2380
rect 7500 2300 7560 2380
rect 7640 2300 7700 2380
rect 7780 2300 7800 2380
rect 7400 1380 7800 2300
rect 26340 2180 26680 6720
rect 10620 2160 26680 2180
rect 10620 2080 10640 2160
rect 10720 2080 10780 2160
rect 10860 2080 10920 2160
rect 11000 2080 26680 2160
rect 10620 1980 26680 2080
rect 10620 1900 10640 1980
rect 10720 1900 10780 1980
rect 10860 1900 10920 1980
rect 11000 1900 26680 1980
rect 10620 1880 26680 1900
rect 7400 1300 7420 1380
rect 7500 1300 7560 1380
rect 7640 1300 7700 1380
rect 7780 1300 7800 1380
rect 7400 1200 7800 1300
rect 7400 1120 7420 1200
rect 7500 1120 7560 1200
rect 7640 1120 7700 1200
rect 7780 1120 7800 1200
rect 7400 220 7800 1120
rect 7400 140 7420 220
rect 7500 140 7540 220
rect 7660 140 7700 220
rect 7780 140 7800 220
rect 7400 0 7800 140
rect 7400 -80 7420 0
rect 7500 -80 7540 0
rect 7660 -80 7700 0
rect 7780 -80 7800 0
rect 7400 -720 7800 -80
rect 7400 -800 7420 -720
rect 7500 -800 7540 -720
rect 7660 -800 7700 -720
rect 7780 -800 7800 -720
rect 7400 -940 7800 -800
rect 7400 -1020 7420 -940
rect 7500 -1020 7540 -940
rect 7660 -1020 7700 -940
rect 7780 -1020 7800 -940
rect 7400 -3560 7800 -1020
use sky130_fd_pr__cap_mim_m3_1_R7S84X  sky130_fd_pr__cap_mim_m3_1_R7S84X_0
timestamp 1769535502
transform 0 1 4740 -1 0 6726
box -2686 -21280 2686 21280
use sky130_fd_pr__nfet_g5v0d10v5_A8KA9K  sky130_fd_pr__nfet_g5v0d10v5_A8KA9K_0
timestamp 1769535502
transform 1 0 5517 0 1 288
box -515 -698 515 698
use sky130_fd_pr__nfet_g5v0d10v5_N5GNFR  sky130_fd_pr__nfet_g5v0d10v5_N5GNFR_0
timestamp 1769529800
transform 1 0 55 0 1 -2663
box -815 -977 815 977
use sky130_fd_pr__nfet_g5v0d10v5_PBQQNH  sky130_fd_pr__nfet_g5v0d10v5_PBQQNH_0
timestamp 1769535502
transform 1 0 3815 0 1 -1102
box -515 -698 515 698
use sky130_fd_pr__nfet_g5v0d10v5_X6KG9Z  sky130_fd_pr__nfet_g5v0d10v5_X6KG9Z_0
timestamp 1769529800
transform 1 0 5515 0 1 -1102
box -515 -698 515 698
use sky130_fd_pr__pfet_g5v0d10v5_RFPNS8  sky130_fd_pr__pfet_g5v0d10v5_RFPNS8_0
timestamp 1769535502
transform 1 0 81 0 1 2422
box -1461 -1262 1461 1262
use sky130_fd_pr__pfet_g5v0d10v5_V6JW4R  sky130_fd_pr__pfet_g5v0d10v5_V6JW4R_0
timestamp 1769571357
transform -1 0 -2133 0 -1 2922
box -467 -762 467 762
use sky130_fd_pr__pfet_g5v0d10v5_V6JW4R  sky130_fd_pr__pfet_g5v0d10v5_V6JW4R_1
timestamp 1769571357
transform -1 0 11447 0 -1 2902
box -467 -762 467 762
use sky130_fd_pr__pfet_g5v0d10v5_S5VYLR  XM2
timestamp 1769535502
transform 1 0 4673 0 1 2462
box -2693 -1202 2693 1202
use sky130_fd_pr__nfet_g5v0d10v5_DC2CKB  XM3
timestamp 1769529800
transform 1 0 3815 0 1 298
box -515 -698 515 698
use sky130_fd_pr__nfet_g5v0d10v5_2899RY  XM5
timestamp 1769535502
transform 1 0 4663 0 1 -2663
box -2663 -977 2663 977
use sky130_fd_pr__pfet_g5v0d10v5_RFPNS8  XM7
timestamp 1769535502
transform 1 0 9281 0 1 2402
box -1461 -1262 1461 1262
use sky130_fd_pr__nfet_g5v0d10v5_N5GNFR  XM8
timestamp 1769529800
transform 1 0 9295 0 1 -2683
box -815 -977 815 977
<< labels >>
flabel metal1 -2600 -3800 -2400 -3600 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 -2600 3600 -2400 3800 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 4560 -4360 4760 -4160 0 FreeSans 256 0 0 0 IBIAS
port 4 nsew
flabel metal1 8000 -4340 8200 -4140 0 FreeSans 256 0 0 0 VP
port 2 nsew
flabel metal1 4540 -5820 4740 -5620 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 1200 -4340 1400 -4140 0 FreeSans 256 0 0 0 VN
port 3 nsew
<< end >>
