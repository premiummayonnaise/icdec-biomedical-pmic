magic
tech sky130A
magscale 1 2
timestamp 1769400417
<< nmos >>
rect -279 -371 -29 309
rect 29 -371 279 309
<< ndiff >>
rect -337 297 -279 309
rect -337 -359 -325 297
rect -291 -359 -279 297
rect -337 -371 -279 -359
rect -29 297 29 309
rect -29 -359 -17 297
rect 17 -359 29 297
rect -29 -371 29 -359
rect 279 297 337 309
rect 279 -359 291 297
rect 325 -359 337 297
rect 279 -371 337 -359
<< ndiffc >>
rect -325 -359 -291 297
rect -17 -359 17 297
rect 291 -359 325 297
<< poly >>
rect -279 381 -29 397
rect -279 347 -263 381
rect -45 347 -29 381
rect -279 309 -29 347
rect 29 381 279 397
rect 29 347 45 381
rect 263 347 279 381
rect 29 309 279 347
rect -279 -397 -29 -371
rect 29 -397 279 -371
<< polycont >>
rect -263 347 -45 381
rect 45 347 263 381
<< locali >>
rect -279 347 -263 381
rect -45 347 -29 381
rect 29 347 45 381
rect 263 347 279 381
rect -325 297 -291 313
rect -325 -375 -291 -359
rect -17 297 17 313
rect -17 -375 17 -359
rect 291 297 325 313
rect 291 -375 325 -359
<< viali >>
rect -263 347 -45 381
rect 45 347 263 381
rect -325 -359 -291 297
rect -17 -359 17 297
rect 291 -359 325 297
<< metal1 >>
rect -275 381 -33 387
rect -275 347 -263 381
rect -45 347 -33 381
rect -275 341 -33 347
rect 33 381 275 387
rect 33 347 45 381
rect 263 347 275 381
rect 33 341 275 347
rect -331 297 -285 309
rect -331 -359 -325 297
rect -291 -359 -285 297
rect -331 -371 -285 -359
rect -23 297 23 309
rect -23 -359 -17 297
rect 17 -359 23 297
rect -23 -371 23 -359
rect 285 297 331 309
rect 285 -359 291 297
rect 325 -359 331 297
rect 285 -371 331 -359
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.4 l 1.25 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
