magic
tech sky130A
magscale 1 2
timestamp 1769535502
<< metal3 >>
rect -2686 21132 2686 21160
rect -2686 16108 2602 21132
rect 2666 16108 2686 21132
rect -2686 16080 2686 16108
rect -2686 15812 2686 15840
rect -2686 10788 2602 15812
rect 2666 10788 2686 15812
rect -2686 10760 2686 10788
rect -2686 10492 2686 10520
rect -2686 5468 2602 10492
rect 2666 5468 2686 10492
rect -2686 5440 2686 5468
rect -2686 5172 2686 5200
rect -2686 148 2602 5172
rect 2666 148 2686 5172
rect -2686 120 2686 148
rect -2686 -148 2686 -120
rect -2686 -5172 2602 -148
rect 2666 -5172 2686 -148
rect -2686 -5200 2686 -5172
rect -2686 -5468 2686 -5440
rect -2686 -10492 2602 -5468
rect 2666 -10492 2686 -5468
rect -2686 -10520 2686 -10492
rect -2686 -10788 2686 -10760
rect -2686 -15812 2602 -10788
rect 2666 -15812 2686 -10788
rect -2686 -15840 2686 -15812
rect -2686 -16108 2686 -16080
rect -2686 -21132 2602 -16108
rect 2666 -21132 2686 -16108
rect -2686 -21160 2686 -21132
<< via3 >>
rect 2602 16108 2666 21132
rect 2602 10788 2666 15812
rect 2602 5468 2666 10492
rect 2602 148 2666 5172
rect 2602 -5172 2666 -148
rect 2602 -10492 2666 -5468
rect 2602 -15812 2666 -10788
rect 2602 -21132 2666 -16108
<< mimcap >>
rect -2646 21080 2354 21120
rect -2646 16160 -2606 21080
rect 2314 16160 2354 21080
rect -2646 16120 2354 16160
rect -2646 15760 2354 15800
rect -2646 10840 -2606 15760
rect 2314 10840 2354 15760
rect -2646 10800 2354 10840
rect -2646 10440 2354 10480
rect -2646 5520 -2606 10440
rect 2314 5520 2354 10440
rect -2646 5480 2354 5520
rect -2646 5120 2354 5160
rect -2646 200 -2606 5120
rect 2314 200 2354 5120
rect -2646 160 2354 200
rect -2646 -200 2354 -160
rect -2646 -5120 -2606 -200
rect 2314 -5120 2354 -200
rect -2646 -5160 2354 -5120
rect -2646 -5520 2354 -5480
rect -2646 -10440 -2606 -5520
rect 2314 -10440 2354 -5520
rect -2646 -10480 2354 -10440
rect -2646 -10840 2354 -10800
rect -2646 -15760 -2606 -10840
rect 2314 -15760 2354 -10840
rect -2646 -15800 2354 -15760
rect -2646 -16160 2354 -16120
rect -2646 -21080 -2606 -16160
rect 2314 -21080 2354 -16160
rect -2646 -21120 2354 -21080
<< mimcapcontact >>
rect -2606 16160 2314 21080
rect -2606 10840 2314 15760
rect -2606 5520 2314 10440
rect -2606 200 2314 5120
rect -2606 -5120 2314 -200
rect -2606 -10440 2314 -5520
rect -2606 -15760 2314 -10840
rect -2606 -21080 2314 -16160
<< metal4 >>
rect -198 21081 -94 21280
rect 2582 21132 2686 21280
rect -2607 21080 2315 21081
rect -2607 16160 -2606 21080
rect 2314 16160 2315 21080
rect -2607 16159 2315 16160
rect -198 15761 -94 16159
rect 2582 16108 2602 21132
rect 2666 16108 2686 21132
rect 2582 15812 2686 16108
rect -2607 15760 2315 15761
rect -2607 10840 -2606 15760
rect 2314 10840 2315 15760
rect -2607 10839 2315 10840
rect -198 10441 -94 10839
rect 2582 10788 2602 15812
rect 2666 10788 2686 15812
rect 2582 10492 2686 10788
rect -2607 10440 2315 10441
rect -2607 5520 -2606 10440
rect 2314 5520 2315 10440
rect -2607 5519 2315 5520
rect -198 5121 -94 5519
rect 2582 5468 2602 10492
rect 2666 5468 2686 10492
rect 2582 5172 2686 5468
rect -2607 5120 2315 5121
rect -2607 200 -2606 5120
rect 2314 200 2315 5120
rect -2607 199 2315 200
rect -198 -199 -94 199
rect 2582 148 2602 5172
rect 2666 148 2686 5172
rect 2582 -148 2686 148
rect -2607 -200 2315 -199
rect -2607 -5120 -2606 -200
rect 2314 -5120 2315 -200
rect -2607 -5121 2315 -5120
rect -198 -5519 -94 -5121
rect 2582 -5172 2602 -148
rect 2666 -5172 2686 -148
rect 2582 -5468 2686 -5172
rect -2607 -5520 2315 -5519
rect -2607 -10440 -2606 -5520
rect 2314 -10440 2315 -5520
rect -2607 -10441 2315 -10440
rect -198 -10839 -94 -10441
rect 2582 -10492 2602 -5468
rect 2666 -10492 2686 -5468
rect 2582 -10788 2686 -10492
rect -2607 -10840 2315 -10839
rect -2607 -15760 -2606 -10840
rect 2314 -15760 2315 -10840
rect -2607 -15761 2315 -15760
rect -198 -16159 -94 -15761
rect 2582 -15812 2602 -10788
rect 2666 -15812 2686 -10788
rect 2582 -16108 2686 -15812
rect -2607 -16160 2315 -16159
rect -2607 -21080 -2606 -16160
rect 2314 -21080 2315 -16160
rect -2607 -21081 2315 -21080
rect -198 -21280 -94 -21081
rect 2582 -21132 2602 -16108
rect 2666 -21132 2686 -16108
rect 2582 -21280 2686 -21132
<< properties >>
string FIXED_BBOX -2686 16080 2394 21160
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 25.0 val 1.269k carea 2.00 cperi 0.19 class capacitor nx 1 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
