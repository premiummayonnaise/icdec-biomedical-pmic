magic
tech sky130A
magscale 1 2
timestamp 1769172933
<< error_p >>
rect -1747 -568 -1717 500
rect -1681 -502 -1651 434
rect 1651 -502 1681 434
rect -1681 -506 -1315 -502
rect -1253 -506 -887 -502
rect -825 -506 -459 -502
rect -397 -506 -31 -502
rect 31 -506 397 -502
rect 459 -506 825 -502
rect 887 -506 1253 -502
rect 1315 -506 1681 -502
rect 1717 -568 1747 500
rect -1747 -572 1747 -568
<< nwell >>
rect -1717 -568 1717 534
<< mvpmos >>
rect -1623 -506 -1373 434
rect -1195 -506 -945 434
rect -767 -506 -517 434
rect -339 -506 -89 434
rect 89 -506 339 434
rect 517 -506 767 434
rect 945 -506 1195 434
rect 1373 -506 1623 434
<< mvpdiff >>
rect -1681 422 -1623 434
rect -1681 -494 -1669 422
rect -1635 -494 -1623 422
rect -1681 -506 -1623 -494
rect -1373 422 -1315 434
rect -1373 -494 -1361 422
rect -1327 -494 -1315 422
rect -1373 -506 -1315 -494
rect -1253 422 -1195 434
rect -1253 -494 -1241 422
rect -1207 -494 -1195 422
rect -1253 -506 -1195 -494
rect -945 422 -887 434
rect -945 -494 -933 422
rect -899 -494 -887 422
rect -945 -506 -887 -494
rect -825 422 -767 434
rect -825 -494 -813 422
rect -779 -494 -767 422
rect -825 -506 -767 -494
rect -517 422 -459 434
rect -517 -494 -505 422
rect -471 -494 -459 422
rect -517 -506 -459 -494
rect -397 422 -339 434
rect -397 -494 -385 422
rect -351 -494 -339 422
rect -397 -506 -339 -494
rect -89 422 -31 434
rect -89 -494 -77 422
rect -43 -494 -31 422
rect -89 -506 -31 -494
rect 31 422 89 434
rect 31 -494 43 422
rect 77 -494 89 422
rect 31 -506 89 -494
rect 339 422 397 434
rect 339 -494 351 422
rect 385 -494 397 422
rect 339 -506 397 -494
rect 459 422 517 434
rect 459 -494 471 422
rect 505 -494 517 422
rect 459 -506 517 -494
rect 767 422 825 434
rect 767 -494 779 422
rect 813 -494 825 422
rect 767 -506 825 -494
rect 887 422 945 434
rect 887 -494 899 422
rect 933 -494 945 422
rect 887 -506 945 -494
rect 1195 422 1253 434
rect 1195 -494 1207 422
rect 1241 -494 1253 422
rect 1195 -506 1253 -494
rect 1315 422 1373 434
rect 1315 -494 1327 422
rect 1361 -494 1373 422
rect 1315 -506 1373 -494
rect 1623 422 1681 434
rect 1623 -494 1635 422
rect 1669 -494 1681 422
rect 1623 -506 1681 -494
<< mvpdiffc >>
rect -1669 -494 -1635 422
rect -1361 -494 -1327 422
rect -1241 -494 -1207 422
rect -933 -494 -899 422
rect -813 -494 -779 422
rect -505 -494 -471 422
rect -385 -494 -351 422
rect -77 -494 -43 422
rect 43 -494 77 422
rect 351 -494 385 422
rect 471 -494 505 422
rect 779 -494 813 422
rect 899 -494 933 422
rect 1207 -494 1241 422
rect 1327 -494 1361 422
rect 1635 -494 1669 422
<< poly >>
rect -1623 515 -1373 531
rect -1623 481 -1607 515
rect -1389 481 -1373 515
rect -1623 434 -1373 481
rect -1195 515 -945 531
rect -1195 481 -1179 515
rect -961 481 -945 515
rect -1195 434 -945 481
rect -767 515 -517 531
rect -767 481 -751 515
rect -533 481 -517 515
rect -767 434 -517 481
rect -339 515 -89 531
rect -339 481 -323 515
rect -105 481 -89 515
rect -339 434 -89 481
rect 89 515 339 531
rect 89 481 105 515
rect 323 481 339 515
rect 89 434 339 481
rect 517 515 767 531
rect 517 481 533 515
rect 751 481 767 515
rect 517 434 767 481
rect 945 515 1195 531
rect 945 481 961 515
rect 1179 481 1195 515
rect 945 434 1195 481
rect 1373 515 1623 531
rect 1373 481 1389 515
rect 1607 481 1623 515
rect 1373 434 1623 481
rect -1623 -532 -1373 -506
rect -1195 -532 -945 -506
rect -767 -532 -517 -506
rect -339 -532 -89 -506
rect 89 -532 339 -506
rect 517 -532 767 -506
rect 945 -532 1195 -506
rect 1373 -532 1623 -506
<< polycont >>
rect -1607 481 -1389 515
rect -1179 481 -961 515
rect -751 481 -533 515
rect -323 481 -105 515
rect 105 481 323 515
rect 533 481 751 515
rect 961 481 1179 515
rect 1389 481 1607 515
<< locali >>
rect -1623 481 -1607 515
rect -1389 481 -1373 515
rect -1195 481 -1179 515
rect -961 481 -945 515
rect -767 481 -751 515
rect -533 481 -517 515
rect -339 481 -323 515
rect -105 481 -89 515
rect 89 481 105 515
rect 323 481 339 515
rect 517 481 533 515
rect 751 481 767 515
rect 945 481 961 515
rect 1179 481 1195 515
rect 1373 481 1389 515
rect 1607 481 1623 515
rect -1669 422 -1635 438
rect -1669 -510 -1635 -494
rect -1361 422 -1327 438
rect -1361 -510 -1327 -494
rect -1241 422 -1207 438
rect -1241 -510 -1207 -494
rect -933 422 -899 438
rect -933 -510 -899 -494
rect -813 422 -779 438
rect -813 -510 -779 -494
rect -505 422 -471 438
rect -505 -510 -471 -494
rect -385 422 -351 438
rect -385 -510 -351 -494
rect -77 422 -43 438
rect -77 -510 -43 -494
rect 43 422 77 438
rect 43 -510 77 -494
rect 351 422 385 438
rect 351 -510 385 -494
rect 471 422 505 438
rect 471 -510 505 -494
rect 779 422 813 438
rect 779 -510 813 -494
rect 899 422 933 438
rect 899 -510 933 -494
rect 1207 422 1241 438
rect 1207 -510 1241 -494
rect 1327 422 1361 438
rect 1327 -510 1361 -494
rect 1635 422 1669 438
rect 1635 -510 1669 -494
<< viali >>
rect -1607 481 -1389 515
rect -1179 481 -961 515
rect -751 481 -533 515
rect -323 481 -105 515
rect 105 481 323 515
rect 533 481 751 515
rect 961 481 1179 515
rect 1389 481 1607 515
rect -1669 -494 -1635 422
rect -1361 -494 -1327 422
rect -1241 -494 -1207 422
rect -933 -494 -899 422
rect -813 -494 -779 422
rect -505 -494 -471 422
rect -385 -494 -351 422
rect -77 -494 -43 422
rect 43 -494 77 422
rect 351 -494 385 422
rect 471 -494 505 422
rect 779 -494 813 422
rect 899 -494 933 422
rect 1207 -494 1241 422
rect 1327 -494 1361 422
rect 1635 -494 1669 422
<< metal1 >>
rect -1619 515 -1377 521
rect -1619 481 -1607 515
rect -1389 481 -1377 515
rect -1619 475 -1377 481
rect -1191 515 -949 521
rect -1191 481 -1179 515
rect -961 481 -949 515
rect -1191 475 -949 481
rect -763 515 -521 521
rect -763 481 -751 515
rect -533 481 -521 515
rect -763 475 -521 481
rect -335 515 -93 521
rect -335 481 -323 515
rect -105 481 -93 515
rect -335 475 -93 481
rect 93 515 335 521
rect 93 481 105 515
rect 323 481 335 515
rect 93 475 335 481
rect 521 515 763 521
rect 521 481 533 515
rect 751 481 763 515
rect 521 475 763 481
rect 949 515 1191 521
rect 949 481 961 515
rect 1179 481 1191 515
rect 949 475 1191 481
rect 1377 515 1619 521
rect 1377 481 1389 515
rect 1607 481 1619 515
rect 1377 475 1619 481
rect -1675 422 -1629 434
rect -1675 -494 -1669 422
rect -1635 -494 -1629 422
rect -1675 -506 -1629 -494
rect -1367 422 -1321 434
rect -1367 -494 -1361 422
rect -1327 -494 -1321 422
rect -1367 -506 -1321 -494
rect -1247 422 -1201 434
rect -1247 -494 -1241 422
rect -1207 -494 -1201 422
rect -1247 -506 -1201 -494
rect -939 422 -893 434
rect -939 -494 -933 422
rect -899 -494 -893 422
rect -939 -506 -893 -494
rect -819 422 -773 434
rect -819 -494 -813 422
rect -779 -494 -773 422
rect -819 -506 -773 -494
rect -511 422 -465 434
rect -511 -494 -505 422
rect -471 -494 -465 422
rect -511 -506 -465 -494
rect -391 422 -345 434
rect -391 -494 -385 422
rect -351 -494 -345 422
rect -391 -506 -345 -494
rect -83 422 -37 434
rect -83 -494 -77 422
rect -43 -494 -37 422
rect -83 -506 -37 -494
rect 37 422 83 434
rect 37 -494 43 422
rect 77 -494 83 422
rect 37 -506 83 -494
rect 345 422 391 434
rect 345 -494 351 422
rect 385 -494 391 422
rect 345 -506 391 -494
rect 465 422 511 434
rect 465 -494 471 422
rect 505 -494 511 422
rect 465 -506 511 -494
rect 773 422 819 434
rect 773 -494 779 422
rect 813 -494 819 422
rect 773 -506 819 -494
rect 893 422 939 434
rect 893 -494 899 422
rect 933 -494 939 422
rect 893 -506 939 -494
rect 1201 422 1247 434
rect 1201 -494 1207 422
rect 1241 -494 1247 422
rect 1201 -506 1247 -494
rect 1321 422 1367 434
rect 1321 -494 1327 422
rect 1361 -494 1367 422
rect 1321 -506 1367 -494
rect 1629 422 1675 434
rect 1629 -494 1635 422
rect 1669 -494 1675 422
rect 1629 -506 1675 -494
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.7 l 1.25 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
