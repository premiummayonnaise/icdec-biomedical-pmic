magic
tech sky130A
timestamp 1770345528
<< psubdiff >>
rect -1995 -7250 -1425 -7125
rect -1995 -7550 -1850 -7250
rect -1550 -7550 -1425 -7250
rect -1995 -7695 -1425 -7550
<< psubdiffcont >>
rect -1850 -7550 -1550 -7250
<< xpolycontact >>
rect -1995 285 -1710 570
rect 1140 -18525 1425 -18240
<< xpolyres >>
rect -1710 285 1425 570
rect 1140 -2565 1425 285
rect -1995 -2850 1425 -2565
rect -1995 -5700 -1710 -2850
rect -1995 -5985 1425 -5700
rect 1140 -8835 1425 -5985
rect -1995 -9120 1425 -8835
rect -1995 -11970 -1710 -9120
rect -1995 -12255 1425 -11970
rect 1140 -15105 1425 -12255
rect -1995 -15390 1425 -15105
rect -1995 -18240 -1710 -15390
rect -1995 -18525 1140 -18240
<< locali >>
rect -1995 -7250 -1425 -7125
rect -1995 -7550 -1850 -7250
rect -1550 -7550 -1425 -7250
rect -1995 -7695 -1425 -7550
<< viali >>
rect -1850 -7550 -1550 -7250
<< metal1 >>
rect -1995 -7250 -1425 -7125
rect -1995 -7550 -1850 -7250
rect -1550 -7550 -1425 -7250
rect -1995 -7695 -1425 -7550
<< labels >>
rlabel xpolycontact -1995 570 -1995 570 1 A
rlabel xpolycontact 1425 -18240 1425 -18240 1 B
<< end >>
