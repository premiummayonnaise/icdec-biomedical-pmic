magic
tech sky130A
magscale 1 2
timestamp 1769535502
<< metal3 >>
rect -22328 2512 -16956 2540
rect -22328 -2512 -17040 2512
rect -16976 -2512 -16956 2512
rect -22328 -2540 -16956 -2512
rect -16716 2512 -11344 2540
rect -16716 -2512 -11428 2512
rect -11364 -2512 -11344 2512
rect -16716 -2540 -11344 -2512
rect -11104 2512 -5732 2540
rect -11104 -2512 -5816 2512
rect -5752 -2512 -5732 2512
rect -11104 -2540 -5732 -2512
rect -5492 2512 -120 2540
rect -5492 -2512 -204 2512
rect -140 -2512 -120 2512
rect -5492 -2540 -120 -2512
rect 120 2512 5492 2540
rect 120 -2512 5408 2512
rect 5472 -2512 5492 2512
rect 120 -2540 5492 -2512
rect 5732 2512 11104 2540
rect 5732 -2512 11020 2512
rect 11084 -2512 11104 2512
rect 5732 -2540 11104 -2512
rect 11344 2512 16716 2540
rect 11344 -2512 16632 2512
rect 16696 -2512 16716 2512
rect 11344 -2540 16716 -2512
rect 16956 2512 22328 2540
rect 16956 -2512 22244 2512
rect 22308 -2512 22328 2512
rect 16956 -2540 22328 -2512
<< via3 >>
rect -17040 -2512 -16976 2512
rect -11428 -2512 -11364 2512
rect -5816 -2512 -5752 2512
rect -204 -2512 -140 2512
rect 5408 -2512 5472 2512
rect 11020 -2512 11084 2512
rect 16632 -2512 16696 2512
rect 22244 -2512 22308 2512
<< mimcap >>
rect -22288 2460 -17288 2500
rect -22288 -2460 -22248 2460
rect -17328 -2460 -17288 2460
rect -22288 -2500 -17288 -2460
rect -16676 2460 -11676 2500
rect -16676 -2460 -16636 2460
rect -11716 -2460 -11676 2460
rect -16676 -2500 -11676 -2460
rect -11064 2460 -6064 2500
rect -11064 -2460 -11024 2460
rect -6104 -2460 -6064 2460
rect -11064 -2500 -6064 -2460
rect -5452 2460 -452 2500
rect -5452 -2460 -5412 2460
rect -492 -2460 -452 2460
rect -5452 -2500 -452 -2460
rect 160 2460 5160 2500
rect 160 -2460 200 2460
rect 5120 -2460 5160 2460
rect 160 -2500 5160 -2460
rect 5772 2460 10772 2500
rect 5772 -2460 5812 2460
rect 10732 -2460 10772 2460
rect 5772 -2500 10772 -2460
rect 11384 2460 16384 2500
rect 11384 -2460 11424 2460
rect 16344 -2460 16384 2460
rect 11384 -2500 16384 -2460
rect 16996 2460 21996 2500
rect 16996 -2460 17036 2460
rect 21956 -2460 21996 2460
rect 16996 -2500 21996 -2460
<< mimcapcontact >>
rect -22248 -2460 -17328 2460
rect -16636 -2460 -11716 2460
rect -11024 -2460 -6104 2460
rect -5412 -2460 -492 2460
rect 200 -2460 5120 2460
rect 5812 -2460 10732 2460
rect 11424 -2460 16344 2460
rect 17036 -2460 21956 2460
<< metal4 >>
rect -17056 2512 -16960 2528
rect -22249 2460 -17327 2461
rect -22249 -2460 -22248 2460
rect -17328 -2460 -17327 2460
rect -22249 -2461 -17327 -2460
rect -17056 -2512 -17040 2512
rect -16976 -2512 -16960 2512
rect -11444 2512 -11348 2528
rect -16637 2460 -11715 2461
rect -16637 -2460 -16636 2460
rect -11716 -2460 -11715 2460
rect -16637 -2461 -11715 -2460
rect -17056 -2528 -16960 -2512
rect -11444 -2512 -11428 2512
rect -11364 -2512 -11348 2512
rect -5832 2512 -5736 2528
rect -11025 2460 -6103 2461
rect -11025 -2460 -11024 2460
rect -6104 -2460 -6103 2460
rect -11025 -2461 -6103 -2460
rect -11444 -2528 -11348 -2512
rect -5832 -2512 -5816 2512
rect -5752 -2512 -5736 2512
rect -220 2512 -124 2528
rect -5413 2460 -491 2461
rect -5413 -2460 -5412 2460
rect -492 -2460 -491 2460
rect -5413 -2461 -491 -2460
rect -5832 -2528 -5736 -2512
rect -220 -2512 -204 2512
rect -140 -2512 -124 2512
rect 5392 2512 5488 2528
rect 199 2460 5121 2461
rect 199 -2460 200 2460
rect 5120 -2460 5121 2460
rect 199 -2461 5121 -2460
rect -220 -2528 -124 -2512
rect 5392 -2512 5408 2512
rect 5472 -2512 5488 2512
rect 11004 2512 11100 2528
rect 5811 2460 10733 2461
rect 5811 -2460 5812 2460
rect 10732 -2460 10733 2460
rect 5811 -2461 10733 -2460
rect 5392 -2528 5488 -2512
rect 11004 -2512 11020 2512
rect 11084 -2512 11100 2512
rect 16616 2512 16712 2528
rect 11423 2460 16345 2461
rect 11423 -2460 11424 2460
rect 16344 -2460 16345 2460
rect 11423 -2461 16345 -2460
rect 11004 -2528 11100 -2512
rect 16616 -2512 16632 2512
rect 16696 -2512 16712 2512
rect 22228 2512 22324 2528
rect 17035 2460 21957 2461
rect 17035 -2460 17036 2460
rect 21956 -2460 21957 2460
rect 17035 -2461 21957 -2460
rect 16616 -2528 16712 -2512
rect 22228 -2512 22244 2512
rect 22308 -2512 22324 2512
rect 22228 -2528 22324 -2512
<< properties >>
string FIXED_BBOX 16956 -2540 22036 2540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 25.0 val 1.269k carea 2.00 cperi 0.19 class capacitor nx 8 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
