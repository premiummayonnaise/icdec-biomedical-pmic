magic
tech sky130A
magscale 1 2
timestamp 1769084796
<< mvnmos >>
rect -239 -269 -89 331
rect 89 -269 239 331
<< mvndiff >>
rect -297 319 -239 331
rect -297 -257 -285 319
rect -251 -257 -239 319
rect -297 -269 -239 -257
rect -89 319 -31 331
rect -89 -257 -77 319
rect -43 -257 -31 319
rect -89 -269 -31 -257
rect 31 319 89 331
rect 31 -257 43 319
rect 77 -257 89 319
rect 31 -269 89 -257
rect 239 319 297 331
rect 239 -257 251 319
rect 285 -257 297 319
rect 239 -269 297 -257
<< mvndiffc >>
rect -285 -257 -251 319
rect -77 -257 -43 319
rect 43 -257 77 319
rect 251 -257 285 319
<< poly >>
rect -239 331 -89 357
rect 89 331 239 357
rect -239 -307 -89 -269
rect -239 -341 -223 -307
rect -105 -341 -89 -307
rect -239 -357 -89 -341
rect 89 -307 239 -269
rect 89 -341 105 -307
rect 223 -341 239 -307
rect 89 -357 239 -341
<< polycont >>
rect -223 -341 -105 -307
rect 105 -341 223 -307
<< locali >>
rect -285 319 -251 335
rect -285 -273 -251 -257
rect -77 319 -43 335
rect -77 -273 -43 -257
rect 43 319 77 335
rect 43 -273 77 -257
rect 251 319 285 335
rect 251 -273 285 -257
rect -239 -341 -223 -307
rect -105 -341 -89 -307
rect 89 -341 105 -307
rect 223 -341 239 -307
<< viali >>
rect -285 -257 -251 319
rect -77 -257 -43 319
rect 43 -257 77 319
rect 251 -257 285 319
rect -223 -341 -105 -307
rect 105 -341 223 -307
<< metal1 >>
rect -291 319 -245 331
rect -291 -257 -285 319
rect -251 -257 -245 319
rect -291 -269 -245 -257
rect -83 319 -37 331
rect -83 -257 -77 319
rect -43 -257 -37 319
rect -83 -269 -37 -257
rect 37 319 83 331
rect 37 -257 43 319
rect 77 -257 83 319
rect 37 -269 83 -257
rect 245 319 291 331
rect 245 -257 251 319
rect 285 -257 291 319
rect 245 -269 291 -257
rect -235 -307 -93 -301
rect -235 -341 -223 -307
rect -105 -341 -93 -307
rect -235 -347 -93 -341
rect 93 -307 235 -301
rect 93 -341 105 -307
rect 223 -341 235 -307
rect 93 -347 235 -341
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 0.75 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
