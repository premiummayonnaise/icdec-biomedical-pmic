magic
tech sky130A
magscale 1 2
timestamp 1770117167
<< nwell >>
rect -1061 -672 1061 672
<< mvpmos >>
rect -803 -375 -653 375
rect -595 -375 -445 375
rect -387 -375 -237 375
rect -179 -375 -29 375
rect 29 -375 179 375
rect 237 -375 387 375
rect 445 -375 595 375
rect 653 -375 803 375
<< mvpdiff >>
rect -861 363 -803 375
rect -861 -363 -849 363
rect -815 -363 -803 363
rect -861 -375 -803 -363
rect -653 363 -595 375
rect -653 -363 -641 363
rect -607 -363 -595 363
rect -653 -375 -595 -363
rect -445 363 -387 375
rect -445 -363 -433 363
rect -399 -363 -387 363
rect -445 -375 -387 -363
rect -237 363 -179 375
rect -237 -363 -225 363
rect -191 -363 -179 363
rect -237 -375 -179 -363
rect -29 363 29 375
rect -29 -363 -17 363
rect 17 -363 29 363
rect -29 -375 29 -363
rect 179 363 237 375
rect 179 -363 191 363
rect 225 -363 237 363
rect 179 -375 237 -363
rect 387 363 445 375
rect 387 -363 399 363
rect 433 -363 445 363
rect 387 -375 445 -363
rect 595 363 653 375
rect 595 -363 607 363
rect 641 -363 653 363
rect 595 -375 653 -363
rect 803 363 861 375
rect 803 -363 815 363
rect 849 -363 861 363
rect 803 -375 861 -363
<< mvpdiffc >>
rect -849 -363 -815 363
rect -641 -363 -607 363
rect -433 -363 -399 363
rect -225 -363 -191 363
rect -17 -363 17 363
rect 191 -363 225 363
rect 399 -363 433 363
rect 607 -363 641 363
rect 815 -363 849 363
<< mvnsubdiff >>
rect -995 594 995 606
rect -995 560 -887 594
rect 887 560 995 594
rect -995 548 995 560
rect -995 -548 -937 548
rect 937 -548 995 548
rect -995 -606 995 -548
<< mvnsubdiffcont >>
rect -887 560 887 594
<< poly >>
rect -803 456 -653 472
rect -803 422 -787 456
rect -669 422 -653 456
rect -803 375 -653 422
rect -595 456 -445 472
rect -595 422 -579 456
rect -461 422 -445 456
rect -595 375 -445 422
rect -387 456 -237 472
rect -387 422 -371 456
rect -253 422 -237 456
rect -387 375 -237 422
rect -179 456 -29 472
rect -179 422 -163 456
rect -45 422 -29 456
rect -179 375 -29 422
rect 29 456 179 472
rect 29 422 45 456
rect 163 422 179 456
rect 29 375 179 422
rect 237 456 387 472
rect 237 422 253 456
rect 371 422 387 456
rect 237 375 387 422
rect 445 456 595 472
rect 445 422 461 456
rect 579 422 595 456
rect 445 375 595 422
rect 653 456 803 472
rect 653 422 669 456
rect 787 422 803 456
rect 653 375 803 422
rect -803 -422 -653 -375
rect -803 -456 -787 -422
rect -669 -456 -653 -422
rect -803 -472 -653 -456
rect -595 -422 -445 -375
rect -595 -456 -579 -422
rect -461 -456 -445 -422
rect -595 -472 -445 -456
rect -387 -422 -237 -375
rect -387 -456 -371 -422
rect -253 -456 -237 -422
rect -387 -472 -237 -456
rect -179 -422 -29 -375
rect -179 -456 -163 -422
rect -45 -456 -29 -422
rect -179 -472 -29 -456
rect 29 -422 179 -375
rect 29 -456 45 -422
rect 163 -456 179 -422
rect 29 -472 179 -456
rect 237 -422 387 -375
rect 237 -456 253 -422
rect 371 -456 387 -422
rect 237 -472 387 -456
rect 445 -422 595 -375
rect 445 -456 461 -422
rect 579 -456 595 -422
rect 445 -472 595 -456
rect 653 -422 803 -375
rect 653 -456 669 -422
rect 787 -456 803 -422
rect 653 -472 803 -456
<< polycont >>
rect -787 422 -669 456
rect -579 422 -461 456
rect -371 422 -253 456
rect -163 422 -45 456
rect 45 422 163 456
rect 253 422 371 456
rect 461 422 579 456
rect 669 422 787 456
rect -787 -456 -669 -422
rect -579 -456 -461 -422
rect -371 -456 -253 -422
rect -163 -456 -45 -422
rect 45 -456 163 -422
rect 253 -456 371 -422
rect 461 -456 579 -422
rect 669 -456 787 -422
<< locali >>
rect -983 560 -887 594
rect 887 560 983 594
rect -983 -560 -949 560
rect -803 422 -787 456
rect -669 422 -653 456
rect -595 422 -579 456
rect -461 422 -445 456
rect -387 422 -371 456
rect -253 422 -237 456
rect -179 422 -163 456
rect -45 422 -29 456
rect 29 422 45 456
rect 163 422 179 456
rect 237 422 253 456
rect 371 422 387 456
rect 445 422 461 456
rect 579 422 595 456
rect 653 422 669 456
rect 787 422 803 456
rect -849 363 -815 379
rect -849 -379 -815 -363
rect -641 363 -607 379
rect -641 -379 -607 -363
rect -433 363 -399 379
rect -433 -379 -399 -363
rect -225 363 -191 379
rect -225 -379 -191 -363
rect -17 363 17 379
rect -17 -379 17 -363
rect 191 363 225 379
rect 191 -379 225 -363
rect 399 363 433 379
rect 399 -379 433 -363
rect 607 363 641 379
rect 607 -379 641 -363
rect 815 363 849 379
rect 815 -379 849 -363
rect -803 -456 -787 -422
rect -669 -456 -653 -422
rect -595 -456 -579 -422
rect -461 -456 -445 -422
rect -387 -456 -371 -422
rect -253 -456 -237 -422
rect -179 -456 -163 -422
rect -45 -456 -29 -422
rect 29 -456 45 -422
rect 163 -456 179 -422
rect 237 -456 253 -422
rect 371 -456 387 -422
rect 445 -456 461 -422
rect 579 -456 595 -422
rect 653 -456 669 -422
rect 787 -456 803 -422
rect 949 -560 983 560
rect -983 -594 983 -560
<< viali >>
rect -787 422 -669 456
rect -579 422 -461 456
rect -371 422 -253 456
rect -163 422 -45 456
rect 45 422 163 456
rect 253 422 371 456
rect 461 422 579 456
rect 669 422 787 456
rect -849 -363 -815 363
rect -641 -363 -607 363
rect -433 -363 -399 363
rect -225 -363 -191 363
rect -17 -363 17 363
rect 191 -363 225 363
rect 399 -363 433 363
rect 607 -363 641 363
rect 815 -363 849 363
rect -787 -456 -669 -422
rect -579 -456 -461 -422
rect -371 -456 -253 -422
rect -163 -456 -45 -422
rect 45 -456 163 -422
rect 253 -456 371 -422
rect 461 -456 579 -422
rect 669 -456 787 -422
<< metal1 >>
rect -799 456 -657 462
rect -799 422 -787 456
rect -669 422 -657 456
rect -799 416 -657 422
rect -591 456 -449 462
rect -591 422 -579 456
rect -461 422 -449 456
rect -591 416 -449 422
rect -383 456 -241 462
rect -383 422 -371 456
rect -253 422 -241 456
rect -383 416 -241 422
rect -175 456 -33 462
rect -175 422 -163 456
rect -45 422 -33 456
rect -175 416 -33 422
rect 33 456 175 462
rect 33 422 45 456
rect 163 422 175 456
rect 33 416 175 422
rect 241 456 383 462
rect 241 422 253 456
rect 371 422 383 456
rect 241 416 383 422
rect 449 456 591 462
rect 449 422 461 456
rect 579 422 591 456
rect 449 416 591 422
rect 657 456 799 462
rect 657 422 669 456
rect 787 422 799 456
rect 657 416 799 422
rect -855 363 -809 375
rect -855 -363 -849 363
rect -815 -363 -809 363
rect -855 -375 -809 -363
rect -647 363 -601 375
rect -647 -363 -641 363
rect -607 -363 -601 363
rect -647 -375 -601 -363
rect -439 363 -393 375
rect -439 -363 -433 363
rect -399 -363 -393 363
rect -439 -375 -393 -363
rect -231 363 -185 375
rect -231 -363 -225 363
rect -191 -363 -185 363
rect -231 -375 -185 -363
rect -23 363 23 375
rect -23 -363 -17 363
rect 17 -363 23 363
rect -23 -375 23 -363
rect 185 363 231 375
rect 185 -363 191 363
rect 225 -363 231 363
rect 185 -375 231 -363
rect 393 363 439 375
rect 393 -363 399 363
rect 433 -363 439 363
rect 393 -375 439 -363
rect 601 363 647 375
rect 601 -363 607 363
rect 641 -363 647 363
rect 601 -375 647 -363
rect 809 363 855 375
rect 809 -363 815 363
rect 849 -363 855 363
rect 809 -375 855 -363
rect -799 -422 -657 -416
rect -799 -456 -787 -422
rect -669 -456 -657 -422
rect -799 -462 -657 -456
rect -591 -422 -449 -416
rect -591 -456 -579 -422
rect -461 -456 -449 -422
rect -591 -462 -449 -456
rect -383 -422 -241 -416
rect -383 -456 -371 -422
rect -253 -456 -241 -422
rect -383 -462 -241 -456
rect -175 -422 -33 -416
rect -175 -456 -163 -422
rect -45 -456 -33 -422
rect -175 -462 -33 -456
rect 33 -422 175 -416
rect 33 -456 45 -422
rect 163 -456 175 -422
rect 33 -462 175 -456
rect 241 -422 383 -416
rect 241 -456 253 -422
rect 371 -456 383 -422
rect 241 -462 383 -456
rect 449 -422 591 -416
rect 449 -456 461 -422
rect 579 -456 591 -422
rect 449 -462 591 -456
rect 657 -422 799 -416
rect 657 -456 669 -422
rect 787 -456 799 -422
rect 657 -462 799 -456
<< labels >>
rlabel mvnsubdiff 0 -577 0 -577 0 B
port 1 nsew
rlabel mvpdiffc -832 0 -832 0 0 D0
port 2 nsew
rlabel polycont -728 439 -728 439 0 G0
port 3 nsew
rlabel mvpdiffc -624 0 -624 0 0 S1
port 4 nsew
rlabel polycont -520 439 -520 439 0 G1
port 5 nsew
rlabel mvpdiffc -416 0 -416 0 0 D2
port 6 nsew
rlabel polycont -312 439 -312 439 0 G2
port 7 nsew
rlabel mvpdiffc -208 0 -208 0 0 S3
port 8 nsew
rlabel polycont -104 439 -104 439 0 G3
port 9 nsew
rlabel mvpdiffc 0 0 0 0 0 D4
port 10 nsew
rlabel polycont 104 439 104 439 0 G4
port 11 nsew
rlabel mvpdiffc 208 0 208 0 0 S5
port 12 nsew
rlabel polycont 312 439 312 439 0 G5
port 13 nsew
rlabel mvpdiffc 416 0 416 0 0 D6
port 14 nsew
rlabel polycont 520 439 520 439 0 G6
port 15 nsew
rlabel mvpdiffc 624 0 624 0 0 S7
port 16 nsew
rlabel polycont 728 439 728 439 0 G7
port 17 nsew
<< properties >>
string FIXED_BBOX -966 -577 966 577
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3.75 l 0.75 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
