magic
tech sky130A
magscale 1 2
timestamp 1770370310
<< nwell >>
rect 9900 -560 16900 420
rect 6760 -3560 20040 -560
rect 6760 -5300 9260 -3560
rect 6760 -9160 7040 -5300
rect 17540 -5300 20040 -3560
rect 19760 -9160 20040 -5300
rect 6760 -9440 10140 -9160
rect 9860 -10160 10140 -9440
rect 16620 -9440 20040 -9160
rect 16620 -10160 16900 -9440
rect 9860 -10440 16900 -10160
<< pwell >>
rect 9300 -5340 17500 -3600
rect 7060 -5360 19760 -5340
rect 7060 -7660 19740 -5360
rect 7060 -7680 17640 -7660
rect 18820 -7680 19740 -7660
rect 7060 -9140 19740 -7680
rect 10140 -10160 16620 -9160
<< psubdiff >>
rect 9500 -3720 17300 -3700
rect 9500 -3780 9620 -3720
rect 17180 -3780 17300 -3720
rect 9500 -3800 17300 -3780
rect 9500 -3820 9600 -3800
rect 7720 -5540 9420 -5520
rect 7720 -5600 7840 -5540
rect 9300 -5600 9420 -5540
rect 7720 -5620 9420 -5600
rect 7720 -5640 7820 -5620
rect 7720 -7400 7740 -5640
rect 7800 -7400 7820 -5640
rect 9320 -5640 9420 -5620
rect 7720 -7420 7820 -7400
rect 9320 -7400 9340 -5640
rect 9400 -7400 9420 -5640
rect 9500 -7080 9520 -3820
rect 9580 -7080 9600 -3820
rect 17200 -3820 17300 -3800
rect 9700 -3920 11300 -3900
rect 9700 -3980 9740 -3920
rect 11260 -3980 11300 -3920
rect 9700 -4000 11300 -3980
rect 9700 -5200 9800 -4000
rect 11200 -5200 11300 -4000
rect 9700 -5300 11300 -5200
rect 11500 -3920 13100 -3900
rect 11500 -3980 11540 -3920
rect 13060 -3980 13100 -3920
rect 11500 -4000 13100 -3980
rect 11500 -5200 11600 -4000
rect 13000 -5200 13100 -4000
rect 11500 -5300 13100 -5200
rect 13700 -3920 15300 -3900
rect 13700 -3980 13740 -3920
rect 15260 -3980 15300 -3920
rect 13700 -4000 15300 -3980
rect 13700 -5200 13800 -4000
rect 15200 -5200 15300 -4000
rect 13700 -5300 15300 -5200
rect 15500 -3920 17100 -3900
rect 15500 -3980 15540 -3920
rect 17060 -3980 17100 -3920
rect 15500 -4000 17100 -3980
rect 15500 -5200 15600 -4000
rect 17000 -5200 17100 -4000
rect 15500 -5300 17100 -5200
rect 9700 -5700 11300 -5600
rect 9700 -6900 9800 -5700
rect 11200 -6900 11300 -5700
rect 9700 -6920 11300 -6900
rect 9700 -6980 9740 -6920
rect 11260 -6980 11300 -6920
rect 9700 -7000 11300 -6980
rect 11500 -5700 13100 -5600
rect 11500 -6900 11600 -5700
rect 13000 -6900 13100 -5700
rect 11500 -6920 13100 -6900
rect 11500 -6980 11540 -6920
rect 13060 -6980 13100 -6920
rect 11500 -7000 13100 -6980
rect 13700 -5700 15300 -5600
rect 13700 -6900 13800 -5700
rect 15200 -6900 15300 -5700
rect 13700 -6920 15300 -6900
rect 13700 -6980 13740 -6920
rect 15260 -6980 15300 -6920
rect 13700 -7000 15300 -6980
rect 15500 -5700 17100 -5600
rect 15500 -6900 15600 -5700
rect 17000 -6900 17100 -5700
rect 15500 -6920 17100 -6900
rect 15500 -6980 15540 -6920
rect 17060 -6980 17100 -6920
rect 15500 -7000 17100 -6980
rect 9500 -7100 9600 -7080
rect 17200 -7080 17220 -3820
rect 17280 -7080 17300 -3820
rect 17200 -7100 17300 -7080
rect 9500 -7120 17300 -7100
rect 9500 -7180 9620 -7120
rect 17180 -7180 17300 -7120
rect 9500 -7200 17300 -7180
rect 17380 -5560 19080 -5540
rect 17380 -5620 17500 -5560
rect 18960 -5620 19080 -5560
rect 17380 -5640 19080 -5620
rect 17380 -5660 17480 -5640
rect 9320 -7420 9420 -7400
rect 7720 -7440 9420 -7420
rect 7720 -7500 7840 -7440
rect 9300 -7500 9420 -7440
rect 7720 -7520 9420 -7500
rect 10200 -7220 10300 -7200
rect 10200 -8980 10220 -7220
rect 10280 -8980 10300 -7220
rect 10200 -9000 10300 -8980
rect 16400 -7220 16500 -7200
rect 16400 -8980 16420 -7220
rect 16480 -8980 16500 -7220
rect 17380 -7400 17400 -5660
rect 17460 -7400 17480 -5660
rect 18980 -5660 19080 -5640
rect 17380 -7420 17480 -7400
rect 18980 -7400 19000 -5660
rect 19060 -7400 19080 -5660
rect 18980 -7420 19080 -7400
rect 17380 -7440 19080 -7420
rect 17380 -7500 17500 -7440
rect 18960 -7500 19080 -7440
rect 17380 -7520 19080 -7500
rect 16400 -9000 16500 -8980
rect 10200 -9020 16500 -9000
rect 10200 -9080 10320 -9020
rect 16380 -9080 16500 -9020
rect 10200 -9100 16500 -9080
<< nsubdiff >>
rect 9940 360 16860 380
rect 9940 -600 9980 360
rect 6800 -620 9980 -600
rect 6800 -780 7000 -620
rect 9920 -780 9980 -620
rect 10100 200 10140 360
rect 16660 200 16700 360
rect 10100 180 16700 200
rect 10100 -780 10140 180
rect 6800 -800 10140 -780
rect 10240 -640 16540 -620
rect 10240 -700 10360 -640
rect 16420 -700 16540 -640
rect 10240 -720 16540 -700
rect 10240 -740 10340 -720
rect 6800 -820 7000 -800
rect 6800 -9180 6820 -820
rect 6980 -9180 7000 -820
rect 7240 -1020 10140 -1000
rect 7240 -1080 7360 -1020
rect 10020 -1080 10140 -1020
rect 7240 -1100 10140 -1080
rect 7240 -1120 7340 -1100
rect 7240 -3380 7260 -1120
rect 7320 -3380 7340 -1120
rect 10040 -1120 10140 -1100
rect 7240 -3400 7340 -3380
rect 10040 -3380 10060 -1120
rect 10120 -3380 10140 -1120
rect 10240 -2900 10260 -740
rect 10320 -2900 10340 -740
rect 10240 -2920 10340 -2900
rect 16440 -740 16540 -720
rect 16440 -2900 16460 -740
rect 16520 -2900 16540 -740
rect 16660 -780 16700 180
rect 16820 -600 16860 360
rect 16820 -620 20000 -600
rect 16820 -780 16860 -620
rect 19780 -780 20000 -620
rect 16660 -800 20000 -780
rect 19800 -820 20000 -800
rect 16440 -2920 16540 -2900
rect 10240 -2940 16540 -2920
rect 10240 -3000 10360 -2940
rect 16420 -3000 16540 -2940
rect 10240 -3020 16540 -3000
rect 16640 -1020 19540 -1000
rect 16640 -1080 16760 -1020
rect 19420 -1080 19540 -1020
rect 16640 -1100 19540 -1080
rect 16640 -1120 16740 -1100
rect 10040 -3400 10140 -3380
rect 7240 -3420 10140 -3400
rect 7240 -3480 7360 -3420
rect 10020 -3480 10140 -3420
rect 7240 -3500 10140 -3480
rect 16640 -3380 16660 -1120
rect 16720 -3380 16740 -1120
rect 19440 -1120 19540 -1100
rect 16640 -3400 16740 -3380
rect 19440 -3380 19460 -1120
rect 19520 -3380 19540 -1120
rect 19440 -3400 19540 -3380
rect 16640 -3420 19540 -3400
rect 16640 -3480 16760 -3420
rect 19420 -3480 19540 -3420
rect 16640 -3500 19540 -3480
rect 8100 -3720 9100 -3700
rect 8100 -3780 8220 -3720
rect 8980 -3780 9100 -3720
rect 8100 -3800 9100 -3780
rect 8100 -3820 8200 -3800
rect 8100 -5080 8120 -3820
rect 8180 -5080 8200 -3820
rect 9000 -3820 9100 -3800
rect 8100 -5100 8200 -5080
rect 9000 -5080 9020 -3820
rect 9080 -5080 9100 -3820
rect 9000 -5100 9100 -5080
rect 8100 -5120 9100 -5100
rect 8100 -5180 8220 -5120
rect 8980 -5180 9100 -5120
rect 8100 -5200 9100 -5180
rect 17700 -3720 18700 -3700
rect 17700 -3780 17820 -3720
rect 18580 -3780 18700 -3720
rect 17700 -3800 18700 -3780
rect 17700 -3820 17800 -3800
rect 17700 -5080 17720 -3820
rect 17780 -5080 17800 -3820
rect 18600 -3820 18700 -3800
rect 17700 -5100 17800 -5080
rect 18600 -5080 18620 -3820
rect 18680 -5080 18700 -3820
rect 18600 -5100 18700 -5080
rect 17700 -5120 18700 -5100
rect 17700 -5180 17820 -5120
rect 18580 -5180 18700 -5120
rect 17700 -5200 18700 -5180
rect 6800 -9200 7000 -9180
rect 19800 -9180 19820 -820
rect 19980 -9180 20000 -820
rect 19800 -9200 20000 -9180
rect 6800 -9220 10100 -9200
rect 6800 -9380 7020 -9220
rect 9880 -9380 9940 -9220
rect 6800 -9400 9940 -9380
rect 9900 -10380 9940 -9400
rect 10060 -10200 10100 -9220
rect 16660 -9220 20000 -9200
rect 16660 -10200 16700 -9220
rect 10060 -10220 16700 -10200
rect 10060 -10380 10100 -10220
rect 16660 -10380 16700 -10220
rect 16820 -9380 16860 -9220
rect 19780 -9380 20000 -9220
rect 16820 -9400 20000 -9380
rect 16820 -10380 16860 -9400
rect 9900 -10400 16860 -10380
<< psubdiffcont >>
rect 9620 -3780 17180 -3720
rect 7840 -5600 9300 -5540
rect 7740 -7400 7800 -5640
rect 9340 -7400 9400 -5640
rect 9520 -7080 9580 -3820
rect 9740 -3980 11260 -3920
rect 11540 -3980 13060 -3920
rect 13740 -3980 15260 -3920
rect 15540 -3980 17060 -3920
rect 9740 -6980 11260 -6920
rect 11540 -6980 13060 -6920
rect 13740 -6980 15260 -6920
rect 15540 -6980 17060 -6920
rect 17220 -7080 17280 -3820
rect 9620 -7180 17180 -7120
rect 17500 -5620 18960 -5560
rect 7840 -7500 9300 -7440
rect 10220 -8980 10280 -7220
rect 16420 -8980 16480 -7220
rect 17400 -7400 17460 -5660
rect 19000 -7400 19060 -5660
rect 17500 -7500 18960 -7440
rect 10320 -9080 16380 -9020
<< nsubdiffcont >>
rect 7000 -780 9920 -620
rect 9980 -780 10100 360
rect 10140 200 16660 360
rect 10360 -700 16420 -640
rect 6820 -9180 6980 -820
rect 7360 -1080 10020 -1020
rect 7260 -3380 7320 -1120
rect 10060 -3380 10120 -1120
rect 10260 -2900 10320 -740
rect 16460 -2900 16520 -740
rect 16700 -780 16820 360
rect 16860 -780 19780 -620
rect 10360 -3000 16420 -2940
rect 16760 -1080 19420 -1020
rect 7360 -3480 10020 -3420
rect 16660 -3380 16720 -1120
rect 19460 -3380 19520 -1120
rect 16760 -3480 19420 -3420
rect 8220 -3780 8980 -3720
rect 8120 -5080 8180 -3820
rect 9020 -5080 9080 -3820
rect 8220 -5180 8980 -5120
rect 17820 -3780 18580 -3720
rect 17720 -5080 17780 -3820
rect 18620 -5080 18680 -3820
rect 17820 -5180 18580 -5120
rect 19820 -9180 19980 -820
rect 7020 -9380 9880 -9220
rect 9940 -10380 10060 -9220
rect 10100 -10380 16660 -10220
rect 16700 -10380 16820 -9220
rect 16860 -9380 19780 -9220
<< poly >>
rect 7360 -3320 7390 -1150
rect 9950 -3320 9980 -1150
rect 16800 -3320 16830 -1160
rect 19390 -3320 19420 -1160
rect 8320 -5020 8350 -3870
rect 8920 -5020 8950 -3870
rect 7840 -7320 7900 -5700
rect 9230 -7320 9290 -5700
rect 17900 -4990 17930 -3840
rect 18500 -4990 18530 -3840
rect 17500 -7340 17560 -5720
rect 18890 -7340 18950 -5720
<< locali >>
rect 9940 360 16860 380
rect 9940 -600 9980 360
rect 6800 -620 9980 -600
rect 6800 -780 7000 -620
rect 9920 -780 9980 -620
rect 10100 200 10140 360
rect 16660 200 16700 360
rect 10100 100 16700 200
rect 10100 20 10160 100
rect 10240 20 10280 100
rect 10360 20 10400 100
rect 10480 20 10520 100
rect 10600 20 10640 100
rect 10720 20 10760 100
rect 10840 20 10880 100
rect 10960 20 11000 100
rect 11080 20 11120 100
rect 11200 20 11240 100
rect 11320 20 11360 100
rect 11440 20 11480 100
rect 11560 20 11600 100
rect 11680 20 11720 100
rect 11800 20 11840 100
rect 11920 20 11960 100
rect 12040 20 12080 100
rect 12160 20 12200 100
rect 12280 20 12320 100
rect 12400 20 12440 100
rect 12520 20 12560 100
rect 12640 20 12680 100
rect 12760 20 12800 100
rect 12880 20 12920 100
rect 13000 20 13040 100
rect 13120 20 13160 100
rect 13240 20 13280 100
rect 13360 20 13400 100
rect 13480 20 13520 100
rect 13600 20 13640 100
rect 13720 20 13760 100
rect 13840 20 13880 100
rect 13960 20 14000 100
rect 14080 20 14120 100
rect 14200 20 14240 100
rect 14320 20 14360 100
rect 14440 20 14480 100
rect 14560 20 14600 100
rect 14680 20 14720 100
rect 14800 20 14840 100
rect 14920 20 14960 100
rect 15040 20 15080 100
rect 15160 20 15200 100
rect 15280 20 15320 100
rect 15400 20 15440 100
rect 15520 20 15560 100
rect 15640 20 15680 100
rect 15760 20 15800 100
rect 15880 20 15920 100
rect 16000 20 16040 100
rect 16120 20 16160 100
rect 16240 20 16280 100
rect 16360 20 16400 100
rect 16480 20 16520 100
rect 16600 20 16700 100
rect 10100 -20 16700 20
rect 10100 -100 10160 -20
rect 10240 -100 10280 -20
rect 10360 -100 10400 -20
rect 10480 -100 10520 -20
rect 10600 -100 10640 -20
rect 10720 -100 10760 -20
rect 10840 -100 10880 -20
rect 10960 -100 11000 -20
rect 11080 -100 11120 -20
rect 11200 -100 11240 -20
rect 11320 -100 11360 -20
rect 11440 -100 11480 -20
rect 11560 -100 11600 -20
rect 11680 -100 11720 -20
rect 11800 -100 11840 -20
rect 11920 -100 11960 -20
rect 12040 -100 12080 -20
rect 12160 -100 12200 -20
rect 12280 -100 12320 -20
rect 12400 -100 12440 -20
rect 12520 -100 12560 -20
rect 12640 -100 12680 -20
rect 12760 -100 12800 -20
rect 12880 -100 12920 -20
rect 13000 -100 13040 -20
rect 13120 -100 13160 -20
rect 13240 -100 13280 -20
rect 13360 -100 13400 -20
rect 13480 -100 13520 -20
rect 13600 -100 13640 -20
rect 13720 -100 13760 -20
rect 13840 -100 13880 -20
rect 13960 -100 14000 -20
rect 14080 -100 14120 -20
rect 14200 -100 14240 -20
rect 14320 -100 14360 -20
rect 14440 -100 14480 -20
rect 14560 -100 14600 -20
rect 14680 -100 14720 -20
rect 14800 -100 14840 -20
rect 14920 -100 14960 -20
rect 15040 -100 15080 -20
rect 15160 -100 15200 -20
rect 15280 -100 15320 -20
rect 15400 -100 15440 -20
rect 15520 -100 15560 -20
rect 15640 -100 15680 -20
rect 15760 -100 15800 -20
rect 15880 -100 15920 -20
rect 16000 -100 16040 -20
rect 16120 -100 16160 -20
rect 16240 -100 16280 -20
rect 16360 -100 16400 -20
rect 16480 -100 16520 -20
rect 16600 -100 16700 -20
rect 10100 -140 16700 -100
rect 10100 -220 10160 -140
rect 10240 -220 10280 -140
rect 10360 -220 10400 -140
rect 10480 -220 10520 -140
rect 10600 -220 10640 -140
rect 10720 -220 10760 -140
rect 10840 -220 10880 -140
rect 10960 -220 11000 -140
rect 11080 -220 11120 -140
rect 11200 -220 11240 -140
rect 11320 -220 11360 -140
rect 11440 -220 11480 -140
rect 11560 -220 11600 -140
rect 11680 -220 11720 -140
rect 11800 -220 11840 -140
rect 11920 -220 11960 -140
rect 12040 -220 12080 -140
rect 12160 -220 12200 -140
rect 12280 -220 12320 -140
rect 12400 -220 12440 -140
rect 12520 -220 12560 -140
rect 12640 -220 12680 -140
rect 12760 -220 12800 -140
rect 12880 -220 12920 -140
rect 13000 -220 13040 -140
rect 13120 -220 13160 -140
rect 13240 -220 13280 -140
rect 13360 -220 13400 -140
rect 13480 -220 13520 -140
rect 13600 -220 13640 -140
rect 13720 -220 13760 -140
rect 13840 -220 13880 -140
rect 13960 -220 14000 -140
rect 14080 -220 14120 -140
rect 14200 -220 14240 -140
rect 14320 -220 14360 -140
rect 14440 -220 14480 -140
rect 14560 -220 14600 -140
rect 14680 -220 14720 -140
rect 14800 -220 14840 -140
rect 14920 -220 14960 -140
rect 15040 -220 15080 -140
rect 15160 -220 15200 -140
rect 15280 -220 15320 -140
rect 15400 -220 15440 -140
rect 15520 -220 15560 -140
rect 15640 -220 15680 -140
rect 15760 -220 15800 -140
rect 15880 -220 15920 -140
rect 16000 -220 16040 -140
rect 16120 -220 16160 -140
rect 16240 -220 16280 -140
rect 16360 -220 16400 -140
rect 16480 -220 16520 -140
rect 16600 -220 16700 -140
rect 10100 -260 16700 -220
rect 10100 -340 10160 -260
rect 10240 -340 10280 -260
rect 10360 -340 10400 -260
rect 10480 -340 10520 -260
rect 10600 -340 10640 -260
rect 10720 -340 10760 -260
rect 10840 -340 10880 -260
rect 10960 -340 11000 -260
rect 11080 -340 11120 -260
rect 11200 -340 11240 -260
rect 11320 -340 11360 -260
rect 11440 -340 11480 -260
rect 11560 -340 11600 -260
rect 11680 -340 11720 -260
rect 11800 -340 11840 -260
rect 11920 -340 11960 -260
rect 12040 -340 12080 -260
rect 12160 -340 12200 -260
rect 12280 -340 12320 -260
rect 12400 -340 12440 -260
rect 12520 -340 12560 -260
rect 12640 -340 12680 -260
rect 12760 -340 12800 -260
rect 12880 -340 12920 -260
rect 13000 -340 13040 -260
rect 13120 -340 13160 -260
rect 13240 -340 13280 -260
rect 13360 -340 13400 -260
rect 13480 -340 13520 -260
rect 13600 -340 13640 -260
rect 13720 -340 13760 -260
rect 13840 -340 13880 -260
rect 13960 -340 14000 -260
rect 14080 -340 14120 -260
rect 14200 -340 14240 -260
rect 14320 -340 14360 -260
rect 14440 -340 14480 -260
rect 14560 -340 14600 -260
rect 14680 -340 14720 -260
rect 14800 -340 14840 -260
rect 14920 -340 14960 -260
rect 15040 -340 15080 -260
rect 15160 -340 15200 -260
rect 15280 -340 15320 -260
rect 15400 -340 15440 -260
rect 15520 -340 15560 -260
rect 15640 -340 15680 -260
rect 15760 -340 15800 -260
rect 15880 -340 15920 -260
rect 16000 -340 16040 -260
rect 16120 -340 16160 -260
rect 16240 -340 16280 -260
rect 16360 -340 16400 -260
rect 16480 -340 16520 -260
rect 16600 -340 16700 -260
rect 10100 -380 16700 -340
rect 10100 -460 10160 -380
rect 10240 -460 10280 -380
rect 10360 -460 10400 -380
rect 10480 -460 10520 -380
rect 10600 -460 10640 -380
rect 10720 -460 10760 -380
rect 10840 -460 10880 -380
rect 10960 -460 11000 -380
rect 11080 -460 11120 -380
rect 11200 -460 11240 -380
rect 11320 -460 11360 -380
rect 11440 -460 11480 -380
rect 11560 -460 11600 -380
rect 11680 -460 11720 -380
rect 11800 -460 11840 -380
rect 11920 -460 11960 -380
rect 12040 -460 12080 -380
rect 12160 -460 12200 -380
rect 12280 -460 12320 -380
rect 12400 -460 12440 -380
rect 12520 -460 12560 -380
rect 12640 -460 12680 -380
rect 12760 -460 12800 -380
rect 12880 -460 12920 -380
rect 13000 -460 13040 -380
rect 13120 -460 13160 -380
rect 13240 -460 13280 -380
rect 13360 -460 13400 -380
rect 13480 -460 13520 -380
rect 13600 -460 13640 -380
rect 13720 -460 13760 -380
rect 13840 -460 13880 -380
rect 13960 -460 14000 -380
rect 14080 -460 14120 -380
rect 14200 -460 14240 -380
rect 14320 -460 14360 -380
rect 14440 -460 14480 -380
rect 14560 -460 14600 -380
rect 14680 -460 14720 -380
rect 14800 -460 14840 -380
rect 14920 -460 14960 -380
rect 15040 -460 15080 -380
rect 15160 -460 15200 -380
rect 15280 -460 15320 -380
rect 15400 -460 15440 -380
rect 15520 -460 15560 -380
rect 15640 -460 15680 -380
rect 15760 -460 15800 -380
rect 15880 -460 15920 -380
rect 16000 -460 16040 -380
rect 16120 -460 16160 -380
rect 16240 -460 16280 -380
rect 16360 -460 16400 -380
rect 16480 -460 16520 -380
rect 16600 -460 16700 -380
rect 10100 -500 16700 -460
rect 10100 -580 10160 -500
rect 10240 -580 10280 -500
rect 10360 -580 10400 -500
rect 10480 -580 10520 -500
rect 10600 -580 10640 -500
rect 10720 -580 10760 -500
rect 10840 -580 10880 -500
rect 10960 -580 11000 -500
rect 11080 -580 11120 -500
rect 11200 -580 11240 -500
rect 11320 -580 11360 -500
rect 11440 -580 11480 -500
rect 11560 -580 11600 -500
rect 11680 -580 11720 -500
rect 11800 -580 11840 -500
rect 11920 -580 11960 -500
rect 12040 -580 12080 -500
rect 12160 -580 12200 -500
rect 12280 -580 12320 -500
rect 12400 -580 12440 -500
rect 12520 -580 12560 -500
rect 12640 -580 12680 -500
rect 12760 -580 12800 -500
rect 12880 -580 12920 -500
rect 13000 -580 13040 -500
rect 13120 -580 13160 -500
rect 13240 -580 13280 -500
rect 13360 -580 13400 -500
rect 13480 -580 13520 -500
rect 13600 -580 13640 -500
rect 13720 -580 13760 -500
rect 13840 -580 13880 -500
rect 13960 -580 14000 -500
rect 14080 -580 14120 -500
rect 14200 -580 14240 -500
rect 14320 -580 14360 -500
rect 14440 -580 14480 -500
rect 14560 -580 14600 -500
rect 14680 -580 14720 -500
rect 14800 -580 14840 -500
rect 14920 -580 14960 -500
rect 15040 -580 15080 -500
rect 15160 -580 15200 -500
rect 15280 -580 15320 -500
rect 15400 -580 15440 -500
rect 15520 -580 15560 -500
rect 15640 -580 15680 -500
rect 15760 -580 15800 -500
rect 15880 -580 15920 -500
rect 16000 -580 16040 -500
rect 16120 -580 16160 -500
rect 16240 -580 16280 -500
rect 16360 -580 16400 -500
rect 16480 -580 16520 -500
rect 16600 -580 16700 -500
rect 10100 -640 16700 -580
rect 10100 -700 10360 -640
rect 16420 -700 16700 -640
rect 10100 -720 16700 -700
rect 10100 -740 10340 -720
rect 10100 -780 10260 -740
rect 6800 -820 10260 -780
rect 6800 -9180 6820 -820
rect 6980 -1020 10260 -820
rect 6980 -1080 7360 -1020
rect 10020 -1080 10260 -1020
rect 6980 -1100 10260 -1080
rect 6980 -1120 7340 -1100
rect 6980 -3380 7260 -1120
rect 7320 -3380 7340 -1120
rect 7660 -3200 7820 -1100
rect 8280 -3200 8440 -1100
rect 8880 -3200 9040 -1100
rect 9500 -3200 9660 -1100
rect 10040 -1120 10260 -1100
rect 6980 -3400 7340 -3380
rect 10040 -3380 10060 -1120
rect 10120 -2900 10260 -1120
rect 10320 -2900 10340 -740
rect 10420 -2760 10480 -720
rect 10580 -2760 10640 -720
rect 10740 -2760 10800 -720
rect 10420 -2820 10800 -2760
rect 10860 -2760 11000 -840
rect 11100 -2620 11240 -720
rect 11720 -2620 11860 -720
rect 12020 -2760 12160 -840
rect 12340 -2620 12480 -720
rect 12960 -2620 13100 -720
rect 13260 -2760 13400 -840
rect 13580 -2620 13720 -720
rect 14180 -2600 14320 -720
rect 14480 -2760 14620 -840
rect 14800 -2600 14940 -720
rect 15420 -2600 15560 -720
rect 15720 -2760 15860 -840
rect 10860 -2820 15860 -2760
rect 15920 -2760 15980 -720
rect 16080 -2760 16140 -720
rect 16240 -2760 16300 -720
rect 15920 -2820 16300 -2760
rect 16440 -740 16700 -720
rect 10120 -2920 10340 -2900
rect 16440 -2900 16460 -740
rect 16520 -780 16700 -740
rect 16820 -600 16860 360
rect 16820 -620 20000 -600
rect 16820 -780 16860 -620
rect 19780 -780 20000 -620
rect 16520 -820 20000 -780
rect 16520 -1020 19820 -820
rect 16520 -1080 16760 -1020
rect 19420 -1080 19820 -1020
rect 16520 -1100 19820 -1080
rect 16520 -1120 16740 -1100
rect 16520 -2900 16660 -1120
rect 16440 -2920 16660 -2900
rect 10120 -2940 16660 -2920
rect 10120 -3000 10360 -2940
rect 16420 -3000 16660 -2940
rect 10120 -3380 16660 -3000
rect 16720 -3380 16740 -1120
rect 17120 -3200 17280 -1100
rect 17720 -3200 17880 -1100
rect 18340 -3200 18500 -1100
rect 18940 -3200 19100 -1100
rect 19440 -1120 19820 -1100
rect 10040 -3400 16740 -3380
rect 19440 -3380 19460 -1120
rect 19520 -3380 19820 -1120
rect 19440 -3400 19820 -3380
rect 6980 -3420 19820 -3400
rect 6980 -3480 7360 -3420
rect 10020 -3480 16760 -3420
rect 19420 -3480 19820 -3420
rect 6980 -3560 19820 -3480
rect 6980 -3720 9260 -3560
rect 6980 -3780 8220 -3720
rect 8980 -3780 9260 -3720
rect 6980 -3800 9260 -3780
rect 6980 -3820 8200 -3800
rect 6980 -5080 8120 -3820
rect 8180 -5080 8200 -3820
rect 6980 -5100 8200 -5080
rect 9000 -3820 9260 -3800
rect 9000 -5080 9020 -3820
rect 9080 -5080 9260 -3820
rect 9000 -5100 9260 -5080
rect 6980 -5120 9260 -5100
rect 6980 -5180 8220 -5120
rect 8980 -5180 9260 -5120
rect 6980 -5300 9260 -5180
rect 9300 -3720 17500 -3600
rect 9300 -3780 9620 -3720
rect 17180 -3780 17500 -3720
rect 9300 -3800 17500 -3780
rect 9300 -3820 13100 -3800
rect 6980 -9180 7000 -5300
rect 9300 -5340 9520 -3820
rect 7040 -5380 9520 -5340
rect 7040 -5460 8440 -5380
rect 8520 -5460 8580 -5380
rect 8680 -5460 8740 -5380
rect 8820 -5460 9520 -5380
rect 7040 -5540 9520 -5460
rect 7040 -5600 7840 -5540
rect 9300 -5600 9520 -5540
rect 7040 -5620 9520 -5600
rect 7040 -5640 7820 -5620
rect 7040 -7400 7740 -5640
rect 7800 -7400 7820 -5640
rect 8180 -7220 8340 -5620
rect 8800 -7220 8960 -5620
rect 9320 -5640 9520 -5620
rect 7040 -7420 7820 -7400
rect 9320 -7400 9340 -5640
rect 9400 -7080 9520 -5640
rect 9580 -3920 13100 -3820
rect 13700 -3820 17500 -3800
rect 9580 -3980 9740 -3920
rect 11260 -3980 11540 -3920
rect 13060 -3980 13100 -3920
rect 9580 -4000 13100 -3980
rect 13140 -3900 13660 -3840
rect 13140 -3980 13220 -3900
rect 13300 -3980 13360 -3900
rect 13440 -3980 13500 -3900
rect 13580 -3980 13660 -3900
rect 9580 -6900 9660 -4000
rect 9860 -5080 9920 -4000
rect 10020 -5080 10080 -4000
rect 10180 -5080 10240 -4000
rect 9860 -5160 10240 -5080
rect 10740 -5080 10800 -4000
rect 10900 -5080 10960 -4000
rect 11060 -5080 11120 -4000
rect 10740 -5160 11120 -5080
rect 11300 -4060 11500 -4040
rect 11300 -4140 11360 -4060
rect 11440 -4140 11500 -4060
rect 11300 -4180 11500 -4140
rect 11300 -4260 11360 -4180
rect 11440 -4260 11500 -4180
rect 11300 -4300 11500 -4260
rect 11300 -4380 11360 -4300
rect 11440 -4380 11500 -4300
rect 11300 -4420 11500 -4380
rect 11300 -4500 11360 -4420
rect 11440 -4500 11500 -4420
rect 11300 -4540 11500 -4500
rect 11300 -4620 11360 -4540
rect 11440 -4620 11500 -4540
rect 11300 -4660 11500 -4620
rect 11300 -4740 11360 -4660
rect 11440 -4740 11500 -4660
rect 11300 -4780 11500 -4740
rect 11300 -4860 11360 -4780
rect 11440 -4860 11500 -4780
rect 11300 -4900 11500 -4860
rect 11300 -4980 11360 -4900
rect 11440 -4980 11500 -4900
rect 11300 -5020 11500 -4980
rect 11300 -5100 11360 -5020
rect 11440 -5100 11500 -5020
rect 11300 -5140 11500 -5100
rect 11300 -5220 11360 -5140
rect 11440 -5220 11500 -5140
rect 11660 -5080 11720 -4000
rect 11820 -5080 11880 -4000
rect 11980 -5080 12040 -4000
rect 11660 -5160 12040 -5080
rect 12540 -5080 12600 -4000
rect 12700 -5080 12760 -4000
rect 12860 -5080 12920 -4000
rect 12540 -5160 12920 -5080
rect 13140 -4020 13660 -3980
rect 13700 -3920 17220 -3820
rect 13700 -3980 13740 -3920
rect 15260 -3980 15540 -3920
rect 17060 -3980 17220 -3920
rect 13700 -4000 17220 -3980
rect 13140 -4100 13220 -4020
rect 13300 -4100 13360 -4020
rect 13440 -4100 13500 -4020
rect 13580 -4100 13660 -4020
rect 13140 -4140 13660 -4100
rect 13140 -4220 13220 -4140
rect 13300 -4220 13360 -4140
rect 13440 -4220 13500 -4140
rect 13580 -4220 13660 -4140
rect 13140 -4260 13660 -4220
rect 13140 -4340 13220 -4260
rect 13300 -4340 13360 -4260
rect 13440 -4340 13500 -4260
rect 13580 -4340 13660 -4260
rect 13140 -4380 13660 -4340
rect 13140 -4460 13220 -4380
rect 13300 -4460 13360 -4380
rect 13440 -4460 13500 -4380
rect 13580 -4460 13660 -4380
rect 13140 -4500 13660 -4460
rect 13140 -4580 13220 -4500
rect 13300 -4580 13360 -4500
rect 13440 -4580 13500 -4500
rect 13580 -4580 13660 -4500
rect 13140 -4620 13660 -4580
rect 13140 -4700 13220 -4620
rect 13300 -4700 13360 -4620
rect 13440 -4700 13500 -4620
rect 13580 -4700 13660 -4620
rect 13140 -4740 13660 -4700
rect 13140 -4820 13220 -4740
rect 13300 -4820 13360 -4740
rect 13440 -4820 13500 -4740
rect 13580 -4820 13660 -4740
rect 13140 -4860 13660 -4820
rect 13140 -4940 13220 -4860
rect 13300 -4940 13360 -4860
rect 13440 -4940 13500 -4860
rect 13580 -4940 13660 -4860
rect 13140 -4980 13660 -4940
rect 13140 -5060 13220 -4980
rect 13300 -5060 13360 -4980
rect 13440 -5060 13500 -4980
rect 13580 -5060 13660 -4980
rect 13140 -5100 13660 -5060
rect 11300 -5260 11500 -5220
rect 11300 -5300 11360 -5260
rect 9700 -5340 11360 -5300
rect 11440 -5300 11500 -5260
rect 13140 -5180 13220 -5100
rect 13300 -5180 13360 -5100
rect 13440 -5180 13500 -5100
rect 13580 -5180 13660 -5100
rect 13860 -5080 13920 -4000
rect 14020 -5080 14080 -4000
rect 14180 -5080 14240 -4000
rect 13860 -5160 14240 -5080
rect 14740 -5080 14800 -4000
rect 14900 -5080 14960 -4000
rect 15060 -5080 15120 -4000
rect 14740 -5160 15120 -5080
rect 15300 -4060 15500 -4040
rect 15300 -4140 15360 -4060
rect 15440 -4140 15500 -4060
rect 15300 -4180 15500 -4140
rect 15300 -4260 15360 -4180
rect 15440 -4260 15500 -4180
rect 15300 -4300 15500 -4260
rect 15300 -4380 15360 -4300
rect 15440 -4380 15500 -4300
rect 15300 -4420 15500 -4380
rect 15300 -4500 15360 -4420
rect 15440 -4500 15500 -4420
rect 15300 -4540 15500 -4500
rect 15300 -4620 15360 -4540
rect 15440 -4620 15500 -4540
rect 15300 -4660 15500 -4620
rect 15300 -4740 15360 -4660
rect 15440 -4740 15500 -4660
rect 15300 -4780 15500 -4740
rect 15300 -4860 15360 -4780
rect 15440 -4860 15500 -4780
rect 15300 -4900 15500 -4860
rect 15300 -4980 15360 -4900
rect 15440 -4980 15500 -4900
rect 15300 -5020 15500 -4980
rect 15300 -5100 15360 -5020
rect 15440 -5100 15500 -5020
rect 15300 -5140 15500 -5100
rect 13140 -5220 13660 -5180
rect 13140 -5300 13220 -5220
rect 13300 -5300 13360 -5220
rect 13440 -5300 13500 -5220
rect 13580 -5300 13660 -5220
rect 15300 -5220 15360 -5140
rect 15440 -5220 15500 -5140
rect 15660 -5080 15720 -4000
rect 15820 -5080 15880 -4000
rect 15980 -5080 16040 -4000
rect 15660 -5160 16040 -5080
rect 16540 -5080 16600 -4000
rect 16700 -5080 16760 -4000
rect 16860 -5080 16920 -4000
rect 16540 -5160 16920 -5080
rect 15300 -5260 15500 -5220
rect 15300 -5300 15360 -5260
rect 11440 -5340 15360 -5300
rect 15440 -5300 15500 -5260
rect 15440 -5340 17100 -5300
rect 9700 -5420 9740 -5340
rect 9820 -5420 9860 -5340
rect 9940 -5420 9980 -5340
rect 10060 -5420 10100 -5340
rect 10180 -5420 10220 -5340
rect 10300 -5420 10340 -5340
rect 10420 -5420 10460 -5340
rect 10540 -5420 10580 -5340
rect 10660 -5420 10700 -5340
rect 10780 -5420 10820 -5340
rect 10900 -5420 10940 -5340
rect 11020 -5420 11060 -5340
rect 11140 -5420 11180 -5340
rect 11260 -5380 11540 -5340
rect 11260 -5420 11360 -5380
rect 9700 -5460 11360 -5420
rect 11440 -5420 11540 -5380
rect 11620 -5420 11660 -5340
rect 11740 -5420 11780 -5340
rect 11860 -5420 11900 -5340
rect 11980 -5420 12020 -5340
rect 12100 -5420 12140 -5340
rect 12220 -5420 12260 -5340
rect 12340 -5420 12380 -5340
rect 12460 -5420 12500 -5340
rect 12580 -5420 12620 -5340
rect 12700 -5420 12740 -5340
rect 12820 -5420 12860 -5340
rect 12940 -5420 12980 -5340
rect 13060 -5420 13100 -5340
rect 13180 -5420 13220 -5340
rect 13300 -5420 13360 -5340
rect 13440 -5420 13500 -5340
rect 13580 -5420 13620 -5340
rect 13700 -5420 13740 -5340
rect 13820 -5420 13860 -5340
rect 13940 -5420 13980 -5340
rect 14060 -5420 14100 -5340
rect 14180 -5420 14220 -5340
rect 14300 -5420 14340 -5340
rect 14420 -5420 14460 -5340
rect 14540 -5420 14580 -5340
rect 14660 -5420 14700 -5340
rect 14780 -5420 14820 -5340
rect 14900 -5420 14940 -5340
rect 15020 -5420 15060 -5340
rect 15140 -5420 15180 -5340
rect 15260 -5380 15540 -5340
rect 15260 -5420 15360 -5380
rect 11440 -5460 15360 -5420
rect 15440 -5420 15540 -5380
rect 15620 -5420 15660 -5340
rect 15740 -5420 15780 -5340
rect 15860 -5420 15900 -5340
rect 15980 -5420 16020 -5340
rect 16100 -5420 16140 -5340
rect 16220 -5420 16260 -5340
rect 16340 -5420 16380 -5340
rect 16460 -5420 16500 -5340
rect 16580 -5420 16620 -5340
rect 16700 -5420 16740 -5340
rect 16820 -5420 16860 -5340
rect 16940 -5420 16980 -5340
rect 17060 -5420 17100 -5340
rect 15440 -5460 17100 -5420
rect 9700 -5480 13220 -5460
rect 9700 -5560 9740 -5480
rect 9820 -5560 9860 -5480
rect 9940 -5560 9980 -5480
rect 10060 -5560 10100 -5480
rect 10180 -5560 10220 -5480
rect 10300 -5560 10340 -5480
rect 10420 -5560 10460 -5480
rect 10540 -5560 10580 -5480
rect 10660 -5560 10700 -5480
rect 10780 -5560 10820 -5480
rect 10900 -5560 10940 -5480
rect 11020 -5560 11060 -5480
rect 11140 -5560 11180 -5480
rect 11260 -5500 11540 -5480
rect 11260 -5560 11360 -5500
rect 9700 -5580 11360 -5560
rect 11440 -5560 11540 -5500
rect 11620 -5560 11660 -5480
rect 11740 -5560 11780 -5480
rect 11860 -5560 11900 -5480
rect 11980 -5560 12020 -5480
rect 12100 -5560 12140 -5480
rect 12220 -5560 12260 -5480
rect 12340 -5560 12380 -5480
rect 12460 -5560 12500 -5480
rect 12580 -5560 12620 -5480
rect 12700 -5560 12740 -5480
rect 12820 -5560 12860 -5480
rect 12940 -5560 12980 -5480
rect 13060 -5560 13100 -5480
rect 13180 -5540 13220 -5480
rect 13300 -5540 13360 -5460
rect 13440 -5540 13500 -5460
rect 13580 -5480 17100 -5460
rect 13580 -5540 13620 -5480
rect 13180 -5560 13620 -5540
rect 13700 -5560 13740 -5480
rect 13820 -5560 13860 -5480
rect 13940 -5560 13980 -5480
rect 14060 -5560 14100 -5480
rect 14180 -5560 14220 -5480
rect 14300 -5560 14340 -5480
rect 14420 -5560 14460 -5480
rect 14540 -5560 14580 -5480
rect 14660 -5560 14700 -5480
rect 14780 -5560 14820 -5480
rect 14900 -5560 14940 -5480
rect 15020 -5560 15060 -5480
rect 15140 -5560 15180 -5480
rect 15260 -5500 15540 -5480
rect 15260 -5560 15360 -5500
rect 11440 -5580 15360 -5560
rect 15440 -5560 15540 -5500
rect 15620 -5560 15660 -5480
rect 15740 -5560 15780 -5480
rect 15860 -5560 15900 -5480
rect 15980 -5560 16020 -5480
rect 16100 -5560 16140 -5480
rect 16220 -5560 16260 -5480
rect 16340 -5560 16380 -5480
rect 16460 -5560 16500 -5480
rect 16580 -5560 16620 -5480
rect 16700 -5560 16740 -5480
rect 16820 -5560 16860 -5480
rect 16940 -5560 16980 -5480
rect 17060 -5560 17100 -5480
rect 15440 -5580 17100 -5560
rect 9700 -5600 13220 -5580
rect 11300 -5620 11500 -5600
rect 11300 -5700 11360 -5620
rect 11440 -5700 11500 -5620
rect 11300 -5740 11500 -5700
rect 13140 -5660 13220 -5600
rect 13300 -5660 13360 -5580
rect 13440 -5660 13500 -5580
rect 13580 -5600 17100 -5580
rect 13580 -5660 13660 -5600
rect 13140 -5700 13660 -5660
rect 9860 -5820 10240 -5740
rect 9860 -6900 9920 -5820
rect 10020 -6900 10080 -5820
rect 10180 -6900 10240 -5820
rect 10740 -5820 11120 -5740
rect 10740 -6900 10800 -5820
rect 10900 -6900 10960 -5820
rect 11060 -6900 11120 -5820
rect 11300 -5820 11360 -5740
rect 11440 -5820 11500 -5740
rect 11300 -5860 11500 -5820
rect 11300 -5940 11360 -5860
rect 11440 -5940 11500 -5860
rect 11300 -5980 11500 -5940
rect 11300 -6060 11360 -5980
rect 11440 -6060 11500 -5980
rect 11300 -6100 11500 -6060
rect 11300 -6180 11360 -6100
rect 11440 -6180 11500 -6100
rect 11300 -6220 11500 -6180
rect 11300 -6300 11360 -6220
rect 11440 -6300 11500 -6220
rect 11300 -6340 11500 -6300
rect 11300 -6420 11360 -6340
rect 11440 -6420 11500 -6340
rect 11300 -6460 11500 -6420
rect 11300 -6540 11360 -6460
rect 11440 -6540 11500 -6460
rect 11300 -6580 11500 -6540
rect 11300 -6660 11360 -6580
rect 11440 -6660 11500 -6580
rect 11300 -6700 11500 -6660
rect 11300 -6780 11360 -6700
rect 11440 -6780 11500 -6700
rect 11300 -6860 11500 -6780
rect 11660 -5820 12040 -5740
rect 11660 -6900 11720 -5820
rect 11820 -6900 11880 -5820
rect 11980 -6900 12040 -5820
rect 12540 -5820 12920 -5740
rect 12540 -6900 12600 -5820
rect 12700 -6900 12760 -5820
rect 12860 -6900 12920 -5820
rect 13140 -5780 13220 -5700
rect 13300 -5780 13360 -5700
rect 13440 -5780 13500 -5700
rect 13580 -5780 13660 -5700
rect 15300 -5620 15500 -5600
rect 15300 -5700 15360 -5620
rect 15440 -5700 15500 -5620
rect 15300 -5740 15500 -5700
rect 13140 -5820 13660 -5780
rect 13140 -5900 13220 -5820
rect 13300 -5900 13360 -5820
rect 13440 -5900 13500 -5820
rect 13580 -5900 13660 -5820
rect 13140 -5940 13660 -5900
rect 13140 -6020 13220 -5940
rect 13300 -6020 13360 -5940
rect 13440 -6020 13500 -5940
rect 13580 -6020 13660 -5940
rect 13140 -6060 13660 -6020
rect 13140 -6140 13220 -6060
rect 13300 -6140 13360 -6060
rect 13440 -6140 13500 -6060
rect 13580 -6140 13660 -6060
rect 13140 -6180 13660 -6140
rect 13140 -6260 13220 -6180
rect 13300 -6260 13360 -6180
rect 13440 -6260 13500 -6180
rect 13580 -6260 13660 -6180
rect 13140 -6300 13660 -6260
rect 13140 -6380 13220 -6300
rect 13300 -6380 13360 -6300
rect 13440 -6380 13500 -6300
rect 13580 -6380 13660 -6300
rect 13140 -6420 13660 -6380
rect 13140 -6500 13220 -6420
rect 13300 -6500 13360 -6420
rect 13440 -6500 13500 -6420
rect 13580 -6500 13660 -6420
rect 13140 -6540 13660 -6500
rect 13140 -6620 13220 -6540
rect 13300 -6620 13360 -6540
rect 13440 -6620 13500 -6540
rect 13580 -6620 13660 -6540
rect 13140 -6660 13660 -6620
rect 13140 -6740 13220 -6660
rect 13300 -6740 13360 -6660
rect 13440 -6740 13500 -6660
rect 13580 -6740 13660 -6660
rect 13140 -6780 13660 -6740
rect 13140 -6860 13220 -6780
rect 13300 -6860 13360 -6780
rect 13440 -6860 13500 -6780
rect 13580 -6860 13660 -6780
rect 13140 -6900 13660 -6860
rect 13860 -5820 14240 -5740
rect 13860 -6900 13920 -5820
rect 14020 -6900 14080 -5820
rect 14180 -6900 14240 -5820
rect 14740 -5820 15120 -5740
rect 14740 -6900 14800 -5820
rect 14900 -6900 14960 -5820
rect 15060 -6900 15120 -5820
rect 15300 -5820 15360 -5740
rect 15440 -5820 15500 -5740
rect 15300 -5860 15500 -5820
rect 15300 -5940 15360 -5860
rect 15440 -5940 15500 -5860
rect 15300 -5980 15500 -5940
rect 15300 -6060 15360 -5980
rect 15440 -6060 15500 -5980
rect 15300 -6100 15500 -6060
rect 15300 -6180 15360 -6100
rect 15440 -6180 15500 -6100
rect 15300 -6220 15500 -6180
rect 15300 -6300 15360 -6220
rect 15440 -6300 15500 -6220
rect 15300 -6340 15500 -6300
rect 15300 -6420 15360 -6340
rect 15440 -6420 15500 -6340
rect 15300 -6460 15500 -6420
rect 15300 -6540 15360 -6460
rect 15440 -6540 15500 -6460
rect 15300 -6580 15500 -6540
rect 15300 -6660 15360 -6580
rect 15440 -6660 15500 -6580
rect 15300 -6700 15500 -6660
rect 15300 -6780 15360 -6700
rect 15440 -6780 15500 -6700
rect 15300 -6860 15500 -6780
rect 15660 -5820 16040 -5740
rect 15660 -6900 15720 -5820
rect 15820 -6900 15880 -5820
rect 15980 -6900 16040 -5820
rect 16540 -5820 16920 -5740
rect 16540 -6900 16600 -5820
rect 16700 -6900 16760 -5820
rect 16860 -6900 16920 -5820
rect 17140 -6900 17220 -4000
rect 9580 -6920 13100 -6900
rect 9580 -6980 9740 -6920
rect 11260 -6980 11540 -6920
rect 13060 -6980 13100 -6920
rect 9580 -7080 13100 -6980
rect 13140 -6980 13220 -6900
rect 13300 -6980 13360 -6900
rect 13440 -6980 13500 -6900
rect 13580 -6980 13660 -6900
rect 13140 -7060 13660 -6980
rect 13700 -6920 17220 -6900
rect 13700 -6980 13740 -6920
rect 15260 -6980 15540 -6920
rect 17060 -6980 17220 -6920
rect 9400 -7100 13100 -7080
rect 13700 -7080 17220 -6980
rect 17280 -5340 17500 -3820
rect 17540 -3720 19820 -3560
rect 17540 -3780 17820 -3720
rect 18580 -3780 19820 -3720
rect 17540 -3800 19820 -3780
rect 17540 -3820 17800 -3800
rect 17540 -5080 17720 -3820
rect 17780 -5080 17800 -3820
rect 17540 -5100 17800 -5080
rect 18600 -3820 19820 -3800
rect 18600 -5080 18620 -3820
rect 18680 -5080 19820 -3820
rect 18600 -5100 19820 -5080
rect 17540 -5120 19820 -5100
rect 17540 -5180 17820 -5120
rect 18580 -5180 19820 -5120
rect 17540 -5300 19820 -5180
rect 17280 -5380 19760 -5340
rect 17280 -5460 18020 -5380
rect 18100 -5460 18140 -5380
rect 18280 -5460 18320 -5380
rect 18400 -5460 19760 -5380
rect 17280 -5560 19760 -5460
rect 17280 -5620 17500 -5560
rect 18960 -5620 19760 -5560
rect 17280 -5640 19760 -5620
rect 17280 -5660 17480 -5640
rect 17280 -7080 17400 -5660
rect 13700 -7100 17400 -7080
rect 9400 -7120 17400 -7100
rect 9400 -7180 9620 -7120
rect 17180 -7180 17400 -7120
rect 9400 -7200 17400 -7180
rect 9400 -7220 10300 -7200
rect 9400 -7400 10220 -7220
rect 9320 -7420 10220 -7400
rect 7040 -7440 10220 -7420
rect 7040 -7500 7840 -7440
rect 9300 -7500 10220 -7440
rect 7040 -8980 10220 -7500
rect 10280 -8980 10300 -7220
rect 16400 -7220 17400 -7200
rect 10880 -7280 15870 -7270
rect 7040 -9000 10300 -8980
rect 10440 -7380 10820 -7300
rect 10440 -9000 10500 -7380
rect 10600 -9000 10660 -7380
rect 10760 -9000 10820 -7380
rect 10880 -7330 15880 -7280
rect 10880 -8940 11040 -7330
rect 11200 -7380 11240 -7370
rect 11810 -7380 11850 -7370
rect 11140 -9000 11280 -7380
rect 11760 -9000 11900 -7380
rect 12060 -8940 12220 -7330
rect 12430 -7380 12470 -7370
rect 12380 -9000 12520 -7380
rect 13000 -9000 13140 -7380
rect 13300 -8940 13460 -7330
rect 13600 -9000 13740 -7380
rect 14240 -9000 14380 -7380
rect 14520 -8940 14680 -7330
rect 14840 -9000 14980 -7380
rect 15440 -9000 15580 -7380
rect 15720 -8940 15880 -7330
rect 15940 -7380 16320 -7300
rect 15940 -9000 16000 -7380
rect 16100 -9000 16160 -7380
rect 16260 -9000 16320 -7380
rect 16400 -8980 16420 -7220
rect 16480 -7400 17400 -7220
rect 17460 -7400 17480 -5660
rect 17840 -7240 18000 -5640
rect 18440 -7240 18600 -5640
rect 18980 -5660 19760 -5640
rect 16480 -7420 17480 -7400
rect 18980 -7400 19000 -5660
rect 19060 -7400 19760 -5660
rect 18980 -7420 19760 -7400
rect 16480 -7440 19760 -7420
rect 16480 -7500 17500 -7440
rect 18960 -7500 19760 -7440
rect 16480 -8980 19760 -7500
rect 16400 -9000 19760 -8980
rect 7040 -9020 19760 -9000
rect 7040 -9080 10320 -9020
rect 16380 -9080 19760 -9020
rect 7040 -9160 19760 -9080
rect 6800 -9200 7000 -9180
rect 6800 -9220 10100 -9200
rect 6800 -9380 7020 -9220
rect 9880 -9380 9940 -9220
rect 6800 -9400 9940 -9380
rect 9900 -10380 9940 -9400
rect 10060 -10200 10100 -9220
rect 10140 -9220 16620 -9160
rect 19800 -9180 19820 -5300
rect 19980 -9180 20000 -820
rect 19800 -9200 20000 -9180
rect 10140 -9300 10160 -9220
rect 10240 -9300 10280 -9220
rect 10360 -9300 10400 -9220
rect 10480 -9300 10520 -9220
rect 10600 -9300 10640 -9220
rect 10720 -9300 10760 -9220
rect 10840 -9300 10880 -9220
rect 10960 -9300 11000 -9220
rect 11080 -9300 11120 -9220
rect 11200 -9300 11240 -9220
rect 11320 -9300 11360 -9220
rect 11440 -9300 11480 -9220
rect 11560 -9300 11600 -9220
rect 11680 -9300 11720 -9220
rect 11800 -9300 11840 -9220
rect 11920 -9300 11960 -9220
rect 12040 -9300 12080 -9220
rect 12160 -9300 12200 -9220
rect 12280 -9300 12320 -9220
rect 12400 -9300 12440 -9220
rect 12520 -9300 12560 -9220
rect 12640 -9300 12680 -9220
rect 12760 -9300 12800 -9220
rect 12880 -9300 12920 -9220
rect 13000 -9300 13040 -9220
rect 13120 -9300 13160 -9220
rect 13240 -9300 13280 -9220
rect 13360 -9300 13400 -9220
rect 13480 -9300 13520 -9220
rect 13600 -9300 13640 -9220
rect 13720 -9300 13760 -9220
rect 13840 -9300 13880 -9220
rect 13960 -9300 14000 -9220
rect 14080 -9300 14120 -9220
rect 14200 -9300 14240 -9220
rect 14320 -9300 14360 -9220
rect 14440 -9300 14480 -9220
rect 14560 -9300 14600 -9220
rect 14680 -9300 14720 -9220
rect 14800 -9300 14840 -9220
rect 14920 -9300 14960 -9220
rect 15040 -9300 15080 -9220
rect 15160 -9300 15200 -9220
rect 15280 -9300 15320 -9220
rect 15400 -9300 15440 -9220
rect 15520 -9300 15560 -9220
rect 15640 -9300 15680 -9220
rect 15760 -9300 15800 -9220
rect 15880 -9300 15920 -9220
rect 16000 -9300 16040 -9220
rect 16120 -9300 16160 -9220
rect 16240 -9300 16280 -9220
rect 16360 -9300 16400 -9220
rect 16480 -9300 16520 -9220
rect 16600 -9300 16620 -9220
rect 10140 -9340 16620 -9300
rect 10140 -9420 10160 -9340
rect 10240 -9420 10280 -9340
rect 10360 -9420 10400 -9340
rect 10480 -9420 10520 -9340
rect 10600 -9420 10640 -9340
rect 10720 -9420 10760 -9340
rect 10840 -9420 10880 -9340
rect 10960 -9420 11000 -9340
rect 11080 -9420 11120 -9340
rect 11200 -9420 11240 -9340
rect 11320 -9420 11360 -9340
rect 11440 -9420 11480 -9340
rect 11560 -9420 11600 -9340
rect 11680 -9420 11720 -9340
rect 11800 -9420 11840 -9340
rect 11920 -9420 11960 -9340
rect 12040 -9420 12080 -9340
rect 12160 -9420 12200 -9340
rect 12280 -9420 12320 -9340
rect 12400 -9420 12440 -9340
rect 12520 -9420 12560 -9340
rect 12640 -9420 12680 -9340
rect 12760 -9420 12800 -9340
rect 12880 -9420 12920 -9340
rect 13000 -9420 13040 -9340
rect 13120 -9420 13160 -9340
rect 13240 -9420 13280 -9340
rect 13360 -9420 13400 -9340
rect 13480 -9420 13520 -9340
rect 13600 -9420 13640 -9340
rect 13720 -9420 13760 -9340
rect 13840 -9420 13880 -9340
rect 13960 -9420 14000 -9340
rect 14080 -9420 14120 -9340
rect 14200 -9420 14240 -9340
rect 14320 -9420 14360 -9340
rect 14440 -9420 14480 -9340
rect 14560 -9420 14600 -9340
rect 14680 -9420 14720 -9340
rect 14800 -9420 14840 -9340
rect 14920 -9420 14960 -9340
rect 15040 -9420 15080 -9340
rect 15160 -9420 15200 -9340
rect 15280 -9420 15320 -9340
rect 15400 -9420 15440 -9340
rect 15520 -9420 15560 -9340
rect 15640 -9420 15680 -9340
rect 15760 -9420 15800 -9340
rect 15880 -9420 15920 -9340
rect 16000 -9420 16040 -9340
rect 16120 -9420 16160 -9340
rect 16240 -9420 16280 -9340
rect 16360 -9420 16400 -9340
rect 16480 -9420 16520 -9340
rect 16600 -9420 16620 -9340
rect 10140 -9460 16620 -9420
rect 10140 -9540 10160 -9460
rect 10240 -9540 10280 -9460
rect 10360 -9540 10400 -9460
rect 10480 -9540 10520 -9460
rect 10600 -9540 10640 -9460
rect 10720 -9540 10760 -9460
rect 10840 -9540 10880 -9460
rect 10960 -9540 11000 -9460
rect 11080 -9540 11120 -9460
rect 11200 -9540 11240 -9460
rect 11320 -9540 11360 -9460
rect 11440 -9540 11480 -9460
rect 11560 -9540 11600 -9460
rect 11680 -9540 11720 -9460
rect 11800 -9540 11840 -9460
rect 11920 -9540 11960 -9460
rect 12040 -9540 12080 -9460
rect 12160 -9540 12200 -9460
rect 12280 -9540 12320 -9460
rect 12400 -9540 12440 -9460
rect 12520 -9540 12560 -9460
rect 12640 -9540 12680 -9460
rect 12760 -9540 12800 -9460
rect 12880 -9540 12920 -9460
rect 13000 -9540 13040 -9460
rect 13120 -9540 13160 -9460
rect 13240 -9540 13280 -9460
rect 13360 -9540 13400 -9460
rect 13480 -9540 13520 -9460
rect 13600 -9540 13640 -9460
rect 13720 -9540 13760 -9460
rect 13840 -9540 13880 -9460
rect 13960 -9540 14000 -9460
rect 14080 -9540 14120 -9460
rect 14200 -9540 14240 -9460
rect 14320 -9540 14360 -9460
rect 14440 -9540 14480 -9460
rect 14560 -9540 14600 -9460
rect 14680 -9540 14720 -9460
rect 14800 -9540 14840 -9460
rect 14920 -9540 14960 -9460
rect 15040 -9540 15080 -9460
rect 15160 -9540 15200 -9460
rect 15280 -9540 15320 -9460
rect 15400 -9540 15440 -9460
rect 15520 -9540 15560 -9460
rect 15640 -9540 15680 -9460
rect 15760 -9540 15800 -9460
rect 15880 -9540 15920 -9460
rect 16000 -9540 16040 -9460
rect 16120 -9540 16160 -9460
rect 16240 -9540 16280 -9460
rect 16360 -9540 16400 -9460
rect 16480 -9540 16520 -9460
rect 16600 -9540 16620 -9460
rect 10140 -9580 16620 -9540
rect 10140 -9660 10160 -9580
rect 10240 -9660 10280 -9580
rect 10360 -9660 10400 -9580
rect 10480 -9660 10520 -9580
rect 10600 -9660 10640 -9580
rect 10720 -9660 10760 -9580
rect 10840 -9660 10880 -9580
rect 10960 -9660 11000 -9580
rect 11080 -9660 11120 -9580
rect 11200 -9660 11240 -9580
rect 11320 -9660 11360 -9580
rect 11440 -9660 11480 -9580
rect 11560 -9660 11600 -9580
rect 11680 -9660 11720 -9580
rect 11800 -9660 11840 -9580
rect 11920 -9660 11960 -9580
rect 12040 -9660 12080 -9580
rect 12160 -9660 12200 -9580
rect 12280 -9660 12320 -9580
rect 12400 -9660 12440 -9580
rect 12520 -9660 12560 -9580
rect 12640 -9660 12680 -9580
rect 12760 -9660 12800 -9580
rect 12880 -9660 12920 -9580
rect 13000 -9660 13040 -9580
rect 13120 -9660 13160 -9580
rect 13240 -9660 13280 -9580
rect 13360 -9660 13400 -9580
rect 13480 -9660 13520 -9580
rect 13600 -9660 13640 -9580
rect 13720 -9660 13760 -9580
rect 13840 -9660 13880 -9580
rect 13960 -9660 14000 -9580
rect 14080 -9660 14120 -9580
rect 14200 -9660 14240 -9580
rect 14320 -9660 14360 -9580
rect 14440 -9660 14480 -9580
rect 14560 -9660 14600 -9580
rect 14680 -9660 14720 -9580
rect 14800 -9660 14840 -9580
rect 14920 -9660 14960 -9580
rect 15040 -9660 15080 -9580
rect 15160 -9660 15200 -9580
rect 15280 -9660 15320 -9580
rect 15400 -9660 15440 -9580
rect 15520 -9660 15560 -9580
rect 15640 -9660 15680 -9580
rect 15760 -9660 15800 -9580
rect 15880 -9660 15920 -9580
rect 16000 -9660 16040 -9580
rect 16120 -9660 16160 -9580
rect 16240 -9660 16280 -9580
rect 16360 -9660 16400 -9580
rect 16480 -9660 16520 -9580
rect 16600 -9660 16620 -9580
rect 10140 -9700 16620 -9660
rect 10140 -9780 10160 -9700
rect 10240 -9780 10280 -9700
rect 10360 -9780 10400 -9700
rect 10480 -9780 10520 -9700
rect 10600 -9780 10640 -9700
rect 10720 -9780 10760 -9700
rect 10840 -9780 10880 -9700
rect 10960 -9780 11000 -9700
rect 11080 -9780 11120 -9700
rect 11200 -9780 11240 -9700
rect 11320 -9780 11360 -9700
rect 11440 -9780 11480 -9700
rect 11560 -9780 11600 -9700
rect 11680 -9780 11720 -9700
rect 11800 -9780 11840 -9700
rect 11920 -9780 11960 -9700
rect 12040 -9780 12080 -9700
rect 12160 -9780 12200 -9700
rect 12280 -9780 12320 -9700
rect 12400 -9780 12440 -9700
rect 12520 -9780 12560 -9700
rect 12640 -9780 12680 -9700
rect 12760 -9780 12800 -9700
rect 12880 -9780 12920 -9700
rect 13000 -9780 13040 -9700
rect 13120 -9780 13160 -9700
rect 13240 -9780 13280 -9700
rect 13360 -9780 13400 -9700
rect 13480 -9780 13520 -9700
rect 13600 -9780 13640 -9700
rect 13720 -9780 13760 -9700
rect 13840 -9780 13880 -9700
rect 13960 -9780 14000 -9700
rect 14080 -9780 14120 -9700
rect 14200 -9780 14240 -9700
rect 14320 -9780 14360 -9700
rect 14440 -9780 14480 -9700
rect 14560 -9780 14600 -9700
rect 14680 -9780 14720 -9700
rect 14800 -9780 14840 -9700
rect 14920 -9780 14960 -9700
rect 15040 -9780 15080 -9700
rect 15160 -9780 15200 -9700
rect 15280 -9780 15320 -9700
rect 15400 -9780 15440 -9700
rect 15520 -9780 15560 -9700
rect 15640 -9780 15680 -9700
rect 15760 -9780 15800 -9700
rect 15880 -9780 15920 -9700
rect 16000 -9780 16040 -9700
rect 16120 -9780 16160 -9700
rect 16240 -9780 16280 -9700
rect 16360 -9780 16400 -9700
rect 16480 -9780 16520 -9700
rect 16600 -9780 16620 -9700
rect 10140 -9820 16620 -9780
rect 10140 -9900 10160 -9820
rect 10240 -9900 10280 -9820
rect 10360 -9900 10400 -9820
rect 10480 -9900 10520 -9820
rect 10600 -9900 10640 -9820
rect 10720 -9900 10760 -9820
rect 10840 -9900 10880 -9820
rect 10960 -9900 11000 -9820
rect 11080 -9900 11120 -9820
rect 11200 -9900 11240 -9820
rect 11320 -9900 11360 -9820
rect 11440 -9900 11480 -9820
rect 11560 -9900 11600 -9820
rect 11680 -9900 11720 -9820
rect 11800 -9900 11840 -9820
rect 11920 -9900 11960 -9820
rect 12040 -9900 12080 -9820
rect 12160 -9900 12200 -9820
rect 12280 -9900 12320 -9820
rect 12400 -9900 12440 -9820
rect 12520 -9900 12560 -9820
rect 12640 -9900 12680 -9820
rect 12760 -9900 12800 -9820
rect 12880 -9900 12920 -9820
rect 13000 -9900 13040 -9820
rect 13120 -9900 13160 -9820
rect 13240 -9900 13280 -9820
rect 13360 -9900 13400 -9820
rect 13480 -9900 13520 -9820
rect 13600 -9900 13640 -9820
rect 13720 -9900 13760 -9820
rect 13840 -9900 13880 -9820
rect 13960 -9900 14000 -9820
rect 14080 -9900 14120 -9820
rect 14200 -9900 14240 -9820
rect 14320 -9900 14360 -9820
rect 14440 -9900 14480 -9820
rect 14560 -9900 14600 -9820
rect 14680 -9900 14720 -9820
rect 14800 -9900 14840 -9820
rect 14920 -9900 14960 -9820
rect 15040 -9900 15080 -9820
rect 15160 -9900 15200 -9820
rect 15280 -9900 15320 -9820
rect 15400 -9900 15440 -9820
rect 15520 -9900 15560 -9820
rect 15640 -9900 15680 -9820
rect 15760 -9900 15800 -9820
rect 15880 -9900 15920 -9820
rect 16000 -9900 16040 -9820
rect 16120 -9900 16160 -9820
rect 16240 -9900 16280 -9820
rect 16360 -9900 16400 -9820
rect 16480 -9900 16520 -9820
rect 16600 -9900 16620 -9820
rect 10140 -9940 16620 -9900
rect 10140 -10020 10160 -9940
rect 10240 -10020 10280 -9940
rect 10360 -10020 10400 -9940
rect 10480 -10020 10520 -9940
rect 10600 -10020 10640 -9940
rect 10720 -10020 10760 -9940
rect 10840 -10020 10880 -9940
rect 10960 -10020 11000 -9940
rect 11080 -10020 11120 -9940
rect 11200 -10020 11240 -9940
rect 11320 -10020 11360 -9940
rect 11440 -10020 11480 -9940
rect 11560 -10020 11600 -9940
rect 11680 -10020 11720 -9940
rect 11800 -10020 11840 -9940
rect 11920 -10020 11960 -9940
rect 12040 -10020 12080 -9940
rect 12160 -10020 12200 -9940
rect 12280 -10020 12320 -9940
rect 12400 -10020 12440 -9940
rect 12520 -10020 12560 -9940
rect 12640 -10020 12680 -9940
rect 12760 -10020 12800 -9940
rect 12880 -10020 12920 -9940
rect 13000 -10020 13040 -9940
rect 13120 -10020 13160 -9940
rect 13240 -10020 13280 -9940
rect 13360 -10020 13400 -9940
rect 13480 -10020 13520 -9940
rect 13600 -10020 13640 -9940
rect 13720 -10020 13760 -9940
rect 13840 -10020 13880 -9940
rect 13960 -10020 14000 -9940
rect 14080 -10020 14120 -9940
rect 14200 -10020 14240 -9940
rect 14320 -10020 14360 -9940
rect 14440 -10020 14480 -9940
rect 14560 -10020 14600 -9940
rect 14680 -10020 14720 -9940
rect 14800 -10020 14840 -9940
rect 14920 -10020 14960 -9940
rect 15040 -10020 15080 -9940
rect 15160 -10020 15200 -9940
rect 15280 -10020 15320 -9940
rect 15400 -10020 15440 -9940
rect 15520 -10020 15560 -9940
rect 15640 -10020 15680 -9940
rect 15760 -10020 15800 -9940
rect 15880 -10020 15920 -9940
rect 16000 -10020 16040 -9940
rect 16120 -10020 16160 -9940
rect 16240 -10020 16280 -9940
rect 16360 -10020 16400 -9940
rect 16480 -10020 16520 -9940
rect 16600 -10020 16620 -9940
rect 10140 -10060 16620 -10020
rect 10140 -10140 10160 -10060
rect 10240 -10140 10280 -10060
rect 10360 -10140 10400 -10060
rect 10480 -10140 10520 -10060
rect 10600 -10140 10640 -10060
rect 10720 -10140 10760 -10060
rect 10840 -10140 10880 -10060
rect 10960 -10140 11000 -10060
rect 11080 -10140 11120 -10060
rect 11200 -10140 11240 -10060
rect 11320 -10140 11360 -10060
rect 11440 -10140 11480 -10060
rect 11560 -10140 11600 -10060
rect 11680 -10140 11720 -10060
rect 11800 -10140 11840 -10060
rect 11920 -10140 11960 -10060
rect 12040 -10140 12080 -10060
rect 12160 -10140 12200 -10060
rect 12280 -10140 12320 -10060
rect 12400 -10140 12440 -10060
rect 12520 -10140 12560 -10060
rect 12640 -10140 12680 -10060
rect 12760 -10140 12800 -10060
rect 12880 -10140 12920 -10060
rect 13000 -10140 13040 -10060
rect 13120 -10140 13160 -10060
rect 13240 -10140 13280 -10060
rect 13360 -10140 13400 -10060
rect 13480 -10140 13520 -10060
rect 13600 -10140 13640 -10060
rect 13720 -10140 13760 -10060
rect 13840 -10140 13880 -10060
rect 13960 -10140 14000 -10060
rect 14080 -10140 14120 -10060
rect 14200 -10140 14240 -10060
rect 14320 -10140 14360 -10060
rect 14440 -10140 14480 -10060
rect 14560 -10140 14600 -10060
rect 14680 -10140 14720 -10060
rect 14800 -10140 14840 -10060
rect 14920 -10140 14960 -10060
rect 15040 -10140 15080 -10060
rect 15160 -10140 15200 -10060
rect 15280 -10140 15320 -10060
rect 15400 -10140 15440 -10060
rect 15520 -10140 15560 -10060
rect 15640 -10140 15680 -10060
rect 15760 -10140 15800 -10060
rect 15880 -10140 15920 -10060
rect 16000 -10140 16040 -10060
rect 16120 -10140 16160 -10060
rect 16240 -10140 16280 -10060
rect 16360 -10140 16400 -10060
rect 16480 -10140 16520 -10060
rect 16600 -10140 16620 -10060
rect 10140 -10160 16620 -10140
rect 16660 -9220 20000 -9200
rect 16660 -10200 16700 -9220
rect 10060 -10220 16700 -10200
rect 10060 -10380 10100 -10220
rect 16660 -10380 16700 -10220
rect 16820 -9380 16860 -9220
rect 19780 -9380 20000 -9220
rect 16820 -9400 20000 -9380
rect 16820 -10380 16860 -9400
rect 9900 -10400 16860 -10380
<< viali >>
rect 10160 20 10240 100
rect 10280 20 10360 100
rect 10400 20 10480 100
rect 10520 20 10600 100
rect 10640 20 10720 100
rect 10760 20 10840 100
rect 10880 20 10960 100
rect 11000 20 11080 100
rect 11120 20 11200 100
rect 11240 20 11320 100
rect 11360 20 11440 100
rect 11480 20 11560 100
rect 11600 20 11680 100
rect 11720 20 11800 100
rect 11840 20 11920 100
rect 11960 20 12040 100
rect 12080 20 12160 100
rect 12200 20 12280 100
rect 12320 20 12400 100
rect 12440 20 12520 100
rect 12560 20 12640 100
rect 12680 20 12760 100
rect 12800 20 12880 100
rect 12920 20 13000 100
rect 13040 20 13120 100
rect 13160 20 13240 100
rect 13280 20 13360 100
rect 13400 20 13480 100
rect 13520 20 13600 100
rect 13640 20 13720 100
rect 13760 20 13840 100
rect 13880 20 13960 100
rect 14000 20 14080 100
rect 14120 20 14200 100
rect 14240 20 14320 100
rect 14360 20 14440 100
rect 14480 20 14560 100
rect 14600 20 14680 100
rect 14720 20 14800 100
rect 14840 20 14920 100
rect 14960 20 15040 100
rect 15080 20 15160 100
rect 15200 20 15280 100
rect 15320 20 15400 100
rect 15440 20 15520 100
rect 15560 20 15640 100
rect 15680 20 15760 100
rect 15800 20 15880 100
rect 15920 20 16000 100
rect 16040 20 16120 100
rect 16160 20 16240 100
rect 16280 20 16360 100
rect 16400 20 16480 100
rect 16520 20 16600 100
rect 10160 -100 10240 -20
rect 10280 -100 10360 -20
rect 10400 -100 10480 -20
rect 10520 -100 10600 -20
rect 10640 -100 10720 -20
rect 10760 -100 10840 -20
rect 10880 -100 10960 -20
rect 11000 -100 11080 -20
rect 11120 -100 11200 -20
rect 11240 -100 11320 -20
rect 11360 -100 11440 -20
rect 11480 -100 11560 -20
rect 11600 -100 11680 -20
rect 11720 -100 11800 -20
rect 11840 -100 11920 -20
rect 11960 -100 12040 -20
rect 12080 -100 12160 -20
rect 12200 -100 12280 -20
rect 12320 -100 12400 -20
rect 12440 -100 12520 -20
rect 12560 -100 12640 -20
rect 12680 -100 12760 -20
rect 12800 -100 12880 -20
rect 12920 -100 13000 -20
rect 13040 -100 13120 -20
rect 13160 -100 13240 -20
rect 13280 -100 13360 -20
rect 13400 -100 13480 -20
rect 13520 -100 13600 -20
rect 13640 -100 13720 -20
rect 13760 -100 13840 -20
rect 13880 -100 13960 -20
rect 14000 -100 14080 -20
rect 14120 -100 14200 -20
rect 14240 -100 14320 -20
rect 14360 -100 14440 -20
rect 14480 -100 14560 -20
rect 14600 -100 14680 -20
rect 14720 -100 14800 -20
rect 14840 -100 14920 -20
rect 14960 -100 15040 -20
rect 15080 -100 15160 -20
rect 15200 -100 15280 -20
rect 15320 -100 15400 -20
rect 15440 -100 15520 -20
rect 15560 -100 15640 -20
rect 15680 -100 15760 -20
rect 15800 -100 15880 -20
rect 15920 -100 16000 -20
rect 16040 -100 16120 -20
rect 16160 -100 16240 -20
rect 16280 -100 16360 -20
rect 16400 -100 16480 -20
rect 16520 -100 16600 -20
rect 10160 -220 10240 -140
rect 10280 -220 10360 -140
rect 10400 -220 10480 -140
rect 10520 -220 10600 -140
rect 10640 -220 10720 -140
rect 10760 -220 10840 -140
rect 10880 -220 10960 -140
rect 11000 -220 11080 -140
rect 11120 -220 11200 -140
rect 11240 -220 11320 -140
rect 11360 -220 11440 -140
rect 11480 -220 11560 -140
rect 11600 -220 11680 -140
rect 11720 -220 11800 -140
rect 11840 -220 11920 -140
rect 11960 -220 12040 -140
rect 12080 -220 12160 -140
rect 12200 -220 12280 -140
rect 12320 -220 12400 -140
rect 12440 -220 12520 -140
rect 12560 -220 12640 -140
rect 12680 -220 12760 -140
rect 12800 -220 12880 -140
rect 12920 -220 13000 -140
rect 13040 -220 13120 -140
rect 13160 -220 13240 -140
rect 13280 -220 13360 -140
rect 13400 -220 13480 -140
rect 13520 -220 13600 -140
rect 13640 -220 13720 -140
rect 13760 -220 13840 -140
rect 13880 -220 13960 -140
rect 14000 -220 14080 -140
rect 14120 -220 14200 -140
rect 14240 -220 14320 -140
rect 14360 -220 14440 -140
rect 14480 -220 14560 -140
rect 14600 -220 14680 -140
rect 14720 -220 14800 -140
rect 14840 -220 14920 -140
rect 14960 -220 15040 -140
rect 15080 -220 15160 -140
rect 15200 -220 15280 -140
rect 15320 -220 15400 -140
rect 15440 -220 15520 -140
rect 15560 -220 15640 -140
rect 15680 -220 15760 -140
rect 15800 -220 15880 -140
rect 15920 -220 16000 -140
rect 16040 -220 16120 -140
rect 16160 -220 16240 -140
rect 16280 -220 16360 -140
rect 16400 -220 16480 -140
rect 16520 -220 16600 -140
rect 10160 -340 10240 -260
rect 10280 -340 10360 -260
rect 10400 -340 10480 -260
rect 10520 -340 10600 -260
rect 10640 -340 10720 -260
rect 10760 -340 10840 -260
rect 10880 -340 10960 -260
rect 11000 -340 11080 -260
rect 11120 -340 11200 -260
rect 11240 -340 11320 -260
rect 11360 -340 11440 -260
rect 11480 -340 11560 -260
rect 11600 -340 11680 -260
rect 11720 -340 11800 -260
rect 11840 -340 11920 -260
rect 11960 -340 12040 -260
rect 12080 -340 12160 -260
rect 12200 -340 12280 -260
rect 12320 -340 12400 -260
rect 12440 -340 12520 -260
rect 12560 -340 12640 -260
rect 12680 -340 12760 -260
rect 12800 -340 12880 -260
rect 12920 -340 13000 -260
rect 13040 -340 13120 -260
rect 13160 -340 13240 -260
rect 13280 -340 13360 -260
rect 13400 -340 13480 -260
rect 13520 -340 13600 -260
rect 13640 -340 13720 -260
rect 13760 -340 13840 -260
rect 13880 -340 13960 -260
rect 14000 -340 14080 -260
rect 14120 -340 14200 -260
rect 14240 -340 14320 -260
rect 14360 -340 14440 -260
rect 14480 -340 14560 -260
rect 14600 -340 14680 -260
rect 14720 -340 14800 -260
rect 14840 -340 14920 -260
rect 14960 -340 15040 -260
rect 15080 -340 15160 -260
rect 15200 -340 15280 -260
rect 15320 -340 15400 -260
rect 15440 -340 15520 -260
rect 15560 -340 15640 -260
rect 15680 -340 15760 -260
rect 15800 -340 15880 -260
rect 15920 -340 16000 -260
rect 16040 -340 16120 -260
rect 16160 -340 16240 -260
rect 16280 -340 16360 -260
rect 16400 -340 16480 -260
rect 16520 -340 16600 -260
rect 10160 -460 10240 -380
rect 10280 -460 10360 -380
rect 10400 -460 10480 -380
rect 10520 -460 10600 -380
rect 10640 -460 10720 -380
rect 10760 -460 10840 -380
rect 10880 -460 10960 -380
rect 11000 -460 11080 -380
rect 11120 -460 11200 -380
rect 11240 -460 11320 -380
rect 11360 -460 11440 -380
rect 11480 -460 11560 -380
rect 11600 -460 11680 -380
rect 11720 -460 11800 -380
rect 11840 -460 11920 -380
rect 11960 -460 12040 -380
rect 12080 -460 12160 -380
rect 12200 -460 12280 -380
rect 12320 -460 12400 -380
rect 12440 -460 12520 -380
rect 12560 -460 12640 -380
rect 12680 -460 12760 -380
rect 12800 -460 12880 -380
rect 12920 -460 13000 -380
rect 13040 -460 13120 -380
rect 13160 -460 13240 -380
rect 13280 -460 13360 -380
rect 13400 -460 13480 -380
rect 13520 -460 13600 -380
rect 13640 -460 13720 -380
rect 13760 -460 13840 -380
rect 13880 -460 13960 -380
rect 14000 -460 14080 -380
rect 14120 -460 14200 -380
rect 14240 -460 14320 -380
rect 14360 -460 14440 -380
rect 14480 -460 14560 -380
rect 14600 -460 14680 -380
rect 14720 -460 14800 -380
rect 14840 -460 14920 -380
rect 14960 -460 15040 -380
rect 15080 -460 15160 -380
rect 15200 -460 15280 -380
rect 15320 -460 15400 -380
rect 15440 -460 15520 -380
rect 15560 -460 15640 -380
rect 15680 -460 15760 -380
rect 15800 -460 15880 -380
rect 15920 -460 16000 -380
rect 16040 -460 16120 -380
rect 16160 -460 16240 -380
rect 16280 -460 16360 -380
rect 16400 -460 16480 -380
rect 16520 -460 16600 -380
rect 10160 -580 10240 -500
rect 10280 -580 10360 -500
rect 10400 -580 10480 -500
rect 10520 -580 10600 -500
rect 10640 -580 10720 -500
rect 10760 -580 10840 -500
rect 10880 -580 10960 -500
rect 11000 -580 11080 -500
rect 11120 -580 11200 -500
rect 11240 -580 11320 -500
rect 11360 -580 11440 -500
rect 11480 -580 11560 -500
rect 11600 -580 11680 -500
rect 11720 -580 11800 -500
rect 11840 -580 11920 -500
rect 11960 -580 12040 -500
rect 12080 -580 12160 -500
rect 12200 -580 12280 -500
rect 12320 -580 12400 -500
rect 12440 -580 12520 -500
rect 12560 -580 12640 -500
rect 12680 -580 12760 -500
rect 12800 -580 12880 -500
rect 12920 -580 13000 -500
rect 13040 -580 13120 -500
rect 13160 -580 13240 -500
rect 13280 -580 13360 -500
rect 13400 -580 13480 -500
rect 13520 -580 13600 -500
rect 13640 -580 13720 -500
rect 13760 -580 13840 -500
rect 13880 -580 13960 -500
rect 14000 -580 14080 -500
rect 14120 -580 14200 -500
rect 14240 -580 14320 -500
rect 14360 -580 14440 -500
rect 14480 -580 14560 -500
rect 14600 -580 14680 -500
rect 14720 -580 14800 -500
rect 14840 -580 14920 -500
rect 14960 -580 15040 -500
rect 15080 -580 15160 -500
rect 15200 -580 15280 -500
rect 15320 -580 15400 -500
rect 15440 -580 15520 -500
rect 15560 -580 15640 -500
rect 15680 -580 15760 -500
rect 15800 -580 15880 -500
rect 15920 -580 16000 -500
rect 16040 -580 16120 -500
rect 16160 -580 16240 -500
rect 16280 -580 16360 -500
rect 16400 -580 16480 -500
rect 16520 -580 16600 -500
rect 8440 -5460 8520 -5380
rect 8580 -5460 8680 -5380
rect 8740 -5460 8820 -5380
rect 13220 -3980 13300 -3900
rect 13360 -3980 13440 -3900
rect 13500 -3980 13580 -3900
rect 11360 -4140 11440 -4060
rect 11360 -4260 11440 -4180
rect 11360 -4380 11440 -4300
rect 11360 -4500 11440 -4420
rect 11360 -4620 11440 -4540
rect 11360 -4740 11440 -4660
rect 11360 -4860 11440 -4780
rect 11360 -4980 11440 -4900
rect 11360 -5100 11440 -5020
rect 11360 -5220 11440 -5140
rect 13220 -4100 13300 -4020
rect 13360 -4100 13440 -4020
rect 13500 -4100 13580 -4020
rect 13220 -4220 13300 -4140
rect 13360 -4220 13440 -4140
rect 13500 -4220 13580 -4140
rect 13220 -4340 13300 -4260
rect 13360 -4340 13440 -4260
rect 13500 -4340 13580 -4260
rect 13220 -4460 13300 -4380
rect 13360 -4460 13440 -4380
rect 13500 -4460 13580 -4380
rect 13220 -4580 13300 -4500
rect 13360 -4580 13440 -4500
rect 13500 -4580 13580 -4500
rect 13220 -4700 13300 -4620
rect 13360 -4700 13440 -4620
rect 13500 -4700 13580 -4620
rect 13220 -4820 13300 -4740
rect 13360 -4820 13440 -4740
rect 13500 -4820 13580 -4740
rect 13220 -4940 13300 -4860
rect 13360 -4940 13440 -4860
rect 13500 -4940 13580 -4860
rect 13220 -5060 13300 -4980
rect 13360 -5060 13440 -4980
rect 13500 -5060 13580 -4980
rect 11360 -5340 11440 -5260
rect 13220 -5180 13300 -5100
rect 13360 -5180 13440 -5100
rect 13500 -5180 13580 -5100
rect 15360 -4140 15440 -4060
rect 15360 -4260 15440 -4180
rect 15360 -4380 15440 -4300
rect 15360 -4500 15440 -4420
rect 15360 -4620 15440 -4540
rect 15360 -4740 15440 -4660
rect 15360 -4860 15440 -4780
rect 15360 -4980 15440 -4900
rect 15360 -5100 15440 -5020
rect 13220 -5300 13300 -5220
rect 13360 -5300 13440 -5220
rect 13500 -5300 13580 -5220
rect 15360 -5220 15440 -5140
rect 15360 -5340 15440 -5260
rect 9740 -5420 9820 -5340
rect 9860 -5420 9940 -5340
rect 9980 -5420 10060 -5340
rect 10100 -5420 10180 -5340
rect 10220 -5420 10300 -5340
rect 10340 -5420 10420 -5340
rect 10460 -5420 10540 -5340
rect 10580 -5420 10660 -5340
rect 10700 -5420 10780 -5340
rect 10820 -5420 10900 -5340
rect 10940 -5420 11020 -5340
rect 11060 -5420 11140 -5340
rect 11180 -5420 11260 -5340
rect 11360 -5460 11440 -5380
rect 11540 -5420 11620 -5340
rect 11660 -5420 11740 -5340
rect 11780 -5420 11860 -5340
rect 11900 -5420 11980 -5340
rect 12020 -5420 12100 -5340
rect 12140 -5420 12220 -5340
rect 12260 -5420 12340 -5340
rect 12380 -5420 12460 -5340
rect 12500 -5420 12580 -5340
rect 12620 -5420 12700 -5340
rect 12740 -5420 12820 -5340
rect 12860 -5420 12940 -5340
rect 12980 -5420 13060 -5340
rect 13100 -5420 13180 -5340
rect 13220 -5420 13300 -5340
rect 13360 -5420 13440 -5340
rect 13500 -5420 13580 -5340
rect 13620 -5420 13700 -5340
rect 13740 -5420 13820 -5340
rect 13860 -5420 13940 -5340
rect 13980 -5420 14060 -5340
rect 14100 -5420 14180 -5340
rect 14220 -5420 14300 -5340
rect 14340 -5420 14420 -5340
rect 14460 -5420 14540 -5340
rect 14580 -5420 14660 -5340
rect 14700 -5420 14780 -5340
rect 14820 -5420 14900 -5340
rect 14940 -5420 15020 -5340
rect 15060 -5420 15140 -5340
rect 15180 -5420 15260 -5340
rect 15360 -5460 15440 -5380
rect 15540 -5420 15620 -5340
rect 15660 -5420 15740 -5340
rect 15780 -5420 15860 -5340
rect 15900 -5420 15980 -5340
rect 16020 -5420 16100 -5340
rect 16140 -5420 16220 -5340
rect 16260 -5420 16340 -5340
rect 16380 -5420 16460 -5340
rect 16500 -5420 16580 -5340
rect 16620 -5420 16700 -5340
rect 16740 -5420 16820 -5340
rect 16860 -5420 16940 -5340
rect 16980 -5420 17060 -5340
rect 9740 -5560 9820 -5480
rect 9860 -5560 9940 -5480
rect 9980 -5560 10060 -5480
rect 10100 -5560 10180 -5480
rect 10220 -5560 10300 -5480
rect 10340 -5560 10420 -5480
rect 10460 -5560 10540 -5480
rect 10580 -5560 10660 -5480
rect 10700 -5560 10780 -5480
rect 10820 -5560 10900 -5480
rect 10940 -5560 11020 -5480
rect 11060 -5560 11140 -5480
rect 11180 -5560 11260 -5480
rect 11360 -5580 11440 -5500
rect 11540 -5560 11620 -5480
rect 11660 -5560 11740 -5480
rect 11780 -5560 11860 -5480
rect 11900 -5560 11980 -5480
rect 12020 -5560 12100 -5480
rect 12140 -5560 12220 -5480
rect 12260 -5560 12340 -5480
rect 12380 -5560 12460 -5480
rect 12500 -5560 12580 -5480
rect 12620 -5560 12700 -5480
rect 12740 -5560 12820 -5480
rect 12860 -5560 12940 -5480
rect 12980 -5560 13060 -5480
rect 13100 -5560 13180 -5480
rect 13220 -5540 13300 -5460
rect 13360 -5540 13440 -5460
rect 13500 -5540 13580 -5460
rect 13620 -5560 13700 -5480
rect 13740 -5560 13820 -5480
rect 13860 -5560 13940 -5480
rect 13980 -5560 14060 -5480
rect 14100 -5560 14180 -5480
rect 14220 -5560 14300 -5480
rect 14340 -5560 14420 -5480
rect 14460 -5560 14540 -5480
rect 14580 -5560 14660 -5480
rect 14700 -5560 14780 -5480
rect 14820 -5560 14900 -5480
rect 14940 -5560 15020 -5480
rect 15060 -5560 15140 -5480
rect 15180 -5560 15260 -5480
rect 15360 -5580 15440 -5500
rect 15540 -5560 15620 -5480
rect 15660 -5560 15740 -5480
rect 15780 -5560 15860 -5480
rect 15900 -5560 15980 -5480
rect 16020 -5560 16100 -5480
rect 16140 -5560 16220 -5480
rect 16260 -5560 16340 -5480
rect 16380 -5560 16460 -5480
rect 16500 -5560 16580 -5480
rect 16620 -5560 16700 -5480
rect 16740 -5560 16820 -5480
rect 16860 -5560 16940 -5480
rect 16980 -5560 17060 -5480
rect 11360 -5700 11440 -5620
rect 13220 -5660 13300 -5580
rect 13360 -5660 13440 -5580
rect 13500 -5660 13580 -5580
rect 11360 -5820 11440 -5740
rect 11360 -5940 11440 -5860
rect 11360 -6060 11440 -5980
rect 11360 -6180 11440 -6100
rect 11360 -6300 11440 -6220
rect 11360 -6420 11440 -6340
rect 11360 -6540 11440 -6460
rect 11360 -6660 11440 -6580
rect 11360 -6780 11440 -6700
rect 13220 -5780 13300 -5700
rect 13360 -5780 13440 -5700
rect 13500 -5780 13580 -5700
rect 15360 -5700 15440 -5620
rect 13220 -5900 13300 -5820
rect 13360 -5900 13440 -5820
rect 13500 -5900 13580 -5820
rect 13220 -6020 13300 -5940
rect 13360 -6020 13440 -5940
rect 13500 -6020 13580 -5940
rect 13220 -6140 13300 -6060
rect 13360 -6140 13440 -6060
rect 13500 -6140 13580 -6060
rect 13220 -6260 13300 -6180
rect 13360 -6260 13440 -6180
rect 13500 -6260 13580 -6180
rect 13220 -6380 13300 -6300
rect 13360 -6380 13440 -6300
rect 13500 -6380 13580 -6300
rect 13220 -6500 13300 -6420
rect 13360 -6500 13440 -6420
rect 13500 -6500 13580 -6420
rect 13220 -6620 13300 -6540
rect 13360 -6620 13440 -6540
rect 13500 -6620 13580 -6540
rect 13220 -6740 13300 -6660
rect 13360 -6740 13440 -6660
rect 13500 -6740 13580 -6660
rect 13220 -6860 13300 -6780
rect 13360 -6860 13440 -6780
rect 13500 -6860 13580 -6780
rect 15360 -5820 15440 -5740
rect 15360 -5940 15440 -5860
rect 15360 -6060 15440 -5980
rect 15360 -6180 15440 -6100
rect 15360 -6300 15440 -6220
rect 15360 -6420 15440 -6340
rect 15360 -6540 15440 -6460
rect 15360 -6660 15440 -6580
rect 15360 -6780 15440 -6700
rect 13220 -6980 13300 -6900
rect 13360 -6980 13440 -6900
rect 13500 -6980 13580 -6900
rect 18020 -5460 18100 -5380
rect 18140 -5460 18280 -5380
rect 18320 -5460 18400 -5380
rect 10160 -9300 10240 -9220
rect 10280 -9300 10360 -9220
rect 10400 -9300 10480 -9220
rect 10520 -9300 10600 -9220
rect 10640 -9300 10720 -9220
rect 10760 -9300 10840 -9220
rect 10880 -9300 10960 -9220
rect 11000 -9300 11080 -9220
rect 11120 -9300 11200 -9220
rect 11240 -9300 11320 -9220
rect 11360 -9300 11440 -9220
rect 11480 -9300 11560 -9220
rect 11600 -9300 11680 -9220
rect 11720 -9300 11800 -9220
rect 11840 -9300 11920 -9220
rect 11960 -9300 12040 -9220
rect 12080 -9300 12160 -9220
rect 12200 -9300 12280 -9220
rect 12320 -9300 12400 -9220
rect 12440 -9300 12520 -9220
rect 12560 -9300 12640 -9220
rect 12680 -9300 12760 -9220
rect 12800 -9300 12880 -9220
rect 12920 -9300 13000 -9220
rect 13040 -9300 13120 -9220
rect 13160 -9300 13240 -9220
rect 13280 -9300 13360 -9220
rect 13400 -9300 13480 -9220
rect 13520 -9300 13600 -9220
rect 13640 -9300 13720 -9220
rect 13760 -9300 13840 -9220
rect 13880 -9300 13960 -9220
rect 14000 -9300 14080 -9220
rect 14120 -9300 14200 -9220
rect 14240 -9300 14320 -9220
rect 14360 -9300 14440 -9220
rect 14480 -9300 14560 -9220
rect 14600 -9300 14680 -9220
rect 14720 -9300 14800 -9220
rect 14840 -9300 14920 -9220
rect 14960 -9300 15040 -9220
rect 15080 -9300 15160 -9220
rect 15200 -9300 15280 -9220
rect 15320 -9300 15400 -9220
rect 15440 -9300 15520 -9220
rect 15560 -9300 15640 -9220
rect 15680 -9300 15760 -9220
rect 15800 -9300 15880 -9220
rect 15920 -9300 16000 -9220
rect 16040 -9300 16120 -9220
rect 16160 -9300 16240 -9220
rect 16280 -9300 16360 -9220
rect 16400 -9300 16480 -9220
rect 16520 -9300 16600 -9220
rect 10160 -9420 10240 -9340
rect 10280 -9420 10360 -9340
rect 10400 -9420 10480 -9340
rect 10520 -9420 10600 -9340
rect 10640 -9420 10720 -9340
rect 10760 -9420 10840 -9340
rect 10880 -9420 10960 -9340
rect 11000 -9420 11080 -9340
rect 11120 -9420 11200 -9340
rect 11240 -9420 11320 -9340
rect 11360 -9420 11440 -9340
rect 11480 -9420 11560 -9340
rect 11600 -9420 11680 -9340
rect 11720 -9420 11800 -9340
rect 11840 -9420 11920 -9340
rect 11960 -9420 12040 -9340
rect 12080 -9420 12160 -9340
rect 12200 -9420 12280 -9340
rect 12320 -9420 12400 -9340
rect 12440 -9420 12520 -9340
rect 12560 -9420 12640 -9340
rect 12680 -9420 12760 -9340
rect 12800 -9420 12880 -9340
rect 12920 -9420 13000 -9340
rect 13040 -9420 13120 -9340
rect 13160 -9420 13240 -9340
rect 13280 -9420 13360 -9340
rect 13400 -9420 13480 -9340
rect 13520 -9420 13600 -9340
rect 13640 -9420 13720 -9340
rect 13760 -9420 13840 -9340
rect 13880 -9420 13960 -9340
rect 14000 -9420 14080 -9340
rect 14120 -9420 14200 -9340
rect 14240 -9420 14320 -9340
rect 14360 -9420 14440 -9340
rect 14480 -9420 14560 -9340
rect 14600 -9420 14680 -9340
rect 14720 -9420 14800 -9340
rect 14840 -9420 14920 -9340
rect 14960 -9420 15040 -9340
rect 15080 -9420 15160 -9340
rect 15200 -9420 15280 -9340
rect 15320 -9420 15400 -9340
rect 15440 -9420 15520 -9340
rect 15560 -9420 15640 -9340
rect 15680 -9420 15760 -9340
rect 15800 -9420 15880 -9340
rect 15920 -9420 16000 -9340
rect 16040 -9420 16120 -9340
rect 16160 -9420 16240 -9340
rect 16280 -9420 16360 -9340
rect 16400 -9420 16480 -9340
rect 16520 -9420 16600 -9340
rect 10160 -9540 10240 -9460
rect 10280 -9540 10360 -9460
rect 10400 -9540 10480 -9460
rect 10520 -9540 10600 -9460
rect 10640 -9540 10720 -9460
rect 10760 -9540 10840 -9460
rect 10880 -9540 10960 -9460
rect 11000 -9540 11080 -9460
rect 11120 -9540 11200 -9460
rect 11240 -9540 11320 -9460
rect 11360 -9540 11440 -9460
rect 11480 -9540 11560 -9460
rect 11600 -9540 11680 -9460
rect 11720 -9540 11800 -9460
rect 11840 -9540 11920 -9460
rect 11960 -9540 12040 -9460
rect 12080 -9540 12160 -9460
rect 12200 -9540 12280 -9460
rect 12320 -9540 12400 -9460
rect 12440 -9540 12520 -9460
rect 12560 -9540 12640 -9460
rect 12680 -9540 12760 -9460
rect 12800 -9540 12880 -9460
rect 12920 -9540 13000 -9460
rect 13040 -9540 13120 -9460
rect 13160 -9540 13240 -9460
rect 13280 -9540 13360 -9460
rect 13400 -9540 13480 -9460
rect 13520 -9540 13600 -9460
rect 13640 -9540 13720 -9460
rect 13760 -9540 13840 -9460
rect 13880 -9540 13960 -9460
rect 14000 -9540 14080 -9460
rect 14120 -9540 14200 -9460
rect 14240 -9540 14320 -9460
rect 14360 -9540 14440 -9460
rect 14480 -9540 14560 -9460
rect 14600 -9540 14680 -9460
rect 14720 -9540 14800 -9460
rect 14840 -9540 14920 -9460
rect 14960 -9540 15040 -9460
rect 15080 -9540 15160 -9460
rect 15200 -9540 15280 -9460
rect 15320 -9540 15400 -9460
rect 15440 -9540 15520 -9460
rect 15560 -9540 15640 -9460
rect 15680 -9540 15760 -9460
rect 15800 -9540 15880 -9460
rect 15920 -9540 16000 -9460
rect 16040 -9540 16120 -9460
rect 16160 -9540 16240 -9460
rect 16280 -9540 16360 -9460
rect 16400 -9540 16480 -9460
rect 16520 -9540 16600 -9460
rect 10160 -9660 10240 -9580
rect 10280 -9660 10360 -9580
rect 10400 -9660 10480 -9580
rect 10520 -9660 10600 -9580
rect 10640 -9660 10720 -9580
rect 10760 -9660 10840 -9580
rect 10880 -9660 10960 -9580
rect 11000 -9660 11080 -9580
rect 11120 -9660 11200 -9580
rect 11240 -9660 11320 -9580
rect 11360 -9660 11440 -9580
rect 11480 -9660 11560 -9580
rect 11600 -9660 11680 -9580
rect 11720 -9660 11800 -9580
rect 11840 -9660 11920 -9580
rect 11960 -9660 12040 -9580
rect 12080 -9660 12160 -9580
rect 12200 -9660 12280 -9580
rect 12320 -9660 12400 -9580
rect 12440 -9660 12520 -9580
rect 12560 -9660 12640 -9580
rect 12680 -9660 12760 -9580
rect 12800 -9660 12880 -9580
rect 12920 -9660 13000 -9580
rect 13040 -9660 13120 -9580
rect 13160 -9660 13240 -9580
rect 13280 -9660 13360 -9580
rect 13400 -9660 13480 -9580
rect 13520 -9660 13600 -9580
rect 13640 -9660 13720 -9580
rect 13760 -9660 13840 -9580
rect 13880 -9660 13960 -9580
rect 14000 -9660 14080 -9580
rect 14120 -9660 14200 -9580
rect 14240 -9660 14320 -9580
rect 14360 -9660 14440 -9580
rect 14480 -9660 14560 -9580
rect 14600 -9660 14680 -9580
rect 14720 -9660 14800 -9580
rect 14840 -9660 14920 -9580
rect 14960 -9660 15040 -9580
rect 15080 -9660 15160 -9580
rect 15200 -9660 15280 -9580
rect 15320 -9660 15400 -9580
rect 15440 -9660 15520 -9580
rect 15560 -9660 15640 -9580
rect 15680 -9660 15760 -9580
rect 15800 -9660 15880 -9580
rect 15920 -9660 16000 -9580
rect 16040 -9660 16120 -9580
rect 16160 -9660 16240 -9580
rect 16280 -9660 16360 -9580
rect 16400 -9660 16480 -9580
rect 16520 -9660 16600 -9580
rect 10160 -9780 10240 -9700
rect 10280 -9780 10360 -9700
rect 10400 -9780 10480 -9700
rect 10520 -9780 10600 -9700
rect 10640 -9780 10720 -9700
rect 10760 -9780 10840 -9700
rect 10880 -9780 10960 -9700
rect 11000 -9780 11080 -9700
rect 11120 -9780 11200 -9700
rect 11240 -9780 11320 -9700
rect 11360 -9780 11440 -9700
rect 11480 -9780 11560 -9700
rect 11600 -9780 11680 -9700
rect 11720 -9780 11800 -9700
rect 11840 -9780 11920 -9700
rect 11960 -9780 12040 -9700
rect 12080 -9780 12160 -9700
rect 12200 -9780 12280 -9700
rect 12320 -9780 12400 -9700
rect 12440 -9780 12520 -9700
rect 12560 -9780 12640 -9700
rect 12680 -9780 12760 -9700
rect 12800 -9780 12880 -9700
rect 12920 -9780 13000 -9700
rect 13040 -9780 13120 -9700
rect 13160 -9780 13240 -9700
rect 13280 -9780 13360 -9700
rect 13400 -9780 13480 -9700
rect 13520 -9780 13600 -9700
rect 13640 -9780 13720 -9700
rect 13760 -9780 13840 -9700
rect 13880 -9780 13960 -9700
rect 14000 -9780 14080 -9700
rect 14120 -9780 14200 -9700
rect 14240 -9780 14320 -9700
rect 14360 -9780 14440 -9700
rect 14480 -9780 14560 -9700
rect 14600 -9780 14680 -9700
rect 14720 -9780 14800 -9700
rect 14840 -9780 14920 -9700
rect 14960 -9780 15040 -9700
rect 15080 -9780 15160 -9700
rect 15200 -9780 15280 -9700
rect 15320 -9780 15400 -9700
rect 15440 -9780 15520 -9700
rect 15560 -9780 15640 -9700
rect 15680 -9780 15760 -9700
rect 15800 -9780 15880 -9700
rect 15920 -9780 16000 -9700
rect 16040 -9780 16120 -9700
rect 16160 -9780 16240 -9700
rect 16280 -9780 16360 -9700
rect 16400 -9780 16480 -9700
rect 16520 -9780 16600 -9700
rect 10160 -9900 10240 -9820
rect 10280 -9900 10360 -9820
rect 10400 -9900 10480 -9820
rect 10520 -9900 10600 -9820
rect 10640 -9900 10720 -9820
rect 10760 -9900 10840 -9820
rect 10880 -9900 10960 -9820
rect 11000 -9900 11080 -9820
rect 11120 -9900 11200 -9820
rect 11240 -9900 11320 -9820
rect 11360 -9900 11440 -9820
rect 11480 -9900 11560 -9820
rect 11600 -9900 11680 -9820
rect 11720 -9900 11800 -9820
rect 11840 -9900 11920 -9820
rect 11960 -9900 12040 -9820
rect 12080 -9900 12160 -9820
rect 12200 -9900 12280 -9820
rect 12320 -9900 12400 -9820
rect 12440 -9900 12520 -9820
rect 12560 -9900 12640 -9820
rect 12680 -9900 12760 -9820
rect 12800 -9900 12880 -9820
rect 12920 -9900 13000 -9820
rect 13040 -9900 13120 -9820
rect 13160 -9900 13240 -9820
rect 13280 -9900 13360 -9820
rect 13400 -9900 13480 -9820
rect 13520 -9900 13600 -9820
rect 13640 -9900 13720 -9820
rect 13760 -9900 13840 -9820
rect 13880 -9900 13960 -9820
rect 14000 -9900 14080 -9820
rect 14120 -9900 14200 -9820
rect 14240 -9900 14320 -9820
rect 14360 -9900 14440 -9820
rect 14480 -9900 14560 -9820
rect 14600 -9900 14680 -9820
rect 14720 -9900 14800 -9820
rect 14840 -9900 14920 -9820
rect 14960 -9900 15040 -9820
rect 15080 -9900 15160 -9820
rect 15200 -9900 15280 -9820
rect 15320 -9900 15400 -9820
rect 15440 -9900 15520 -9820
rect 15560 -9900 15640 -9820
rect 15680 -9900 15760 -9820
rect 15800 -9900 15880 -9820
rect 15920 -9900 16000 -9820
rect 16040 -9900 16120 -9820
rect 16160 -9900 16240 -9820
rect 16280 -9900 16360 -9820
rect 16400 -9900 16480 -9820
rect 16520 -9900 16600 -9820
rect 10160 -10020 10240 -9940
rect 10280 -10020 10360 -9940
rect 10400 -10020 10480 -9940
rect 10520 -10020 10600 -9940
rect 10640 -10020 10720 -9940
rect 10760 -10020 10840 -9940
rect 10880 -10020 10960 -9940
rect 11000 -10020 11080 -9940
rect 11120 -10020 11200 -9940
rect 11240 -10020 11320 -9940
rect 11360 -10020 11440 -9940
rect 11480 -10020 11560 -9940
rect 11600 -10020 11680 -9940
rect 11720 -10020 11800 -9940
rect 11840 -10020 11920 -9940
rect 11960 -10020 12040 -9940
rect 12080 -10020 12160 -9940
rect 12200 -10020 12280 -9940
rect 12320 -10020 12400 -9940
rect 12440 -10020 12520 -9940
rect 12560 -10020 12640 -9940
rect 12680 -10020 12760 -9940
rect 12800 -10020 12880 -9940
rect 12920 -10020 13000 -9940
rect 13040 -10020 13120 -9940
rect 13160 -10020 13240 -9940
rect 13280 -10020 13360 -9940
rect 13400 -10020 13480 -9940
rect 13520 -10020 13600 -9940
rect 13640 -10020 13720 -9940
rect 13760 -10020 13840 -9940
rect 13880 -10020 13960 -9940
rect 14000 -10020 14080 -9940
rect 14120 -10020 14200 -9940
rect 14240 -10020 14320 -9940
rect 14360 -10020 14440 -9940
rect 14480 -10020 14560 -9940
rect 14600 -10020 14680 -9940
rect 14720 -10020 14800 -9940
rect 14840 -10020 14920 -9940
rect 14960 -10020 15040 -9940
rect 15080 -10020 15160 -9940
rect 15200 -10020 15280 -9940
rect 15320 -10020 15400 -9940
rect 15440 -10020 15520 -9940
rect 15560 -10020 15640 -9940
rect 15680 -10020 15760 -9940
rect 15800 -10020 15880 -9940
rect 15920 -10020 16000 -9940
rect 16040 -10020 16120 -9940
rect 16160 -10020 16240 -9940
rect 16280 -10020 16360 -9940
rect 16400 -10020 16480 -9940
rect 16520 -10020 16600 -9940
rect 10160 -10140 10240 -10060
rect 10280 -10140 10360 -10060
rect 10400 -10140 10480 -10060
rect 10520 -10140 10600 -10060
rect 10640 -10140 10720 -10060
rect 10760 -10140 10840 -10060
rect 10880 -10140 10960 -10060
rect 11000 -10140 11080 -10060
rect 11120 -10140 11200 -10060
rect 11240 -10140 11320 -10060
rect 11360 -10140 11440 -10060
rect 11480 -10140 11560 -10060
rect 11600 -10140 11680 -10060
rect 11720 -10140 11800 -10060
rect 11840 -10140 11920 -10060
rect 11960 -10140 12040 -10060
rect 12080 -10140 12160 -10060
rect 12200 -10140 12280 -10060
rect 12320 -10140 12400 -10060
rect 12440 -10140 12520 -10060
rect 12560 -10140 12640 -10060
rect 12680 -10140 12760 -10060
rect 12800 -10140 12880 -10060
rect 12920 -10140 13000 -10060
rect 13040 -10140 13120 -10060
rect 13160 -10140 13240 -10060
rect 13280 -10140 13360 -10060
rect 13400 -10140 13480 -10060
rect 13520 -10140 13600 -10060
rect 13640 -10140 13720 -10060
rect 13760 -10140 13840 -10060
rect 13880 -10140 13960 -10060
rect 14000 -10140 14080 -10060
rect 14120 -10140 14200 -10060
rect 14240 -10140 14320 -10060
rect 14360 -10140 14440 -10060
rect 14480 -10140 14560 -10060
rect 14600 -10140 14680 -10060
rect 14720 -10140 14800 -10060
rect 14840 -10140 14920 -10060
rect 14960 -10140 15040 -10060
rect 15080 -10140 15160 -10060
rect 15200 -10140 15280 -10060
rect 15320 -10140 15400 -10060
rect 15440 -10140 15520 -10060
rect 15560 -10140 15640 -10060
rect 15680 -10140 15760 -10060
rect 15800 -10140 15880 -10060
rect 15920 -10140 16000 -10060
rect 16040 -10140 16120 -10060
rect 16160 -10140 16240 -10060
rect 16280 -10140 16360 -10060
rect 16400 -10140 16480 -10060
rect 16520 -10140 16600 -10060
<< metal1 >>
rect 10140 100 16660 120
rect 10140 20 10160 100
rect 10240 20 10280 100
rect 10360 20 10400 100
rect 10480 20 10520 100
rect 10600 20 10640 100
rect 10720 20 10760 100
rect 10840 20 10880 100
rect 10960 20 11000 100
rect 11080 20 11120 100
rect 11200 20 11240 100
rect 11320 20 11360 100
rect 11440 20 11480 100
rect 11560 20 11600 100
rect 11680 20 11720 100
rect 11800 20 11840 100
rect 11920 20 11960 100
rect 12040 20 12080 100
rect 12160 20 12200 100
rect 12280 20 12320 100
rect 12400 20 12440 100
rect 12520 20 12560 100
rect 12640 20 12680 100
rect 12760 20 12800 100
rect 12880 20 12920 100
rect 13000 20 13040 100
rect 13120 20 13160 100
rect 13240 20 13280 100
rect 13360 20 13400 100
rect 13480 20 13520 100
rect 13600 20 13640 100
rect 13720 20 13760 100
rect 13840 20 13880 100
rect 13960 20 14000 100
rect 14080 20 14120 100
rect 14200 20 14240 100
rect 14320 20 14360 100
rect 14440 20 14480 100
rect 14560 20 14600 100
rect 14680 20 14720 100
rect 14800 20 14840 100
rect 14920 20 14960 100
rect 15040 20 15080 100
rect 15160 20 15200 100
rect 15280 20 15320 100
rect 15400 20 15440 100
rect 15520 20 15560 100
rect 15640 20 15680 100
rect 15760 20 15800 100
rect 15880 20 15920 100
rect 16000 20 16040 100
rect 16120 20 16160 100
rect 16240 20 16280 100
rect 16360 20 16400 100
rect 16480 20 16520 100
rect 16600 20 16660 100
rect 10140 -20 16660 20
rect 10140 -100 10160 -20
rect 10240 -100 10280 -20
rect 10360 -100 10400 -20
rect 10480 -100 10520 -20
rect 10600 -100 10640 -20
rect 10720 -100 10760 -20
rect 10840 -100 10880 -20
rect 10960 -100 11000 -20
rect 11080 -100 11120 -20
rect 11200 -100 11240 -20
rect 11320 -100 11360 -20
rect 11440 -100 11480 -20
rect 11560 -100 11600 -20
rect 11680 -100 11720 -20
rect 11800 -100 11840 -20
rect 11920 -100 11960 -20
rect 12040 -100 12080 -20
rect 12160 -100 12200 -20
rect 12280 -100 12320 -20
rect 12400 -100 12440 -20
rect 12520 -100 12560 -20
rect 12640 -100 12680 -20
rect 12760 -100 12800 -20
rect 12880 -100 12920 -20
rect 13000 -100 13040 -20
rect 13120 -100 13160 -20
rect 13240 -100 13280 -20
rect 13360 -100 13400 -20
rect 13480 -100 13520 -20
rect 13600 -100 13640 -20
rect 13720 -100 13760 -20
rect 13840 -100 13880 -20
rect 13960 -100 14000 -20
rect 14080 -100 14120 -20
rect 14200 -100 14240 -20
rect 14320 -100 14360 -20
rect 14440 -100 14480 -20
rect 14560 -100 14600 -20
rect 14680 -100 14720 -20
rect 14800 -100 14840 -20
rect 14920 -100 14960 -20
rect 15040 -100 15080 -20
rect 15160 -100 15200 -20
rect 15280 -100 15320 -20
rect 15400 -100 15440 -20
rect 15520 -100 15560 -20
rect 15640 -100 15680 -20
rect 15760 -100 15800 -20
rect 15880 -100 15920 -20
rect 16000 -100 16040 -20
rect 16120 -100 16160 -20
rect 16240 -100 16280 -20
rect 16360 -100 16400 -20
rect 16480 -100 16520 -20
rect 16600 -100 16660 -20
rect 10140 -140 16660 -100
rect 10140 -220 10160 -140
rect 10240 -220 10280 -140
rect 10360 -220 10400 -140
rect 10480 -220 10520 -140
rect 10600 -220 10640 -140
rect 10720 -220 10760 -140
rect 10840 -220 10880 -140
rect 10960 -220 11000 -140
rect 11080 -220 11120 -140
rect 11200 -220 11240 -140
rect 11320 -220 11360 -140
rect 11440 -220 11480 -140
rect 11560 -220 11600 -140
rect 11680 -220 11720 -140
rect 11800 -220 11840 -140
rect 11920 -220 11960 -140
rect 12040 -220 12080 -140
rect 12160 -220 12200 -140
rect 12280 -220 12320 -140
rect 12400 -220 12440 -140
rect 12520 -220 12560 -140
rect 12640 -220 12680 -140
rect 12760 -220 12800 -140
rect 12880 -220 12920 -140
rect 13000 -220 13040 -140
rect 13120 -220 13160 -140
rect 13240 -220 13280 -140
rect 13360 -220 13400 -140
rect 13480 -220 13520 -140
rect 13600 -220 13640 -140
rect 13720 -220 13760 -140
rect 13840 -220 13880 -140
rect 13960 -220 14000 -140
rect 14080 -220 14120 -140
rect 14200 -220 14240 -140
rect 14320 -220 14360 -140
rect 14440 -220 14480 -140
rect 14560 -220 14600 -140
rect 14680 -220 14720 -140
rect 14800 -220 14840 -140
rect 14920 -220 14960 -140
rect 15040 -220 15080 -140
rect 15160 -220 15200 -140
rect 15280 -220 15320 -140
rect 15400 -220 15440 -140
rect 15520 -220 15560 -140
rect 15640 -220 15680 -140
rect 15760 -220 15800 -140
rect 15880 -220 15920 -140
rect 16000 -220 16040 -140
rect 16120 -220 16160 -140
rect 16240 -220 16280 -140
rect 16360 -220 16400 -140
rect 16480 -220 16520 -140
rect 16600 -220 16660 -140
rect 10140 -260 16660 -220
rect 10140 -340 10160 -260
rect 10240 -340 10280 -260
rect 10360 -340 10400 -260
rect 10480 -340 10520 -260
rect 10600 -340 10640 -260
rect 10720 -340 10760 -260
rect 10840 -340 10880 -260
rect 10960 -340 11000 -260
rect 11080 -340 11120 -260
rect 11200 -340 11240 -260
rect 11320 -340 11360 -260
rect 11440 -340 11480 -260
rect 11560 -340 11600 -260
rect 11680 -340 11720 -260
rect 11800 -340 11840 -260
rect 11920 -340 11960 -260
rect 12040 -340 12080 -260
rect 12160 -340 12200 -260
rect 12280 -340 12320 -260
rect 12400 -340 12440 -260
rect 12520 -340 12560 -260
rect 12640 -340 12680 -260
rect 12760 -340 12800 -260
rect 12880 -340 12920 -260
rect 13000 -340 13040 -260
rect 13120 -340 13160 -260
rect 13240 -340 13280 -260
rect 13360 -340 13400 -260
rect 13480 -340 13520 -260
rect 13600 -340 13640 -260
rect 13720 -340 13760 -260
rect 13840 -340 13880 -260
rect 13960 -340 14000 -260
rect 14080 -340 14120 -260
rect 14200 -340 14240 -260
rect 14320 -340 14360 -260
rect 14440 -340 14480 -260
rect 14560 -340 14600 -260
rect 14680 -340 14720 -260
rect 14800 -340 14840 -260
rect 14920 -340 14960 -260
rect 15040 -340 15080 -260
rect 15160 -340 15200 -260
rect 15280 -340 15320 -260
rect 15400 -340 15440 -260
rect 15520 -340 15560 -260
rect 15640 -340 15680 -260
rect 15760 -340 15800 -260
rect 15880 -340 15920 -260
rect 16000 -340 16040 -260
rect 16120 -340 16160 -260
rect 16240 -340 16280 -260
rect 16360 -340 16400 -260
rect 16480 -340 16520 -260
rect 16600 -340 16660 -260
rect 10140 -380 16660 -340
rect 10140 -460 10160 -380
rect 10240 -460 10280 -380
rect 10360 -460 10400 -380
rect 10480 -460 10520 -380
rect 10600 -460 10640 -380
rect 10720 -460 10760 -380
rect 10840 -460 10880 -380
rect 10960 -460 11000 -380
rect 11080 -460 11120 -380
rect 11200 -460 11240 -380
rect 11320 -460 11360 -380
rect 11440 -460 11480 -380
rect 11560 -460 11600 -380
rect 11680 -460 11720 -380
rect 11800 -460 11840 -380
rect 11920 -460 11960 -380
rect 12040 -460 12080 -380
rect 12160 -460 12200 -380
rect 12280 -460 12320 -380
rect 12400 -460 12440 -380
rect 12520 -460 12560 -380
rect 12640 -460 12680 -380
rect 12760 -460 12800 -380
rect 12880 -460 12920 -380
rect 13000 -460 13040 -380
rect 13120 -460 13160 -380
rect 13240 -460 13280 -380
rect 13360 -460 13400 -380
rect 13480 -460 13520 -380
rect 13600 -460 13640 -380
rect 13720 -460 13760 -380
rect 13840 -460 13880 -380
rect 13960 -460 14000 -380
rect 14080 -460 14120 -380
rect 14200 -460 14240 -380
rect 14320 -460 14360 -380
rect 14440 -460 14480 -380
rect 14560 -460 14600 -380
rect 14680 -460 14720 -380
rect 14800 -460 14840 -380
rect 14920 -460 14960 -380
rect 15040 -460 15080 -380
rect 15160 -460 15200 -380
rect 15280 -460 15320 -380
rect 15400 -460 15440 -380
rect 15520 -460 15560 -380
rect 15640 -460 15680 -380
rect 15760 -460 15800 -380
rect 15880 -460 15920 -380
rect 16000 -460 16040 -380
rect 16120 -460 16160 -380
rect 16240 -460 16280 -380
rect 16360 -460 16400 -380
rect 16480 -460 16520 -380
rect 16600 -460 16660 -380
rect 10140 -500 16660 -460
rect 10140 -580 10160 -500
rect 10240 -580 10280 -500
rect 10360 -580 10400 -500
rect 10480 -580 10520 -500
rect 10600 -580 10640 -500
rect 10720 -580 10760 -500
rect 10840 -580 10880 -500
rect 10960 -580 11000 -500
rect 11080 -580 11120 -500
rect 11200 -580 11240 -500
rect 11320 -580 11360 -500
rect 11440 -580 11480 -500
rect 11560 -580 11600 -500
rect 11680 -580 11720 -500
rect 11800 -580 11840 -500
rect 11920 -580 11960 -500
rect 12040 -580 12080 -500
rect 12160 -580 12200 -500
rect 12280 -580 12320 -500
rect 12400 -580 12440 -500
rect 12520 -580 12560 -500
rect 12640 -580 12680 -500
rect 12760 -580 12800 -500
rect 12880 -580 12920 -500
rect 13000 -580 13040 -500
rect 13120 -580 13160 -500
rect 13240 -580 13280 -500
rect 13360 -580 13400 -500
rect 13480 -580 13520 -500
rect 13600 -580 13640 -500
rect 13720 -580 13760 -500
rect 13840 -580 13880 -500
rect 13960 -580 14000 -500
rect 14080 -580 14120 -500
rect 14200 -580 14240 -500
rect 14320 -580 14360 -500
rect 14440 -580 14480 -500
rect 14560 -580 14600 -500
rect 14680 -580 14720 -500
rect 14800 -580 14840 -500
rect 14920 -580 14960 -500
rect 15040 -580 15080 -500
rect 15160 -580 15200 -500
rect 15280 -580 15320 -500
rect 15400 -580 15440 -500
rect 15520 -580 15560 -500
rect 15640 -580 15680 -500
rect 15760 -580 15800 -500
rect 15880 -580 15920 -500
rect 16000 -580 16040 -500
rect 16120 -580 16160 -500
rect 16240 -580 16280 -500
rect 16360 -580 16400 -500
rect 16480 -580 16520 -500
rect 16600 -580 16660 -500
rect 10140 -600 16660 -580
rect 11380 -1980 11580 -1960
rect 11380 -2040 11400 -1980
rect 11460 -2040 11500 -1980
rect 11560 -2040 11580 -1980
rect 11380 -2060 11580 -2040
rect 11380 -2120 11400 -2060
rect 11460 -2120 11500 -2060
rect 11560 -2120 11580 -2060
rect 11380 -2180 11580 -2120
rect 11380 -2240 11400 -2180
rect 11460 -2240 11500 -2180
rect 11560 -2240 11580 -2180
rect 11380 -2260 11580 -2240
rect 11380 -2320 11400 -2260
rect 11460 -2320 11500 -2260
rect 11560 -2320 11580 -2260
rect 11380 -2340 11580 -2320
rect 12620 -1980 12820 -1960
rect 12620 -2040 12640 -1980
rect 12700 -2040 12740 -1980
rect 12800 -2040 12820 -1980
rect 12620 -2060 12820 -2040
rect 12620 -2120 12640 -2060
rect 12700 -2120 12740 -2060
rect 12800 -2120 12820 -2060
rect 12620 -2180 12820 -2120
rect 12620 -2240 12640 -2180
rect 12700 -2240 12740 -2180
rect 12800 -2240 12820 -2180
rect 12620 -2260 12820 -2240
rect 12620 -2320 12640 -2260
rect 12700 -2320 12740 -2260
rect 12800 -2320 12820 -2260
rect 12620 -2340 12820 -2320
rect 13840 -1980 14040 -1960
rect 13840 -2040 13860 -1980
rect 13920 -2040 13960 -1980
rect 14020 -2040 14040 -1980
rect 13840 -2060 14040 -2040
rect 13840 -2120 13860 -2060
rect 13920 -2120 13960 -2060
rect 14020 -2120 14040 -2060
rect 13840 -2180 14040 -2120
rect 13840 -2240 13860 -2180
rect 13920 -2240 13960 -2180
rect 14020 -2240 14040 -2180
rect 13840 -2260 14040 -2240
rect 13840 -2320 13860 -2260
rect 13920 -2320 13960 -2260
rect 14020 -2320 14040 -2260
rect 13840 -2340 14040 -2320
rect 15080 -1980 15280 -1960
rect 15080 -2040 15100 -1980
rect 15160 -2040 15200 -1980
rect 15260 -2040 15280 -1980
rect 15080 -2060 15280 -2040
rect 15080 -2120 15100 -2060
rect 15160 -2120 15200 -2060
rect 15260 -2120 15280 -2060
rect 15080 -2180 15280 -2120
rect 15080 -2240 15100 -2180
rect 15160 -2240 15200 -2180
rect 15260 -2240 15280 -2180
rect 15080 -2260 15280 -2240
rect 15080 -2320 15100 -2260
rect 15160 -2320 15200 -2260
rect 15260 -2320 15280 -2260
rect 15080 -2340 15280 -2320
rect 10860 -2820 15860 -2620
rect 7380 -2880 7500 -2860
rect 7380 -2940 7400 -2880
rect 7460 -2940 7500 -2880
rect 7380 -3060 7500 -2940
rect 7380 -3120 7400 -3060
rect 7460 -3120 7500 -3060
rect 7380 -3140 7500 -3120
rect 7980 -2880 8100 -2860
rect 7980 -2940 8000 -2880
rect 8060 -2940 8100 -2880
rect 7980 -3060 8100 -2940
rect 7980 -3120 8000 -3060
rect 8060 -3120 8100 -3060
rect 7980 -3140 8100 -3120
rect 8600 -2880 8720 -2860
rect 8600 -2940 8640 -2880
rect 8700 -2940 8720 -2880
rect 8600 -3060 8720 -2940
rect 8600 -3120 8640 -3060
rect 8700 -3120 8720 -3060
rect 8600 -3140 8720 -3120
rect 9220 -2880 9340 -2860
rect 9220 -2940 9240 -2880
rect 9300 -2940 9340 -2880
rect 9220 -3060 9340 -2940
rect 9220 -3120 9240 -3060
rect 9300 -3120 9340 -3060
rect 9220 -3140 9340 -3120
rect 9840 -2880 9960 -2860
rect 9840 -2940 9880 -2880
rect 9940 -2940 9960 -2880
rect 9840 -3060 9960 -2940
rect 9840 -3120 9880 -3060
rect 9940 -3120 9960 -3060
rect 9840 -3140 9960 -3120
rect 11120 -2940 15680 -2820
rect 11120 -3020 11140 -2940
rect 11220 -3020 11260 -2940
rect 11340 -3020 11380 -2940
rect 11460 -3020 11500 -2940
rect 11580 -3020 11620 -2940
rect 11700 -3020 11740 -2940
rect 11820 -3020 11860 -2940
rect 11940 -3020 11980 -2940
rect 12060 -3020 12100 -2940
rect 12180 -3020 12220 -2940
rect 12300 -3020 12340 -2940
rect 12420 -3020 12460 -2940
rect 12540 -3020 12580 -2940
rect 12660 -3020 12700 -2940
rect 12780 -3020 12820 -2940
rect 12900 -3020 12940 -2940
rect 13020 -3020 13060 -2940
rect 13140 -3020 13180 -2940
rect 13260 -3020 13300 -2940
rect 13380 -3020 13420 -2940
rect 13500 -3020 13540 -2940
rect 13620 -3020 13660 -2940
rect 13740 -3020 13780 -2940
rect 13860 -3020 13900 -2940
rect 13980 -3020 14020 -2940
rect 14100 -3020 14140 -2940
rect 14220 -3020 14260 -2940
rect 14340 -3020 14380 -2940
rect 14460 -3020 14500 -2940
rect 14580 -3020 14620 -2940
rect 14700 -3020 14740 -2940
rect 14820 -3020 14860 -2940
rect 14940 -3020 14980 -2940
rect 15060 -3020 15100 -2940
rect 15180 -3020 15220 -2940
rect 15300 -3020 15340 -2940
rect 15420 -3020 15460 -2940
rect 15540 -3020 15580 -2940
rect 15660 -3020 15680 -2940
rect 11120 -3080 15680 -3020
rect 11120 -3160 11140 -3080
rect 11220 -3160 11260 -3080
rect 11340 -3160 11380 -3080
rect 11460 -3160 11500 -3080
rect 11580 -3160 11620 -3080
rect 11700 -3160 11740 -3080
rect 11820 -3160 11860 -3080
rect 11940 -3160 11980 -3080
rect 12060 -3160 12100 -3080
rect 12180 -3160 12220 -3080
rect 12300 -3160 12340 -3080
rect 12420 -3160 12460 -3080
rect 12540 -3160 12580 -3080
rect 12660 -3160 12700 -3080
rect 12780 -3160 12820 -3080
rect 12900 -3160 12940 -3080
rect 13020 -3160 13060 -3080
rect 13140 -3160 13180 -3080
rect 13260 -3160 13300 -3080
rect 13380 -3160 13420 -3080
rect 13500 -3160 13540 -3080
rect 13620 -3160 13660 -3080
rect 13740 -3160 13780 -3080
rect 13860 -3160 13900 -3080
rect 13980 -3160 14020 -3080
rect 14100 -3160 14140 -3080
rect 14220 -3160 14260 -3080
rect 14340 -3160 14380 -3080
rect 14460 -3160 14500 -3080
rect 14580 -3160 14620 -3080
rect 14700 -3160 14740 -3080
rect 14820 -3160 14860 -3080
rect 14940 -3160 14980 -3080
rect 15060 -3160 15100 -3080
rect 15180 -3160 15220 -3080
rect 15300 -3160 15340 -3080
rect 15420 -3160 15460 -3080
rect 15540 -3160 15580 -3080
rect 15660 -3160 15680 -3080
rect 16820 -2880 16940 -2860
rect 16820 -2940 16840 -2880
rect 16900 -2940 16940 -2880
rect 16820 -3060 16940 -2940
rect 16820 -3120 16840 -3060
rect 16900 -3120 16940 -3060
rect 16820 -3140 16940 -3120
rect 17420 -2880 17540 -2860
rect 17420 -2940 17440 -2880
rect 17500 -2940 17540 -2880
rect 17420 -3060 17540 -2940
rect 17420 -3120 17440 -3060
rect 17500 -3120 17540 -3060
rect 17420 -3140 17540 -3120
rect 18040 -2880 18160 -2860
rect 18040 -2940 18080 -2880
rect 18140 -2940 18160 -2880
rect 18040 -3060 18160 -2940
rect 18040 -3120 18080 -3060
rect 18140 -3120 18160 -3060
rect 18040 -3140 18160 -3120
rect 18660 -2880 18780 -2860
rect 18660 -2940 18680 -2880
rect 18740 -2940 18780 -2880
rect 18660 -3060 18780 -2940
rect 18660 -3120 18680 -3060
rect 18740 -3120 18780 -3060
rect 18660 -3140 18780 -3120
rect 19280 -2880 19400 -2860
rect 19280 -2940 19300 -2880
rect 19360 -2940 19400 -2880
rect 19280 -3060 19400 -2940
rect 19280 -3120 19300 -3060
rect 19360 -3120 19400 -3060
rect 19280 -3140 19400 -3120
rect 11120 -3220 15680 -3160
rect 7460 -3420 9880 -3260
rect 11120 -3300 11140 -3220
rect 11220 -3300 11260 -3220
rect 11340 -3300 11380 -3220
rect 11460 -3300 11500 -3220
rect 11580 -3300 11620 -3220
rect 11700 -3300 11740 -3220
rect 11820 -3300 11860 -3220
rect 11940 -3300 11980 -3220
rect 12060 -3300 12100 -3220
rect 12180 -3300 12220 -3220
rect 12300 -3300 12340 -3220
rect 12420 -3300 12460 -3220
rect 12540 -3300 12580 -3220
rect 12660 -3300 12700 -3220
rect 12780 -3300 12820 -3220
rect 12900 -3300 12940 -3220
rect 13020 -3300 13060 -3220
rect 13140 -3300 13180 -3220
rect 13260 -3300 13300 -3220
rect 13380 -3300 13420 -3220
rect 13500 -3300 13540 -3220
rect 13620 -3300 13660 -3220
rect 13740 -3300 13780 -3220
rect 13860 -3300 13900 -3220
rect 13980 -3300 14020 -3220
rect 14100 -3300 14140 -3220
rect 14220 -3300 14260 -3220
rect 14340 -3300 14380 -3220
rect 14460 -3300 14500 -3220
rect 14580 -3300 14620 -3220
rect 14700 -3300 14740 -3220
rect 14820 -3300 14860 -3220
rect 14940 -3300 14980 -3220
rect 15060 -3300 15100 -3220
rect 15180 -3300 15220 -3220
rect 15300 -3300 15340 -3220
rect 15420 -3300 15460 -3220
rect 15540 -3300 15580 -3220
rect 15660 -3300 15680 -3220
rect 11120 -3320 15680 -3300
rect 7460 -3500 7480 -3420
rect 7560 -3500 7580 -3420
rect 7660 -3500 7680 -3420
rect 7760 -3500 7780 -3420
rect 7860 -3500 7880 -3420
rect 7960 -3500 7980 -3420
rect 8060 -3500 8080 -3420
rect 8160 -3500 8180 -3420
rect 8260 -3500 8280 -3420
rect 8360 -3500 8380 -3420
rect 8460 -3500 8480 -3420
rect 8560 -3500 8580 -3420
rect 8660 -3500 8680 -3420
rect 8760 -3500 8780 -3420
rect 8860 -3500 8880 -3420
rect 8960 -3500 8980 -3420
rect 9060 -3500 9080 -3420
rect 9160 -3500 9180 -3420
rect 9260 -3500 9280 -3420
rect 9360 -3500 9380 -3420
rect 9460 -3500 9480 -3420
rect 9560 -3500 9580 -3420
rect 9660 -3500 9680 -3420
rect 9760 -3500 9780 -3420
rect 9860 -3500 9880 -3420
rect 7460 -3560 9880 -3500
rect 7460 -3640 7480 -3560
rect 7560 -3640 7580 -3560
rect 7660 -3640 7680 -3560
rect 7760 -3640 7780 -3560
rect 7860 -3640 7880 -3560
rect 7960 -3640 7980 -3560
rect 8060 -3640 8080 -3560
rect 8160 -3640 8180 -3560
rect 8260 -3640 8280 -3560
rect 8360 -3640 8380 -3560
rect 8460 -3640 8480 -3560
rect 8560 -3640 8580 -3560
rect 8660 -3640 8680 -3560
rect 8760 -3640 8780 -3560
rect 8860 -3640 8880 -3560
rect 8960 -3640 8980 -3560
rect 9060 -3640 9080 -3560
rect 9160 -3640 9180 -3560
rect 9260 -3640 9280 -3560
rect 9360 -3640 9380 -3560
rect 9460 -3640 9480 -3560
rect 9560 -3640 9580 -3560
rect 9660 -3640 9680 -3560
rect 9760 -3640 9780 -3560
rect 9860 -3640 9880 -3560
rect 7460 -3700 9880 -3640
rect 7460 -3780 7480 -3700
rect 7560 -3780 7580 -3700
rect 7660 -3780 7680 -3700
rect 7760 -3780 7780 -3700
rect 7860 -3780 7880 -3700
rect 7960 -3780 7980 -3700
rect 8060 -3780 8080 -3700
rect 8160 -3780 8180 -3700
rect 8260 -3780 8280 -3700
rect 8360 -3780 8380 -3700
rect 8460 -3780 8480 -3700
rect 8560 -3780 8580 -3700
rect 8660 -3780 8680 -3700
rect 8760 -3780 8780 -3700
rect 8860 -3780 8880 -3700
rect 8960 -3780 8980 -3700
rect 9060 -3780 9080 -3700
rect 9160 -3780 9180 -3700
rect 9260 -3780 9280 -3700
rect 9360 -3780 9380 -3700
rect 9460 -3780 9480 -3700
rect 9560 -3780 9580 -3700
rect 9660 -3780 9680 -3700
rect 9760 -3780 9780 -3700
rect 9860 -3780 9880 -3700
rect 7460 -3800 9880 -3780
rect 16900 -3420 19320 -3260
rect 16900 -3500 16920 -3420
rect 17000 -3500 17020 -3420
rect 17100 -3500 17120 -3420
rect 17200 -3500 17220 -3420
rect 17300 -3500 17320 -3420
rect 17400 -3500 17420 -3420
rect 17500 -3500 17520 -3420
rect 17600 -3500 17620 -3420
rect 17700 -3500 17720 -3420
rect 17800 -3500 17820 -3420
rect 17900 -3500 17920 -3420
rect 18000 -3500 18020 -3420
rect 18100 -3500 18120 -3420
rect 18200 -3500 18220 -3420
rect 18300 -3500 18320 -3420
rect 18400 -3500 18420 -3420
rect 18500 -3500 18520 -3420
rect 18600 -3500 18620 -3420
rect 18700 -3500 18720 -3420
rect 18800 -3500 18820 -3420
rect 18900 -3500 18920 -3420
rect 19000 -3500 19020 -3420
rect 19100 -3500 19120 -3420
rect 19200 -3500 19220 -3420
rect 19300 -3500 19320 -3420
rect 16900 -3560 19320 -3500
rect 16900 -3640 16920 -3560
rect 17000 -3640 17020 -3560
rect 17100 -3640 17120 -3560
rect 17200 -3640 17220 -3560
rect 17300 -3640 17320 -3560
rect 17400 -3640 17420 -3560
rect 17500 -3640 17520 -3560
rect 17600 -3640 17620 -3560
rect 17700 -3640 17720 -3560
rect 17800 -3640 17820 -3560
rect 17900 -3640 17920 -3560
rect 18000 -3640 18020 -3560
rect 18100 -3640 18120 -3560
rect 18200 -3640 18220 -3560
rect 18300 -3640 18320 -3560
rect 18400 -3640 18420 -3560
rect 18500 -3640 18520 -3560
rect 18600 -3640 18620 -3560
rect 18700 -3640 18720 -3560
rect 18800 -3640 18820 -3560
rect 18900 -3640 18920 -3560
rect 19000 -3640 19020 -3560
rect 19100 -3640 19120 -3560
rect 19200 -3640 19220 -3560
rect 19300 -3640 19320 -3560
rect 16900 -3700 19320 -3640
rect 16900 -3780 16920 -3700
rect 17000 -3780 17020 -3700
rect 17100 -3780 17120 -3700
rect 17200 -3780 17220 -3700
rect 17300 -3780 17320 -3700
rect 17400 -3780 17420 -3700
rect 17500 -3780 17520 -3700
rect 17600 -3780 17620 -3700
rect 17700 -3780 17720 -3700
rect 17800 -3780 17820 -3700
rect 17900 -3780 17920 -3700
rect 18000 -3780 18020 -3700
rect 18100 -3780 18120 -3700
rect 18200 -3780 18220 -3700
rect 18300 -3780 18320 -3700
rect 18400 -3780 18420 -3700
rect 18500 -3780 18520 -3700
rect 18600 -3780 18620 -3700
rect 18700 -3780 18720 -3700
rect 18800 -3780 18820 -3700
rect 18900 -3780 18920 -3700
rect 19000 -3780 19020 -3700
rect 19100 -3780 19120 -3700
rect 19200 -3780 19220 -3700
rect 19300 -3780 19320 -3700
rect 16900 -3800 19320 -3780
rect 13200 -3900 13600 -3880
rect 8320 -3960 8460 -3940
rect 8320 -4020 8360 -3960
rect 8420 -4020 8460 -3960
rect 8320 -4140 8460 -4020
rect 8320 -4200 8360 -4140
rect 8420 -4200 8460 -4140
rect 8320 -4220 8460 -4200
rect 8780 -3960 8920 -3940
rect 8780 -4020 8820 -3960
rect 8880 -4020 8920 -3960
rect 13200 -3980 13220 -3900
rect 13300 -3980 13360 -3900
rect 13440 -3980 13500 -3900
rect 13580 -3980 13600 -3900
rect 17940 -3960 18080 -3940
rect 8780 -4140 8920 -4020
rect 8780 -4200 8820 -4140
rect 8880 -4200 8920 -4140
rect 8780 -4220 8920 -4200
rect 10420 -4060 12360 -3980
rect 10420 -4080 11360 -4060
rect 8560 -4440 8700 -4420
rect 8560 -4500 8620 -4440
rect 8680 -4500 8700 -4440
rect 8560 -4540 8700 -4500
rect 8560 -4600 8620 -4540
rect 8680 -4600 8700 -4540
rect 8560 -4620 8700 -4600
rect 10280 -4440 10380 -4420
rect 10280 -4500 10300 -4440
rect 10360 -4500 10380 -4440
rect 10280 -4520 10380 -4500
rect 10280 -4580 10300 -4520
rect 10360 -4580 10380 -4520
rect 10280 -4600 10380 -4580
rect 10280 -4660 10300 -4600
rect 10360 -4660 10380 -4600
rect 10280 -4680 10380 -4660
rect 8420 -5380 8840 -4960
rect 10420 -5060 10560 -4080
rect 11320 -4140 11360 -4080
rect 11440 -4080 12360 -4060
rect 11440 -4140 11480 -4080
rect 11320 -4180 11480 -4140
rect 11320 -4260 11360 -4180
rect 11440 -4260 11480 -4180
rect 11320 -4300 11480 -4260
rect 11320 -4380 11360 -4300
rect 11440 -4380 11480 -4300
rect 11320 -4420 11480 -4380
rect 10600 -4440 10700 -4420
rect 10600 -4500 10620 -4440
rect 10680 -4500 10700 -4440
rect 10600 -4520 10700 -4500
rect 10600 -4580 10620 -4520
rect 10680 -4580 10700 -4520
rect 10600 -4600 10700 -4580
rect 10600 -4660 10620 -4600
rect 10680 -4660 10700 -4600
rect 10600 -4680 10700 -4660
rect 11320 -4500 11360 -4420
rect 11440 -4500 11480 -4420
rect 11320 -4540 11480 -4500
rect 11320 -4620 11360 -4540
rect 11440 -4620 11480 -4540
rect 11320 -4660 11480 -4620
rect 11320 -4740 11360 -4660
rect 11440 -4740 11480 -4660
rect 12080 -4440 12180 -4420
rect 12080 -4500 12100 -4440
rect 12160 -4500 12180 -4440
rect 12080 -4520 12180 -4500
rect 12080 -4580 12100 -4520
rect 12160 -4580 12180 -4520
rect 12080 -4600 12180 -4580
rect 12080 -4660 12100 -4600
rect 12160 -4660 12180 -4600
rect 12080 -4680 12180 -4660
rect 11320 -4780 11480 -4740
rect 11320 -4860 11360 -4780
rect 11440 -4860 11480 -4780
rect 11320 -4900 11480 -4860
rect 11320 -4980 11360 -4900
rect 11440 -4980 11480 -4900
rect 11320 -5020 11480 -4980
rect 11320 -5100 11360 -5020
rect 11440 -5100 11480 -5020
rect 12220 -5060 12360 -4080
rect 13200 -4020 13600 -3980
rect 13200 -4100 13220 -4020
rect 13300 -4100 13360 -4020
rect 13440 -4100 13500 -4020
rect 13580 -4100 13600 -4020
rect 13200 -4140 13600 -4100
rect 13200 -4220 13220 -4140
rect 13300 -4220 13360 -4140
rect 13440 -4220 13500 -4140
rect 13580 -4220 13600 -4140
rect 13200 -4260 13600 -4220
rect 13200 -4340 13220 -4260
rect 13300 -4340 13360 -4260
rect 13440 -4340 13500 -4260
rect 13580 -4340 13600 -4260
rect 13200 -4380 13600 -4340
rect 12400 -4440 12500 -4420
rect 12400 -4500 12420 -4440
rect 12480 -4500 12500 -4440
rect 12400 -4520 12500 -4500
rect 12400 -4580 12420 -4520
rect 12480 -4580 12500 -4520
rect 12400 -4600 12500 -4580
rect 12400 -4660 12420 -4600
rect 12480 -4660 12500 -4600
rect 12400 -4680 12500 -4660
rect 13200 -4460 13220 -4380
rect 13300 -4460 13360 -4380
rect 13440 -4460 13500 -4380
rect 13580 -4460 13600 -4380
rect 14420 -4060 16360 -3980
rect 14420 -4080 15360 -4060
rect 13200 -4500 13600 -4460
rect 13200 -4580 13220 -4500
rect 13300 -4580 13360 -4500
rect 13440 -4580 13500 -4500
rect 13580 -4580 13600 -4500
rect 13200 -4620 13600 -4580
rect 13200 -4700 13220 -4620
rect 13300 -4700 13360 -4620
rect 13440 -4700 13500 -4620
rect 13580 -4700 13600 -4620
rect 14280 -4440 14380 -4420
rect 14280 -4500 14300 -4440
rect 14360 -4500 14380 -4440
rect 14280 -4520 14380 -4500
rect 14280 -4580 14300 -4520
rect 14360 -4580 14380 -4520
rect 14280 -4600 14380 -4580
rect 14280 -4660 14300 -4600
rect 14360 -4660 14380 -4600
rect 14280 -4680 14380 -4660
rect 13200 -4740 13600 -4700
rect 13200 -4820 13220 -4740
rect 13300 -4820 13360 -4740
rect 13440 -4820 13500 -4740
rect 13580 -4820 13600 -4740
rect 13200 -4860 13600 -4820
rect 13200 -4940 13220 -4860
rect 13300 -4940 13360 -4860
rect 13440 -4940 13500 -4860
rect 13580 -4940 13600 -4860
rect 13200 -4980 13600 -4940
rect 13200 -5060 13220 -4980
rect 13300 -5060 13360 -4980
rect 13440 -5060 13500 -4980
rect 13580 -5060 13600 -4980
rect 14420 -5060 14560 -4080
rect 15320 -4140 15360 -4080
rect 15440 -4080 16360 -4060
rect 15440 -4140 15480 -4080
rect 15320 -4180 15480 -4140
rect 15320 -4260 15360 -4180
rect 15440 -4260 15480 -4180
rect 15320 -4300 15480 -4260
rect 15320 -4380 15360 -4300
rect 15440 -4380 15480 -4300
rect 15320 -4420 15480 -4380
rect 14600 -4440 14700 -4420
rect 14600 -4500 14620 -4440
rect 14680 -4500 14700 -4440
rect 14600 -4520 14700 -4500
rect 14600 -4580 14620 -4520
rect 14680 -4580 14700 -4520
rect 14600 -4600 14700 -4580
rect 14600 -4660 14620 -4600
rect 14680 -4660 14700 -4600
rect 14600 -4680 14700 -4660
rect 15320 -4500 15360 -4420
rect 15440 -4500 15480 -4420
rect 15320 -4540 15480 -4500
rect 15320 -4620 15360 -4540
rect 15440 -4620 15480 -4540
rect 15320 -4660 15480 -4620
rect 15320 -4740 15360 -4660
rect 15440 -4740 15480 -4660
rect 16080 -4440 16180 -4420
rect 16080 -4500 16100 -4440
rect 16160 -4500 16180 -4440
rect 16080 -4520 16180 -4500
rect 16080 -4580 16100 -4520
rect 16160 -4580 16180 -4520
rect 16080 -4600 16180 -4580
rect 16080 -4660 16100 -4600
rect 16160 -4660 16180 -4600
rect 16080 -4680 16180 -4660
rect 15320 -4780 15480 -4740
rect 15320 -4860 15360 -4780
rect 15440 -4860 15480 -4780
rect 15320 -4900 15480 -4860
rect 15320 -4980 15360 -4900
rect 15440 -4980 15480 -4900
rect 15320 -5020 15480 -4980
rect 13200 -5100 13600 -5060
rect 15320 -5100 15360 -5020
rect 15440 -5100 15480 -5020
rect 16220 -5060 16360 -4080
rect 17940 -4020 17960 -3960
rect 18020 -4020 18080 -3960
rect 17940 -4140 18080 -4020
rect 17940 -4200 17960 -4140
rect 18020 -4200 18080 -4140
rect 17940 -4220 18080 -4200
rect 18380 -3960 18520 -3940
rect 18380 -4020 18420 -3960
rect 18480 -4020 18520 -3960
rect 18380 -4140 18520 -4020
rect 18380 -4200 18420 -4140
rect 18480 -4200 18520 -4140
rect 18380 -4220 18520 -4200
rect 16400 -4440 16500 -4420
rect 16400 -4500 16420 -4440
rect 16480 -4500 16500 -4440
rect 16400 -4520 16500 -4500
rect 16400 -4580 16420 -4520
rect 16480 -4580 16500 -4520
rect 16400 -4600 16500 -4580
rect 16400 -4660 16420 -4600
rect 16480 -4660 16500 -4600
rect 18120 -4440 18260 -4420
rect 18120 -4500 18140 -4440
rect 18200 -4500 18260 -4440
rect 18120 -4540 18260 -4500
rect 18120 -4600 18140 -4540
rect 18200 -4600 18260 -4540
rect 18120 -4620 18260 -4600
rect 16400 -4680 16500 -4660
rect 10360 -5120 10620 -5100
rect 10360 -5180 10380 -5120
rect 10440 -5180 10540 -5120
rect 10600 -5180 10620 -5120
rect 10360 -5240 10620 -5180
rect 11320 -5140 11480 -5100
rect 11320 -5220 11360 -5140
rect 11440 -5220 11480 -5140
rect 11320 -5260 11480 -5220
rect 12160 -5120 12420 -5100
rect 12160 -5180 12180 -5120
rect 12240 -5180 12340 -5120
rect 12400 -5180 12420 -5120
rect 12160 -5240 12420 -5180
rect 13200 -5180 13220 -5100
rect 13300 -5180 13360 -5100
rect 13440 -5180 13500 -5100
rect 13580 -5180 13600 -5100
rect 13200 -5220 13600 -5180
rect 11320 -5320 11360 -5260
rect 8420 -5460 8440 -5380
rect 8520 -5460 8580 -5380
rect 8680 -5460 8740 -5380
rect 8820 -5460 8840 -5380
rect 8420 -5500 8840 -5460
rect 9720 -5340 11360 -5320
rect 11440 -5320 11480 -5260
rect 13200 -5300 13220 -5220
rect 13300 -5300 13360 -5220
rect 13440 -5300 13500 -5220
rect 13580 -5300 13600 -5220
rect 14360 -5120 14620 -5100
rect 14360 -5180 14380 -5120
rect 14440 -5180 14540 -5120
rect 14600 -5180 14620 -5120
rect 14360 -5240 14620 -5180
rect 15320 -5140 15480 -5100
rect 15320 -5220 15360 -5140
rect 15440 -5220 15480 -5140
rect 13200 -5320 13600 -5300
rect 15320 -5260 15480 -5220
rect 16160 -5120 16420 -5110
rect 16160 -5180 16180 -5120
rect 16240 -5180 16340 -5120
rect 16400 -5180 16420 -5120
rect 16160 -5250 16420 -5180
rect 15320 -5320 15360 -5260
rect 11440 -5340 15360 -5320
rect 15440 -5320 15480 -5260
rect 15440 -5340 17080 -5320
rect 9720 -5420 9740 -5340
rect 9820 -5420 9860 -5340
rect 9940 -5420 9980 -5340
rect 10060 -5420 10100 -5340
rect 10180 -5420 10220 -5340
rect 10300 -5420 10340 -5340
rect 10420 -5420 10460 -5340
rect 10540 -5420 10580 -5340
rect 10660 -5420 10700 -5340
rect 10780 -5420 10820 -5340
rect 10900 -5420 10940 -5340
rect 11020 -5420 11060 -5340
rect 11140 -5420 11180 -5340
rect 11260 -5380 11540 -5340
rect 11260 -5420 11360 -5380
rect 9720 -5460 11360 -5420
rect 11440 -5420 11540 -5380
rect 11620 -5420 11660 -5340
rect 11740 -5420 11780 -5340
rect 11860 -5420 11900 -5340
rect 11980 -5420 12020 -5340
rect 12100 -5420 12140 -5340
rect 12220 -5420 12260 -5340
rect 12340 -5420 12380 -5340
rect 12460 -5420 12500 -5340
rect 12580 -5420 12620 -5340
rect 12700 -5420 12740 -5340
rect 12820 -5420 12860 -5340
rect 12940 -5420 12980 -5340
rect 13060 -5420 13100 -5340
rect 13180 -5420 13220 -5340
rect 13300 -5420 13360 -5340
rect 13440 -5420 13500 -5340
rect 13580 -5420 13620 -5340
rect 13700 -5420 13740 -5340
rect 13820 -5420 13860 -5340
rect 13940 -5420 13980 -5340
rect 14060 -5420 14100 -5340
rect 14180 -5420 14220 -5340
rect 14300 -5420 14340 -5340
rect 14420 -5420 14460 -5340
rect 14540 -5420 14580 -5340
rect 14660 -5420 14700 -5340
rect 14780 -5420 14820 -5340
rect 14900 -5420 14940 -5340
rect 15020 -5420 15060 -5340
rect 15140 -5420 15180 -5340
rect 15260 -5380 15540 -5340
rect 15260 -5420 15360 -5380
rect 11440 -5460 15360 -5420
rect 15440 -5420 15540 -5380
rect 15620 -5420 15660 -5340
rect 15740 -5420 15780 -5340
rect 15860 -5420 15900 -5340
rect 15980 -5420 16020 -5340
rect 16100 -5420 16140 -5340
rect 16220 -5420 16260 -5340
rect 16340 -5420 16380 -5340
rect 16460 -5420 16500 -5340
rect 16580 -5420 16620 -5340
rect 16700 -5420 16740 -5340
rect 16820 -5420 16860 -5340
rect 16940 -5420 16980 -5340
rect 17060 -5420 17080 -5340
rect 15440 -5460 17080 -5420
rect 9720 -5480 13220 -5460
rect 9720 -5560 9740 -5480
rect 9820 -5560 9860 -5480
rect 9940 -5560 9980 -5480
rect 10060 -5560 10100 -5480
rect 10180 -5560 10220 -5480
rect 10300 -5560 10340 -5480
rect 10420 -5560 10460 -5480
rect 10540 -5560 10580 -5480
rect 10660 -5560 10700 -5480
rect 10780 -5560 10820 -5480
rect 10900 -5560 10940 -5480
rect 11020 -5560 11060 -5480
rect 11140 -5560 11180 -5480
rect 11260 -5500 11540 -5480
rect 11260 -5560 11360 -5500
rect 9720 -5580 11360 -5560
rect 11440 -5560 11540 -5500
rect 11620 -5560 11660 -5480
rect 11740 -5560 11780 -5480
rect 11860 -5560 11900 -5480
rect 11980 -5560 12020 -5480
rect 12100 -5560 12140 -5480
rect 12220 -5560 12260 -5480
rect 12340 -5560 12380 -5480
rect 12460 -5560 12500 -5480
rect 12580 -5560 12620 -5480
rect 12700 -5560 12740 -5480
rect 12820 -5560 12860 -5480
rect 12940 -5560 12980 -5480
rect 13060 -5560 13100 -5480
rect 13180 -5540 13220 -5480
rect 13300 -5540 13360 -5460
rect 13440 -5540 13500 -5460
rect 13580 -5480 17080 -5460
rect 13580 -5540 13620 -5480
rect 13180 -5560 13620 -5540
rect 13700 -5560 13740 -5480
rect 13820 -5560 13860 -5480
rect 13940 -5560 13980 -5480
rect 14060 -5560 14100 -5480
rect 14180 -5560 14220 -5480
rect 14300 -5560 14340 -5480
rect 14420 -5560 14460 -5480
rect 14540 -5560 14580 -5480
rect 14660 -5560 14700 -5480
rect 14780 -5560 14820 -5480
rect 14900 -5560 14940 -5480
rect 15020 -5560 15060 -5480
rect 15140 -5560 15180 -5480
rect 15260 -5500 15540 -5480
rect 15260 -5560 15360 -5500
rect 11440 -5580 15360 -5560
rect 15440 -5560 15540 -5500
rect 15620 -5560 15660 -5480
rect 15740 -5560 15780 -5480
rect 15860 -5560 15900 -5480
rect 15980 -5560 16020 -5480
rect 16100 -5560 16140 -5480
rect 16220 -5560 16260 -5480
rect 16340 -5560 16380 -5480
rect 16460 -5560 16500 -5480
rect 16580 -5560 16620 -5480
rect 16700 -5560 16740 -5480
rect 16820 -5560 16860 -5480
rect 16940 -5560 16980 -5480
rect 17060 -5560 17080 -5480
rect 18000 -5380 18420 -4960
rect 18000 -5460 18020 -5380
rect 18100 -5460 18140 -5380
rect 18280 -5460 18320 -5380
rect 18400 -5460 18420 -5380
rect 18000 -5500 18420 -5460
rect 15440 -5580 17080 -5560
rect 11320 -5620 11480 -5580
rect 10360 -5720 10620 -5650
rect 10360 -5780 10380 -5720
rect 10440 -5780 10540 -5720
rect 10600 -5780 10620 -5720
rect 10360 -5790 10620 -5780
rect 11320 -5700 11360 -5620
rect 11440 -5700 11480 -5620
rect 11320 -5740 11480 -5700
rect 11320 -5820 11360 -5740
rect 11440 -5820 11480 -5740
rect 12160 -5720 12420 -5650
rect 12160 -5780 12180 -5720
rect 12240 -5780 12340 -5720
rect 12400 -5780 12420 -5720
rect 12160 -5790 12420 -5780
rect 13200 -5660 13220 -5580
rect 13300 -5660 13360 -5580
rect 13440 -5660 13500 -5580
rect 13580 -5660 13600 -5580
rect 15320 -5620 15480 -5580
rect 13200 -5700 13600 -5660
rect 13200 -5780 13220 -5700
rect 13300 -5780 13360 -5700
rect 13440 -5780 13500 -5700
rect 13580 -5780 13600 -5700
rect 10280 -5940 10380 -5920
rect 7860 -5960 8040 -5940
rect 7860 -6020 7920 -5960
rect 7980 -6020 8040 -5960
rect 7860 -6140 8040 -6020
rect 7860 -6200 7920 -6140
rect 7980 -6200 8040 -6140
rect 7860 -6220 8040 -6200
rect 8480 -5960 8660 -5940
rect 8480 -6020 8540 -5960
rect 8600 -6020 8660 -5960
rect 8480 -6140 8660 -6020
rect 8480 -6200 8540 -6140
rect 8600 -6200 8660 -6140
rect 8480 -6220 8660 -6200
rect 9100 -5960 9280 -5940
rect 9100 -6020 9140 -5960
rect 9200 -6020 9280 -5960
rect 9100 -6140 9280 -6020
rect 9100 -6200 9140 -6140
rect 9200 -6200 9280 -6140
rect 10280 -6000 10300 -5940
rect 10360 -6000 10380 -5940
rect 10280 -6020 10380 -6000
rect 10280 -6080 10300 -6020
rect 10360 -6080 10380 -6020
rect 10280 -6100 10380 -6080
rect 10280 -6160 10300 -6100
rect 10360 -6160 10380 -6100
rect 10280 -6180 10380 -6160
rect 9100 -6220 9280 -6200
rect 10420 -6820 10560 -5840
rect 11320 -5860 11480 -5820
rect 13200 -5820 13600 -5780
rect 14360 -5720 14620 -5650
rect 14360 -5780 14380 -5720
rect 14440 -5780 14540 -5720
rect 14600 -5780 14620 -5720
rect 14360 -5790 14620 -5780
rect 15320 -5700 15360 -5620
rect 15440 -5700 15480 -5620
rect 15320 -5740 15480 -5700
rect 10600 -5940 10700 -5920
rect 10600 -6000 10620 -5940
rect 10680 -6000 10700 -5940
rect 10600 -6020 10700 -6000
rect 10600 -6080 10620 -6020
rect 10680 -6080 10700 -6020
rect 10600 -6100 10700 -6080
rect 10600 -6160 10620 -6100
rect 10680 -6160 10700 -6100
rect 10600 -6180 10700 -6160
rect 11320 -5940 11360 -5860
rect 11440 -5940 11480 -5860
rect 11320 -5980 11480 -5940
rect 11320 -6060 11360 -5980
rect 11440 -6060 11480 -5980
rect 11320 -6100 11480 -6060
rect 11320 -6180 11360 -6100
rect 11440 -6180 11480 -6100
rect 11320 -6220 11480 -6180
rect 11320 -6300 11360 -6220
rect 11440 -6300 11480 -6220
rect 11320 -6340 11480 -6300
rect 11320 -6420 11360 -6340
rect 11440 -6420 11480 -6340
rect 11320 -6460 11480 -6420
rect 11320 -6540 11360 -6460
rect 11440 -6540 11480 -6460
rect 11320 -6580 11480 -6540
rect 11320 -6660 11360 -6580
rect 11440 -6660 11480 -6580
rect 11320 -6700 11480 -6660
rect 11320 -6780 11360 -6700
rect 11440 -6780 11480 -6700
rect 12080 -6540 12180 -6520
rect 12080 -6600 12100 -6540
rect 12160 -6600 12180 -6540
rect 12080 -6620 12180 -6600
rect 12080 -6680 12100 -6620
rect 12160 -6680 12180 -6620
rect 12080 -6700 12180 -6680
rect 12080 -6760 12100 -6700
rect 12160 -6760 12180 -6700
rect 12080 -6780 12180 -6760
rect 11320 -6820 11480 -6780
rect 12220 -6820 12360 -5840
rect 13200 -5900 13220 -5820
rect 13300 -5900 13360 -5820
rect 13440 -5900 13500 -5820
rect 13580 -5900 13600 -5820
rect 15320 -5820 15360 -5740
rect 15440 -5820 15480 -5740
rect 16160 -5720 16420 -5650
rect 16160 -5780 16180 -5720
rect 16240 -5780 16340 -5720
rect 16400 -5780 16420 -5720
rect 16160 -5790 16420 -5780
rect 13200 -5940 13600 -5900
rect 13200 -6020 13220 -5940
rect 13300 -6020 13360 -5940
rect 13440 -6020 13500 -5940
rect 13580 -6020 13600 -5940
rect 13200 -6060 13600 -6020
rect 13200 -6140 13220 -6060
rect 13300 -6140 13360 -6060
rect 13440 -6140 13500 -6060
rect 13580 -6140 13600 -6060
rect 13200 -6180 13600 -6140
rect 13200 -6260 13220 -6180
rect 13300 -6260 13360 -6180
rect 13440 -6260 13500 -6180
rect 13580 -6260 13600 -6180
rect 13200 -6300 13600 -6260
rect 13200 -6380 13220 -6300
rect 13300 -6380 13360 -6300
rect 13440 -6380 13500 -6300
rect 13580 -6380 13600 -6300
rect 13200 -6420 13600 -6380
rect 13200 -6500 13220 -6420
rect 13300 -6500 13360 -6420
rect 13440 -6500 13500 -6420
rect 13580 -6500 13600 -6420
rect 12400 -6540 12500 -6520
rect 12400 -6600 12420 -6540
rect 12480 -6600 12500 -6540
rect 12400 -6620 12500 -6600
rect 12400 -6680 12420 -6620
rect 12480 -6680 12500 -6620
rect 12400 -6700 12500 -6680
rect 12400 -6760 12420 -6700
rect 12480 -6760 12500 -6700
rect 12400 -6780 12500 -6760
rect 13200 -6540 13600 -6500
rect 13200 -6620 13220 -6540
rect 13300 -6620 13360 -6540
rect 13440 -6620 13500 -6540
rect 13580 -6620 13600 -6540
rect 13200 -6660 13600 -6620
rect 13200 -6740 13220 -6660
rect 13300 -6740 13360 -6660
rect 13440 -6740 13500 -6660
rect 13580 -6740 13600 -6660
rect 13200 -6780 13600 -6740
rect 14280 -6540 14380 -6520
rect 14280 -6600 14300 -6540
rect 14360 -6600 14380 -6540
rect 14280 -6620 14380 -6600
rect 14280 -6680 14300 -6620
rect 14360 -6680 14380 -6620
rect 14280 -6700 14380 -6680
rect 14280 -6760 14300 -6700
rect 14360 -6760 14380 -6700
rect 14280 -6780 14380 -6760
rect 10420 -6920 12360 -6820
rect 13200 -6860 13220 -6780
rect 13300 -6860 13360 -6780
rect 13440 -6860 13500 -6780
rect 13580 -6860 13600 -6780
rect 13200 -6900 13600 -6860
rect 13200 -6980 13220 -6900
rect 13300 -6980 13360 -6900
rect 13440 -6980 13500 -6900
rect 13580 -6980 13600 -6900
rect 14420 -6820 14560 -5840
rect 15320 -5860 15480 -5820
rect 15040 -6180 15140 -5920
rect 15320 -5940 15360 -5860
rect 15440 -5940 15480 -5860
rect 15320 -5980 15480 -5940
rect 15320 -6060 15360 -5980
rect 15440 -6060 15480 -5980
rect 15320 -6100 15480 -6060
rect 15320 -6180 15360 -6100
rect 15440 -6180 15480 -6100
rect 16080 -5940 16180 -5920
rect 16080 -6000 16100 -5940
rect 16160 -6000 16180 -5940
rect 16080 -6020 16180 -6000
rect 16080 -6080 16100 -6020
rect 16160 -6080 16180 -6020
rect 16080 -6100 16180 -6080
rect 16080 -6160 16100 -6100
rect 16160 -6160 16180 -6100
rect 16080 -6180 16180 -6160
rect 15320 -6220 15480 -6180
rect 15320 -6300 15360 -6220
rect 15440 -6300 15480 -6220
rect 15320 -6340 15480 -6300
rect 15320 -6420 15360 -6340
rect 15440 -6420 15480 -6340
rect 15320 -6460 15480 -6420
rect 14600 -6540 14700 -6520
rect 14600 -6600 14620 -6540
rect 14680 -6600 14700 -6540
rect 14600 -6620 14700 -6600
rect 14600 -6680 14620 -6620
rect 14680 -6680 14700 -6620
rect 14600 -6700 14700 -6680
rect 14600 -6760 14620 -6700
rect 14680 -6760 14700 -6700
rect 14600 -6780 14700 -6760
rect 15320 -6540 15360 -6460
rect 15440 -6540 15480 -6460
rect 15320 -6580 15480 -6540
rect 15320 -6660 15360 -6580
rect 15440 -6660 15480 -6580
rect 15320 -6700 15480 -6660
rect 15320 -6780 15360 -6700
rect 15440 -6780 15480 -6700
rect 15320 -6820 15480 -6780
rect 16220 -6820 16360 -5840
rect 16400 -5940 16500 -5920
rect 16400 -6000 16420 -5940
rect 16480 -6000 16500 -5940
rect 16400 -6020 16500 -6000
rect 16400 -6080 16420 -6020
rect 16480 -6080 16500 -6020
rect 16400 -6100 16500 -6080
rect 16400 -6160 16420 -6100
rect 16480 -6160 16500 -6100
rect 16400 -6180 16500 -6160
rect 17520 -5960 17700 -5940
rect 17520 -6020 17580 -5960
rect 17640 -6020 17700 -5960
rect 17520 -6140 17700 -6020
rect 17520 -6200 17580 -6140
rect 17640 -6200 17700 -6140
rect 17520 -6220 17700 -6200
rect 18160 -5960 18340 -5940
rect 18160 -6020 18200 -5960
rect 18260 -6020 18340 -5960
rect 18160 -6140 18340 -6020
rect 18160 -6200 18200 -6140
rect 18260 -6200 18340 -6140
rect 18160 -6220 18340 -6200
rect 18740 -5960 18920 -5940
rect 18740 -6020 18800 -5960
rect 18860 -6020 18920 -5960
rect 18740 -6140 18920 -6020
rect 18740 -6200 18800 -6140
rect 18860 -6200 18920 -6140
rect 18740 -6220 18920 -6200
rect 14420 -6920 16360 -6820
rect 13200 -7020 13600 -6980
rect 7980 -7480 9160 -7280
rect 7980 -7540 8000 -7480
rect 8060 -7540 8080 -7480
rect 8140 -7540 8160 -7480
rect 8220 -7540 8240 -7480
rect 8300 -7540 8320 -7480
rect 8380 -7540 8400 -7480
rect 8460 -7540 8480 -7480
rect 8540 -7540 8560 -7480
rect 8620 -7540 8640 -7480
rect 8700 -7540 8720 -7480
rect 8780 -7540 8800 -7480
rect 8860 -7540 8880 -7480
rect 8940 -7540 8960 -7480
rect 9060 -7540 9080 -7480
rect 9140 -7540 9160 -7480
rect 7980 -7580 9160 -7540
rect 7980 -7640 8000 -7580
rect 8060 -7640 8080 -7580
rect 8140 -7640 8160 -7580
rect 8220 -7640 8240 -7580
rect 8300 -7640 8320 -7580
rect 8380 -7640 8400 -7580
rect 8460 -7640 8480 -7580
rect 8540 -7640 8560 -7580
rect 8620 -7640 8640 -7580
rect 8700 -7640 8720 -7580
rect 8780 -7640 8800 -7580
rect 8860 -7640 8880 -7580
rect 8940 -7640 8960 -7580
rect 9060 -7640 9080 -7580
rect 9140 -7640 9160 -7580
rect 7980 -7660 9160 -7640
rect 10880 -7480 11040 -7460
rect 10940 -7540 10980 -7480
rect 10880 -7560 11040 -7540
rect 10940 -7620 10980 -7560
rect 10880 -7740 11040 -7620
rect 10940 -7800 10980 -7740
rect 10880 -7820 11040 -7800
rect 10940 -7880 10980 -7820
rect 10880 -7900 11040 -7880
rect 11440 -7500 11620 -7460
rect 11440 -7560 11460 -7500
rect 11520 -7560 11540 -7500
rect 11600 -7560 11620 -7500
rect 11440 -7580 11620 -7560
rect 11440 -7640 11460 -7580
rect 11520 -7640 11540 -7580
rect 11600 -7640 11620 -7580
rect 11440 -7660 11620 -7640
rect 11440 -7720 11460 -7660
rect 11520 -7720 11540 -7660
rect 11600 -7720 11620 -7660
rect 11440 -7740 11620 -7720
rect 11440 -7800 11460 -7740
rect 11520 -7800 11540 -7740
rect 11600 -7800 11620 -7740
rect 11440 -7820 11620 -7800
rect 11440 -7880 11460 -7820
rect 11520 -7880 11540 -7820
rect 11600 -7880 11620 -7820
rect 11440 -7900 11620 -7880
rect 12660 -7500 12840 -7460
rect 12660 -7560 12680 -7500
rect 12740 -7560 12760 -7500
rect 12820 -7560 12840 -7500
rect 12660 -7580 12840 -7560
rect 12660 -7640 12680 -7580
rect 12740 -7640 12760 -7580
rect 12820 -7640 12840 -7580
rect 12660 -7660 12840 -7640
rect 12660 -7720 12680 -7660
rect 12740 -7720 12760 -7660
rect 12820 -7720 12840 -7660
rect 12660 -7740 12840 -7720
rect 12660 -7800 12680 -7740
rect 12740 -7800 12760 -7740
rect 12820 -7800 12840 -7740
rect 12660 -7820 12840 -7800
rect 12660 -7880 12680 -7820
rect 12740 -7880 12760 -7820
rect 12820 -7880 12840 -7820
rect 12660 -7900 12840 -7880
rect 13900 -7500 14080 -7460
rect 13900 -7560 13920 -7500
rect 13980 -7560 14000 -7500
rect 14060 -7560 14080 -7500
rect 13900 -7580 14080 -7560
rect 13900 -7640 13920 -7580
rect 13980 -7640 14000 -7580
rect 14060 -7640 14080 -7580
rect 13900 -7660 14080 -7640
rect 13900 -7720 13920 -7660
rect 13980 -7720 14000 -7660
rect 14060 -7720 14080 -7660
rect 13900 -7740 14080 -7720
rect 13900 -7800 13920 -7740
rect 13980 -7800 14000 -7740
rect 14060 -7800 14080 -7740
rect 13900 -7820 14080 -7800
rect 13900 -7880 13920 -7820
rect 13980 -7880 14000 -7820
rect 14060 -7880 14080 -7820
rect 13900 -7900 14080 -7880
rect 15120 -7500 15300 -7460
rect 15120 -7560 15140 -7500
rect 15200 -7560 15220 -7500
rect 15280 -7560 15300 -7500
rect 15120 -7580 15300 -7560
rect 15120 -7640 15140 -7580
rect 15200 -7640 15220 -7580
rect 15280 -7640 15300 -7580
rect 15120 -7660 15300 -7640
rect 15120 -7720 15140 -7660
rect 15200 -7720 15220 -7660
rect 15280 -7720 15300 -7660
rect 15120 -7740 15300 -7720
rect 15120 -7800 15140 -7740
rect 15200 -7800 15220 -7740
rect 15280 -7800 15300 -7740
rect 15120 -7820 15300 -7800
rect 15120 -7880 15140 -7820
rect 15200 -7880 15220 -7820
rect 15280 -7880 15300 -7820
rect 15120 -7900 15300 -7880
rect 15720 -7480 15880 -7460
rect 15780 -7540 15820 -7480
rect 15720 -7560 15880 -7540
rect 15780 -7620 15820 -7560
rect 15720 -7740 15880 -7620
rect 17640 -7480 18820 -7300
rect 17640 -7540 17660 -7480
rect 17720 -7540 17740 -7480
rect 17840 -7540 17860 -7480
rect 17920 -7540 17940 -7480
rect 18000 -7540 18020 -7480
rect 18080 -7540 18100 -7480
rect 18160 -7540 18180 -7480
rect 18240 -7540 18260 -7480
rect 18320 -7540 18340 -7480
rect 18400 -7540 18420 -7480
rect 18480 -7540 18500 -7480
rect 18560 -7540 18580 -7480
rect 18640 -7540 18660 -7480
rect 18720 -7540 18740 -7480
rect 18800 -7540 18820 -7480
rect 17640 -7580 18820 -7540
rect 17640 -7640 17660 -7580
rect 17720 -7640 17740 -7580
rect 17840 -7640 17860 -7580
rect 17920 -7640 17940 -7580
rect 18000 -7640 18020 -7580
rect 18080 -7640 18100 -7580
rect 18160 -7640 18180 -7580
rect 18240 -7640 18260 -7580
rect 18320 -7640 18340 -7580
rect 18400 -7640 18420 -7580
rect 18480 -7640 18500 -7580
rect 18560 -7640 18580 -7580
rect 18640 -7640 18660 -7580
rect 18720 -7640 18740 -7580
rect 18800 -7640 18820 -7580
rect 17640 -7660 18820 -7640
rect 15780 -7800 15820 -7740
rect 15720 -7820 15880 -7800
rect 15780 -7880 15820 -7820
rect 15720 -7900 15880 -7880
rect 10880 -8100 11040 -8080
rect 10940 -8160 10980 -8100
rect 10880 -8180 11040 -8160
rect 10940 -8240 10980 -8180
rect 10880 -8320 11040 -8240
rect 10940 -8380 10980 -8320
rect 10880 -8400 11040 -8380
rect 10940 -8460 10980 -8400
rect 10880 -8480 11040 -8460
rect 12060 -8100 12220 -8080
rect 12120 -8160 12160 -8100
rect 12060 -8180 12220 -8160
rect 12120 -8240 12160 -8180
rect 12060 -8320 12220 -8240
rect 12120 -8380 12160 -8320
rect 12060 -8400 12220 -8380
rect 12120 -8460 12160 -8400
rect 12060 -8480 12220 -8460
rect 13300 -8100 13460 -8080
rect 13360 -8160 13400 -8100
rect 13300 -8180 13460 -8160
rect 13360 -8240 13400 -8180
rect 13300 -8320 13460 -8240
rect 13360 -8380 13400 -8320
rect 13300 -8400 13460 -8380
rect 13360 -8460 13400 -8400
rect 13300 -8480 13460 -8460
rect 14520 -8100 14680 -8080
rect 14580 -8160 14620 -8100
rect 14520 -8180 14680 -8160
rect 14580 -8240 14620 -8180
rect 14520 -8320 14680 -8240
rect 14580 -8380 14620 -8320
rect 14520 -8400 14680 -8380
rect 14580 -8460 14620 -8400
rect 14520 -8480 14680 -8460
rect 15720 -8100 15880 -8080
rect 15780 -8160 15820 -8100
rect 15720 -8180 15880 -8160
rect 15780 -8240 15820 -8180
rect 15720 -8320 15880 -8240
rect 15780 -8380 15820 -8320
rect 15720 -8400 15880 -8380
rect 15780 -8460 15820 -8400
rect 15720 -8480 15880 -8460
rect 10140 -9220 16620 -9160
rect 10140 -9300 10160 -9220
rect 10240 -9300 10280 -9220
rect 10360 -9300 10400 -9220
rect 10480 -9300 10520 -9220
rect 10600 -9300 10640 -9220
rect 10720 -9300 10760 -9220
rect 10840 -9300 10880 -9220
rect 10960 -9300 11000 -9220
rect 11080 -9300 11120 -9220
rect 11200 -9300 11240 -9220
rect 11320 -9300 11360 -9220
rect 11440 -9300 11480 -9220
rect 11560 -9300 11600 -9220
rect 11680 -9300 11720 -9220
rect 11800 -9300 11840 -9220
rect 11920 -9300 11960 -9220
rect 12040 -9300 12080 -9220
rect 12160 -9300 12200 -9220
rect 12280 -9300 12320 -9220
rect 12400 -9300 12440 -9220
rect 12520 -9300 12560 -9220
rect 12640 -9300 12680 -9220
rect 12760 -9300 12800 -9220
rect 12880 -9300 12920 -9220
rect 13000 -9300 13040 -9220
rect 13120 -9300 13160 -9220
rect 13240 -9300 13280 -9220
rect 13360 -9300 13400 -9220
rect 13480 -9300 13520 -9220
rect 13600 -9300 13640 -9220
rect 13720 -9300 13760 -9220
rect 13840 -9300 13880 -9220
rect 13960 -9300 14000 -9220
rect 14080 -9300 14120 -9220
rect 14200 -9300 14240 -9220
rect 14320 -9300 14360 -9220
rect 14440 -9300 14480 -9220
rect 14560 -9300 14600 -9220
rect 14680 -9300 14720 -9220
rect 14800 -9300 14840 -9220
rect 14920 -9300 14960 -9220
rect 15040 -9300 15080 -9220
rect 15160 -9300 15200 -9220
rect 15280 -9300 15320 -9220
rect 15400 -9300 15440 -9220
rect 15520 -9300 15560 -9220
rect 15640 -9300 15680 -9220
rect 15760 -9300 15800 -9220
rect 15880 -9300 15920 -9220
rect 16000 -9300 16040 -9220
rect 16120 -9300 16160 -9220
rect 16240 -9300 16280 -9220
rect 16360 -9300 16400 -9220
rect 16480 -9300 16520 -9220
rect 16600 -9300 16620 -9220
rect 10140 -9340 16620 -9300
rect 10140 -9420 10160 -9340
rect 10240 -9420 10280 -9340
rect 10360 -9420 10400 -9340
rect 10480 -9420 10520 -9340
rect 10600 -9420 10640 -9340
rect 10720 -9420 10760 -9340
rect 10840 -9420 10880 -9340
rect 10960 -9420 11000 -9340
rect 11080 -9420 11120 -9340
rect 11200 -9420 11240 -9340
rect 11320 -9420 11360 -9340
rect 11440 -9420 11480 -9340
rect 11560 -9420 11600 -9340
rect 11680 -9420 11720 -9340
rect 11800 -9420 11840 -9340
rect 11920 -9420 11960 -9340
rect 12040 -9420 12080 -9340
rect 12160 -9420 12200 -9340
rect 12280 -9420 12320 -9340
rect 12400 -9420 12440 -9340
rect 12520 -9420 12560 -9340
rect 12640 -9420 12680 -9340
rect 12760 -9420 12800 -9340
rect 12880 -9420 12920 -9340
rect 13000 -9420 13040 -9340
rect 13120 -9420 13160 -9340
rect 13240 -9420 13280 -9340
rect 13360 -9420 13400 -9340
rect 13480 -9420 13520 -9340
rect 13600 -9420 13640 -9340
rect 13720 -9420 13760 -9340
rect 13840 -9420 13880 -9340
rect 13960 -9420 14000 -9340
rect 14080 -9420 14120 -9340
rect 14200 -9420 14240 -9340
rect 14320 -9420 14360 -9340
rect 14440 -9420 14480 -9340
rect 14560 -9420 14600 -9340
rect 14680 -9420 14720 -9340
rect 14800 -9420 14840 -9340
rect 14920 -9420 14960 -9340
rect 15040 -9420 15080 -9340
rect 15160 -9420 15200 -9340
rect 15280 -9420 15320 -9340
rect 15400 -9420 15440 -9340
rect 15520 -9420 15560 -9340
rect 15640 -9420 15680 -9340
rect 15760 -9420 15800 -9340
rect 15880 -9420 15920 -9340
rect 16000 -9420 16040 -9340
rect 16120 -9420 16160 -9340
rect 16240 -9420 16280 -9340
rect 16360 -9420 16400 -9340
rect 16480 -9420 16520 -9340
rect 16600 -9420 16620 -9340
rect 10140 -9460 16620 -9420
rect 10140 -9540 10160 -9460
rect 10240 -9540 10280 -9460
rect 10360 -9540 10400 -9460
rect 10480 -9540 10520 -9460
rect 10600 -9540 10640 -9460
rect 10720 -9540 10760 -9460
rect 10840 -9540 10880 -9460
rect 10960 -9540 11000 -9460
rect 11080 -9540 11120 -9460
rect 11200 -9540 11240 -9460
rect 11320 -9540 11360 -9460
rect 11440 -9540 11480 -9460
rect 11560 -9540 11600 -9460
rect 11680 -9540 11720 -9460
rect 11800 -9540 11840 -9460
rect 11920 -9540 11960 -9460
rect 12040 -9540 12080 -9460
rect 12160 -9540 12200 -9460
rect 12280 -9540 12320 -9460
rect 12400 -9540 12440 -9460
rect 12520 -9540 12560 -9460
rect 12640 -9540 12680 -9460
rect 12760 -9540 12800 -9460
rect 12880 -9540 12920 -9460
rect 13000 -9540 13040 -9460
rect 13120 -9540 13160 -9460
rect 13240 -9540 13280 -9460
rect 13360 -9540 13400 -9460
rect 13480 -9540 13520 -9460
rect 13600 -9540 13640 -9460
rect 13720 -9540 13760 -9460
rect 13840 -9540 13880 -9460
rect 13960 -9540 14000 -9460
rect 14080 -9540 14120 -9460
rect 14200 -9540 14240 -9460
rect 14320 -9540 14360 -9460
rect 14440 -9540 14480 -9460
rect 14560 -9540 14600 -9460
rect 14680 -9540 14720 -9460
rect 14800 -9540 14840 -9460
rect 14920 -9540 14960 -9460
rect 15040 -9540 15080 -9460
rect 15160 -9540 15200 -9460
rect 15280 -9540 15320 -9460
rect 15400 -9540 15440 -9460
rect 15520 -9540 15560 -9460
rect 15640 -9540 15680 -9460
rect 15760 -9540 15800 -9460
rect 15880 -9540 15920 -9460
rect 16000 -9540 16040 -9460
rect 16120 -9540 16160 -9460
rect 16240 -9540 16280 -9460
rect 16360 -9540 16400 -9460
rect 16480 -9540 16520 -9460
rect 16600 -9540 16620 -9460
rect 10140 -9580 16620 -9540
rect 10140 -9660 10160 -9580
rect 10240 -9660 10280 -9580
rect 10360 -9660 10400 -9580
rect 10480 -9660 10520 -9580
rect 10600 -9660 10640 -9580
rect 10720 -9660 10760 -9580
rect 10840 -9660 10880 -9580
rect 10960 -9660 11000 -9580
rect 11080 -9660 11120 -9580
rect 11200 -9660 11240 -9580
rect 11320 -9660 11360 -9580
rect 11440 -9660 11480 -9580
rect 11560 -9660 11600 -9580
rect 11680 -9660 11720 -9580
rect 11800 -9660 11840 -9580
rect 11920 -9660 11960 -9580
rect 12040 -9660 12080 -9580
rect 12160 -9660 12200 -9580
rect 12280 -9660 12320 -9580
rect 12400 -9660 12440 -9580
rect 12520 -9660 12560 -9580
rect 12640 -9660 12680 -9580
rect 12760 -9660 12800 -9580
rect 12880 -9660 12920 -9580
rect 13000 -9660 13040 -9580
rect 13120 -9660 13160 -9580
rect 13240 -9660 13280 -9580
rect 13360 -9660 13400 -9580
rect 13480 -9660 13520 -9580
rect 13600 -9660 13640 -9580
rect 13720 -9660 13760 -9580
rect 13840 -9660 13880 -9580
rect 13960 -9660 14000 -9580
rect 14080 -9660 14120 -9580
rect 14200 -9660 14240 -9580
rect 14320 -9660 14360 -9580
rect 14440 -9660 14480 -9580
rect 14560 -9660 14600 -9580
rect 14680 -9660 14720 -9580
rect 14800 -9660 14840 -9580
rect 14920 -9660 14960 -9580
rect 15040 -9660 15080 -9580
rect 15160 -9660 15200 -9580
rect 15280 -9660 15320 -9580
rect 15400 -9660 15440 -9580
rect 15520 -9660 15560 -9580
rect 15640 -9660 15680 -9580
rect 15760 -9660 15800 -9580
rect 15880 -9660 15920 -9580
rect 16000 -9660 16040 -9580
rect 16120 -9660 16160 -9580
rect 16240 -9660 16280 -9580
rect 16360 -9660 16400 -9580
rect 16480 -9660 16520 -9580
rect 16600 -9660 16620 -9580
rect 10140 -9700 16620 -9660
rect 10140 -9780 10160 -9700
rect 10240 -9780 10280 -9700
rect 10360 -9780 10400 -9700
rect 10480 -9780 10520 -9700
rect 10600 -9780 10640 -9700
rect 10720 -9780 10760 -9700
rect 10840 -9780 10880 -9700
rect 10960 -9780 11000 -9700
rect 11080 -9780 11120 -9700
rect 11200 -9780 11240 -9700
rect 11320 -9780 11360 -9700
rect 11440 -9780 11480 -9700
rect 11560 -9780 11600 -9700
rect 11680 -9780 11720 -9700
rect 11800 -9780 11840 -9700
rect 11920 -9780 11960 -9700
rect 12040 -9780 12080 -9700
rect 12160 -9780 12200 -9700
rect 12280 -9780 12320 -9700
rect 12400 -9780 12440 -9700
rect 12520 -9780 12560 -9700
rect 12640 -9780 12680 -9700
rect 12760 -9780 12800 -9700
rect 12880 -9780 12920 -9700
rect 13000 -9780 13040 -9700
rect 13120 -9780 13160 -9700
rect 13240 -9780 13280 -9700
rect 13360 -9780 13400 -9700
rect 13480 -9780 13520 -9700
rect 13600 -9780 13640 -9700
rect 13720 -9780 13760 -9700
rect 13840 -9780 13880 -9700
rect 13960 -9780 14000 -9700
rect 14080 -9780 14120 -9700
rect 14200 -9780 14240 -9700
rect 14320 -9780 14360 -9700
rect 14440 -9780 14480 -9700
rect 14560 -9780 14600 -9700
rect 14680 -9780 14720 -9700
rect 14800 -9780 14840 -9700
rect 14920 -9780 14960 -9700
rect 15040 -9780 15080 -9700
rect 15160 -9780 15200 -9700
rect 15280 -9780 15320 -9700
rect 15400 -9780 15440 -9700
rect 15520 -9780 15560 -9700
rect 15640 -9780 15680 -9700
rect 15760 -9780 15800 -9700
rect 15880 -9780 15920 -9700
rect 16000 -9780 16040 -9700
rect 16120 -9780 16160 -9700
rect 16240 -9780 16280 -9700
rect 16360 -9780 16400 -9700
rect 16480 -9780 16520 -9700
rect 16600 -9780 16620 -9700
rect 10140 -9820 16620 -9780
rect 10140 -9900 10160 -9820
rect 10240 -9900 10280 -9820
rect 10360 -9900 10400 -9820
rect 10480 -9900 10520 -9820
rect 10600 -9900 10640 -9820
rect 10720 -9900 10760 -9820
rect 10840 -9900 10880 -9820
rect 10960 -9900 11000 -9820
rect 11080 -9900 11120 -9820
rect 11200 -9900 11240 -9820
rect 11320 -9900 11360 -9820
rect 11440 -9900 11480 -9820
rect 11560 -9900 11600 -9820
rect 11680 -9900 11720 -9820
rect 11800 -9900 11840 -9820
rect 11920 -9900 11960 -9820
rect 12040 -9900 12080 -9820
rect 12160 -9900 12200 -9820
rect 12280 -9900 12320 -9820
rect 12400 -9900 12440 -9820
rect 12520 -9900 12560 -9820
rect 12640 -9900 12680 -9820
rect 12760 -9900 12800 -9820
rect 12880 -9900 12920 -9820
rect 13000 -9900 13040 -9820
rect 13120 -9900 13160 -9820
rect 13240 -9900 13280 -9820
rect 13360 -9900 13400 -9820
rect 13480 -9900 13520 -9820
rect 13600 -9900 13640 -9820
rect 13720 -9900 13760 -9820
rect 13840 -9900 13880 -9820
rect 13960 -9900 14000 -9820
rect 14080 -9900 14120 -9820
rect 14200 -9900 14240 -9820
rect 14320 -9900 14360 -9820
rect 14440 -9900 14480 -9820
rect 14560 -9900 14600 -9820
rect 14680 -9900 14720 -9820
rect 14800 -9900 14840 -9820
rect 14920 -9900 14960 -9820
rect 15040 -9900 15080 -9820
rect 15160 -9900 15200 -9820
rect 15280 -9900 15320 -9820
rect 15400 -9900 15440 -9820
rect 15520 -9900 15560 -9820
rect 15640 -9900 15680 -9820
rect 15760 -9900 15800 -9820
rect 15880 -9900 15920 -9820
rect 16000 -9900 16040 -9820
rect 16120 -9900 16160 -9820
rect 16240 -9900 16280 -9820
rect 16360 -9900 16400 -9820
rect 16480 -9900 16520 -9820
rect 16600 -9900 16620 -9820
rect 10140 -9940 16620 -9900
rect 9300 -10020 9700 -10000
rect 9300 -10100 9320 -10020
rect 9400 -10100 9460 -10020
rect 9540 -10100 9600 -10020
rect 9680 -10100 9700 -10020
rect 9300 -10160 9700 -10100
rect 10140 -10020 10160 -9940
rect 10240 -10020 10280 -9940
rect 10360 -10020 10400 -9940
rect 10480 -10020 10520 -9940
rect 10600 -10020 10640 -9940
rect 10720 -10020 10760 -9940
rect 10840 -10020 10880 -9940
rect 10960 -10020 11000 -9940
rect 11080 -10020 11120 -9940
rect 11200 -10020 11240 -9940
rect 11320 -10020 11360 -9940
rect 11440 -10020 11480 -9940
rect 11560 -10020 11600 -9940
rect 11680 -10020 11720 -9940
rect 11800 -10020 11840 -9940
rect 11920 -10020 11960 -9940
rect 12040 -10020 12080 -9940
rect 12160 -10020 12200 -9940
rect 12280 -10020 12320 -9940
rect 12400 -10020 12440 -9940
rect 12520 -10020 12560 -9940
rect 12640 -10020 12680 -9940
rect 12760 -10020 12800 -9940
rect 12880 -10020 12920 -9940
rect 13000 -10020 13040 -9940
rect 13120 -10020 13160 -9940
rect 13240 -10020 13280 -9940
rect 13360 -10020 13400 -9940
rect 13480 -10020 13520 -9940
rect 13600 -10020 13640 -9940
rect 13720 -10020 13760 -9940
rect 13840 -10020 13880 -9940
rect 13960 -10020 14000 -9940
rect 14080 -10020 14120 -9940
rect 14200 -10020 14240 -9940
rect 14320 -10020 14360 -9940
rect 14440 -10020 14480 -9940
rect 14560 -10020 14600 -9940
rect 14680 -10020 14720 -9940
rect 14800 -10020 14840 -9940
rect 14920 -10020 14960 -9940
rect 15040 -10020 15080 -9940
rect 15160 -10020 15200 -9940
rect 15280 -10020 15320 -9940
rect 15400 -10020 15440 -9940
rect 15520 -10020 15560 -9940
rect 15640 -10020 15680 -9940
rect 15760 -10020 15800 -9940
rect 15880 -10020 15920 -9940
rect 16000 -10020 16040 -9940
rect 16120 -10020 16160 -9940
rect 16240 -10020 16280 -9940
rect 16360 -10020 16400 -9940
rect 16480 -10020 16520 -9940
rect 16600 -10020 16620 -9940
rect 10140 -10060 16620 -10020
rect 10140 -10140 10160 -10060
rect 10240 -10140 10280 -10060
rect 10360 -10140 10400 -10060
rect 10480 -10140 10520 -10060
rect 10600 -10140 10640 -10060
rect 10720 -10140 10760 -10060
rect 10840 -10140 10880 -10060
rect 10960 -10140 11000 -10060
rect 11080 -10140 11120 -10060
rect 11200 -10140 11240 -10060
rect 11320 -10140 11360 -10060
rect 11440 -10140 11480 -10060
rect 11560 -10140 11600 -10060
rect 11680 -10140 11720 -10060
rect 11800 -10140 11840 -10060
rect 11920 -10140 11960 -10060
rect 12040 -10140 12080 -10060
rect 12160 -10140 12200 -10060
rect 12280 -10140 12320 -10060
rect 12400 -10140 12440 -10060
rect 12520 -10140 12560 -10060
rect 12640 -10140 12680 -10060
rect 12760 -10140 12800 -10060
rect 12880 -10140 12920 -10060
rect 13000 -10140 13040 -10060
rect 13120 -10140 13160 -10060
rect 13240 -10140 13280 -10060
rect 13360 -10140 13400 -10060
rect 13480 -10140 13520 -10060
rect 13600 -10140 13640 -10060
rect 13720 -10140 13760 -10060
rect 13840 -10140 13880 -10060
rect 13960 -10140 14000 -10060
rect 14080 -10140 14120 -10060
rect 14200 -10140 14240 -10060
rect 14320 -10140 14360 -10060
rect 14440 -10140 14480 -10060
rect 14560 -10140 14600 -10060
rect 14680 -10140 14720 -10060
rect 14800 -10140 14840 -10060
rect 14920 -10140 14960 -10060
rect 15040 -10140 15080 -10060
rect 15160 -10140 15200 -10060
rect 15280 -10140 15320 -10060
rect 15400 -10140 15440 -10060
rect 15520 -10140 15560 -10060
rect 15640 -10140 15680 -10060
rect 15760 -10140 15800 -10060
rect 15880 -10140 15920 -10060
rect 16000 -10140 16040 -10060
rect 16120 -10140 16160 -10060
rect 16240 -10140 16280 -10060
rect 16360 -10140 16400 -10060
rect 16480 -10140 16520 -10060
rect 16600 -10140 16620 -10060
rect 10140 -10160 16620 -10140
rect 17100 -10020 17500 -10000
rect 17100 -10100 17120 -10020
rect 17200 -10100 17260 -10020
rect 17340 -10100 17400 -10020
rect 17480 -10100 17500 -10020
rect 17100 -10160 17500 -10100
rect 9300 -10240 9320 -10160
rect 9400 -10240 9460 -10160
rect 9540 -10240 9600 -10160
rect 9680 -10240 9700 -10160
rect 9300 -10300 9700 -10240
rect 9300 -10380 9320 -10300
rect 9400 -10380 9460 -10300
rect 9540 -10380 9600 -10300
rect 9680 -10380 9700 -10300
rect 9300 -10400 9700 -10380
rect 17100 -10240 17120 -10160
rect 17200 -10240 17260 -10160
rect 17340 -10240 17400 -10160
rect 17480 -10240 17500 -10160
rect 17100 -10300 17500 -10240
rect 17100 -10380 17120 -10300
rect 17200 -10380 17260 -10300
rect 17340 -10380 17400 -10300
rect 17480 -10380 17500 -10300
rect 17100 -10400 17500 -10380
rect 13200 -10620 13600 -10600
rect 13200 -10680 13220 -10620
rect 13280 -10680 13320 -10620
rect 13380 -10680 13420 -10620
rect 13480 -10680 13520 -10620
rect 13580 -10680 13600 -10620
rect 13200 -10720 13600 -10680
rect 13200 -10780 13220 -10720
rect 13280 -10780 13320 -10720
rect 13380 -10780 13420 -10720
rect 13480 -10780 13520 -10720
rect 13580 -10780 13600 -10720
rect 13200 -10820 13600 -10780
rect 13200 -10880 13220 -10820
rect 13280 -10880 13320 -10820
rect 13380 -10880 13420 -10820
rect 13480 -10880 13520 -10820
rect 13580 -10880 13600 -10820
rect 13200 -10920 13600 -10880
rect 13200 -10980 13220 -10920
rect 13280 -10980 13320 -10920
rect 13380 -10980 13420 -10920
rect 13480 -10980 13520 -10920
rect 13580 -10980 13600 -10920
rect 13200 -11000 13600 -10980
rect 8240 -11420 8640 -11400
rect 8240 -11480 8260 -11420
rect 8320 -11480 8360 -11420
rect 8420 -11480 8460 -11420
rect 8520 -11480 8560 -11420
rect 8620 -11480 8640 -11420
rect 8240 -11500 8640 -11480
rect 8240 -11560 8260 -11500
rect 8320 -11560 8360 -11500
rect 8420 -11560 8460 -11500
rect 8520 -11560 8560 -11500
rect 8620 -11560 8640 -11500
rect 8240 -11600 8640 -11560
rect 8240 -11660 8260 -11600
rect 8320 -11660 8360 -11600
rect 8420 -11660 8460 -11600
rect 8520 -11660 8560 -11600
rect 8620 -11660 8640 -11600
rect 8240 -11700 8640 -11660
rect 8240 -11760 8260 -11700
rect 8320 -11760 8360 -11700
rect 8420 -11760 8460 -11700
rect 8520 -11760 8560 -11700
rect 8620 -11760 8640 -11700
rect 8240 -11780 8640 -11760
rect 18160 -11420 18560 -11400
rect 18160 -11480 18180 -11420
rect 18240 -11480 18280 -11420
rect 18340 -11480 18380 -11420
rect 18440 -11480 18480 -11420
rect 18540 -11480 18560 -11420
rect 18160 -11500 18560 -11480
rect 18160 -11560 18180 -11500
rect 18240 -11560 18280 -11500
rect 18340 -11560 18380 -11500
rect 18440 -11560 18480 -11500
rect 18540 -11560 18560 -11500
rect 18160 -11600 18560 -11560
rect 18160 -11660 18180 -11600
rect 18240 -11660 18280 -11600
rect 18340 -11660 18380 -11600
rect 18440 -11660 18480 -11600
rect 18540 -11660 18560 -11600
rect 18160 -11700 18560 -11660
rect 18160 -11760 18180 -11700
rect 18240 -11760 18280 -11700
rect 18340 -11760 18380 -11700
rect 18440 -11760 18480 -11700
rect 18540 -11760 18560 -11700
rect 18160 -11780 18560 -11760
<< via1 >>
rect 11400 -2040 11460 -1980
rect 11500 -2040 11560 -1980
rect 11400 -2120 11460 -2060
rect 11500 -2120 11560 -2060
rect 11400 -2240 11460 -2180
rect 11500 -2240 11560 -2180
rect 11400 -2320 11460 -2260
rect 11500 -2320 11560 -2260
rect 12640 -2040 12700 -1980
rect 12740 -2040 12800 -1980
rect 12640 -2120 12700 -2060
rect 12740 -2120 12800 -2060
rect 12640 -2240 12700 -2180
rect 12740 -2240 12800 -2180
rect 12640 -2320 12700 -2260
rect 12740 -2320 12800 -2260
rect 13860 -2040 13920 -1980
rect 13960 -2040 14020 -1980
rect 13860 -2120 13920 -2060
rect 13960 -2120 14020 -2060
rect 13860 -2240 13920 -2180
rect 13960 -2240 14020 -2180
rect 13860 -2320 13920 -2260
rect 13960 -2320 14020 -2260
rect 15100 -2040 15160 -1980
rect 15200 -2040 15260 -1980
rect 15100 -2120 15160 -2060
rect 15200 -2120 15260 -2060
rect 15100 -2240 15160 -2180
rect 15200 -2240 15260 -2180
rect 15100 -2320 15160 -2260
rect 15200 -2320 15260 -2260
rect 7400 -2940 7460 -2880
rect 7400 -3120 7460 -3060
rect 8000 -2940 8060 -2880
rect 8000 -3120 8060 -3060
rect 8640 -2940 8700 -2880
rect 8640 -3120 8700 -3060
rect 9240 -2940 9300 -2880
rect 9240 -3120 9300 -3060
rect 9880 -2940 9940 -2880
rect 9880 -3120 9940 -3060
rect 11140 -3020 11220 -2940
rect 11260 -3020 11340 -2940
rect 11380 -3020 11460 -2940
rect 11500 -3020 11580 -2940
rect 11620 -3020 11700 -2940
rect 11740 -3020 11820 -2940
rect 11860 -3020 11940 -2940
rect 11980 -3020 12060 -2940
rect 12100 -3020 12180 -2940
rect 12220 -3020 12300 -2940
rect 12340 -3020 12420 -2940
rect 12460 -3020 12540 -2940
rect 12580 -3020 12660 -2940
rect 12700 -3020 12780 -2940
rect 12820 -3020 12900 -2940
rect 12940 -3020 13020 -2940
rect 13060 -3020 13140 -2940
rect 13180 -3020 13260 -2940
rect 13300 -3020 13380 -2940
rect 13420 -3020 13500 -2940
rect 13540 -3020 13620 -2940
rect 13660 -3020 13740 -2940
rect 13780 -3020 13860 -2940
rect 13900 -3020 13980 -2940
rect 14020 -3020 14100 -2940
rect 14140 -3020 14220 -2940
rect 14260 -3020 14340 -2940
rect 14380 -3020 14460 -2940
rect 14500 -3020 14580 -2940
rect 14620 -3020 14700 -2940
rect 14740 -3020 14820 -2940
rect 14860 -3020 14940 -2940
rect 14980 -3020 15060 -2940
rect 15100 -3020 15180 -2940
rect 15220 -3020 15300 -2940
rect 15340 -3020 15420 -2940
rect 15460 -3020 15540 -2940
rect 15580 -3020 15660 -2940
rect 11140 -3160 11220 -3080
rect 11260 -3160 11340 -3080
rect 11380 -3160 11460 -3080
rect 11500 -3160 11580 -3080
rect 11620 -3160 11700 -3080
rect 11740 -3160 11820 -3080
rect 11860 -3160 11940 -3080
rect 11980 -3160 12060 -3080
rect 12100 -3160 12180 -3080
rect 12220 -3160 12300 -3080
rect 12340 -3160 12420 -3080
rect 12460 -3160 12540 -3080
rect 12580 -3160 12660 -3080
rect 12700 -3160 12780 -3080
rect 12820 -3160 12900 -3080
rect 12940 -3160 13020 -3080
rect 13060 -3160 13140 -3080
rect 13180 -3160 13260 -3080
rect 13300 -3160 13380 -3080
rect 13420 -3160 13500 -3080
rect 13540 -3160 13620 -3080
rect 13660 -3160 13740 -3080
rect 13780 -3160 13860 -3080
rect 13900 -3160 13980 -3080
rect 14020 -3160 14100 -3080
rect 14140 -3160 14220 -3080
rect 14260 -3160 14340 -3080
rect 14380 -3160 14460 -3080
rect 14500 -3160 14580 -3080
rect 14620 -3160 14700 -3080
rect 14740 -3160 14820 -3080
rect 14860 -3160 14940 -3080
rect 14980 -3160 15060 -3080
rect 15100 -3160 15180 -3080
rect 15220 -3160 15300 -3080
rect 15340 -3160 15420 -3080
rect 15460 -3160 15540 -3080
rect 15580 -3160 15660 -3080
rect 16840 -2940 16900 -2880
rect 16840 -3120 16900 -3060
rect 17440 -2940 17500 -2880
rect 17440 -3120 17500 -3060
rect 18080 -2940 18140 -2880
rect 18080 -3120 18140 -3060
rect 18680 -2940 18740 -2880
rect 18680 -3120 18740 -3060
rect 19300 -2940 19360 -2880
rect 19300 -3120 19360 -3060
rect 11140 -3300 11220 -3220
rect 11260 -3300 11340 -3220
rect 11380 -3300 11460 -3220
rect 11500 -3300 11580 -3220
rect 11620 -3300 11700 -3220
rect 11740 -3300 11820 -3220
rect 11860 -3300 11940 -3220
rect 11980 -3300 12060 -3220
rect 12100 -3300 12180 -3220
rect 12220 -3300 12300 -3220
rect 12340 -3300 12420 -3220
rect 12460 -3300 12540 -3220
rect 12580 -3300 12660 -3220
rect 12700 -3300 12780 -3220
rect 12820 -3300 12900 -3220
rect 12940 -3300 13020 -3220
rect 13060 -3300 13140 -3220
rect 13180 -3300 13260 -3220
rect 13300 -3300 13380 -3220
rect 13420 -3300 13500 -3220
rect 13540 -3300 13620 -3220
rect 13660 -3300 13740 -3220
rect 13780 -3300 13860 -3220
rect 13900 -3300 13980 -3220
rect 14020 -3300 14100 -3220
rect 14140 -3300 14220 -3220
rect 14260 -3300 14340 -3220
rect 14380 -3300 14460 -3220
rect 14500 -3300 14580 -3220
rect 14620 -3300 14700 -3220
rect 14740 -3300 14820 -3220
rect 14860 -3300 14940 -3220
rect 14980 -3300 15060 -3220
rect 15100 -3300 15180 -3220
rect 15220 -3300 15300 -3220
rect 15340 -3300 15420 -3220
rect 15460 -3300 15540 -3220
rect 15580 -3300 15660 -3220
rect 7480 -3500 7560 -3420
rect 7580 -3500 7660 -3420
rect 7680 -3500 7760 -3420
rect 7780 -3500 7860 -3420
rect 7880 -3500 7960 -3420
rect 7980 -3500 8060 -3420
rect 8080 -3500 8160 -3420
rect 8180 -3500 8260 -3420
rect 8280 -3500 8360 -3420
rect 8380 -3500 8460 -3420
rect 8480 -3500 8560 -3420
rect 8580 -3500 8660 -3420
rect 8680 -3500 8760 -3420
rect 8780 -3500 8860 -3420
rect 8880 -3500 8960 -3420
rect 8980 -3500 9060 -3420
rect 9080 -3500 9160 -3420
rect 9180 -3500 9260 -3420
rect 9280 -3500 9360 -3420
rect 9380 -3500 9460 -3420
rect 9480 -3500 9560 -3420
rect 9580 -3500 9660 -3420
rect 9680 -3500 9760 -3420
rect 9780 -3500 9860 -3420
rect 7480 -3640 7560 -3560
rect 7580 -3640 7660 -3560
rect 7680 -3640 7760 -3560
rect 7780 -3640 7860 -3560
rect 7880 -3640 7960 -3560
rect 7980 -3640 8060 -3560
rect 8080 -3640 8160 -3560
rect 8180 -3640 8260 -3560
rect 8280 -3640 8360 -3560
rect 8380 -3640 8460 -3560
rect 8480 -3640 8560 -3560
rect 8580 -3640 8660 -3560
rect 8680 -3640 8760 -3560
rect 8780 -3640 8860 -3560
rect 8880 -3640 8960 -3560
rect 8980 -3640 9060 -3560
rect 9080 -3640 9160 -3560
rect 9180 -3640 9260 -3560
rect 9280 -3640 9360 -3560
rect 9380 -3640 9460 -3560
rect 9480 -3640 9560 -3560
rect 9580 -3640 9660 -3560
rect 9680 -3640 9760 -3560
rect 9780 -3640 9860 -3560
rect 7480 -3780 7560 -3700
rect 7580 -3780 7660 -3700
rect 7680 -3780 7760 -3700
rect 7780 -3780 7860 -3700
rect 7880 -3780 7960 -3700
rect 7980 -3780 8060 -3700
rect 8080 -3780 8160 -3700
rect 8180 -3780 8260 -3700
rect 8280 -3780 8360 -3700
rect 8380 -3780 8460 -3700
rect 8480 -3780 8560 -3700
rect 8580 -3780 8660 -3700
rect 8680 -3780 8760 -3700
rect 8780 -3780 8860 -3700
rect 8880 -3780 8960 -3700
rect 8980 -3780 9060 -3700
rect 9080 -3780 9160 -3700
rect 9180 -3780 9260 -3700
rect 9280 -3780 9360 -3700
rect 9380 -3780 9460 -3700
rect 9480 -3780 9560 -3700
rect 9580 -3780 9660 -3700
rect 9680 -3780 9760 -3700
rect 9780 -3780 9860 -3700
rect 16920 -3500 17000 -3420
rect 17020 -3500 17100 -3420
rect 17120 -3500 17200 -3420
rect 17220 -3500 17300 -3420
rect 17320 -3500 17400 -3420
rect 17420 -3500 17500 -3420
rect 17520 -3500 17600 -3420
rect 17620 -3500 17700 -3420
rect 17720 -3500 17800 -3420
rect 17820 -3500 17900 -3420
rect 17920 -3500 18000 -3420
rect 18020 -3500 18100 -3420
rect 18120 -3500 18200 -3420
rect 18220 -3500 18300 -3420
rect 18320 -3500 18400 -3420
rect 18420 -3500 18500 -3420
rect 18520 -3500 18600 -3420
rect 18620 -3500 18700 -3420
rect 18720 -3500 18800 -3420
rect 18820 -3500 18900 -3420
rect 18920 -3500 19000 -3420
rect 19020 -3500 19100 -3420
rect 19120 -3500 19200 -3420
rect 19220 -3500 19300 -3420
rect 16920 -3640 17000 -3560
rect 17020 -3640 17100 -3560
rect 17120 -3640 17200 -3560
rect 17220 -3640 17300 -3560
rect 17320 -3640 17400 -3560
rect 17420 -3640 17500 -3560
rect 17520 -3640 17600 -3560
rect 17620 -3640 17700 -3560
rect 17720 -3640 17800 -3560
rect 17820 -3640 17900 -3560
rect 17920 -3640 18000 -3560
rect 18020 -3640 18100 -3560
rect 18120 -3640 18200 -3560
rect 18220 -3640 18300 -3560
rect 18320 -3640 18400 -3560
rect 18420 -3640 18500 -3560
rect 18520 -3640 18600 -3560
rect 18620 -3640 18700 -3560
rect 18720 -3640 18800 -3560
rect 18820 -3640 18900 -3560
rect 18920 -3640 19000 -3560
rect 19020 -3640 19100 -3560
rect 19120 -3640 19200 -3560
rect 19220 -3640 19300 -3560
rect 16920 -3780 17000 -3700
rect 17020 -3780 17100 -3700
rect 17120 -3780 17200 -3700
rect 17220 -3780 17300 -3700
rect 17320 -3780 17400 -3700
rect 17420 -3780 17500 -3700
rect 17520 -3780 17600 -3700
rect 17620 -3780 17700 -3700
rect 17720 -3780 17800 -3700
rect 17820 -3780 17900 -3700
rect 17920 -3780 18000 -3700
rect 18020 -3780 18100 -3700
rect 18120 -3780 18200 -3700
rect 18220 -3780 18300 -3700
rect 18320 -3780 18400 -3700
rect 18420 -3780 18500 -3700
rect 18520 -3780 18600 -3700
rect 18620 -3780 18700 -3700
rect 18720 -3780 18800 -3700
rect 18820 -3780 18900 -3700
rect 18920 -3780 19000 -3700
rect 19020 -3780 19100 -3700
rect 19120 -3780 19200 -3700
rect 19220 -3780 19300 -3700
rect 8360 -4020 8420 -3960
rect 8360 -4200 8420 -4140
rect 8820 -4020 8880 -3960
rect 13220 -3980 13300 -3900
rect 13360 -3980 13440 -3900
rect 13500 -3980 13580 -3900
rect 8820 -4200 8880 -4140
rect 8620 -4500 8680 -4440
rect 8620 -4600 8680 -4540
rect 10300 -4500 10360 -4440
rect 10300 -4580 10360 -4520
rect 10300 -4660 10360 -4600
rect 10620 -4500 10680 -4440
rect 10620 -4580 10680 -4520
rect 10620 -4660 10680 -4600
rect 12100 -4500 12160 -4440
rect 12100 -4580 12160 -4520
rect 12100 -4660 12160 -4600
rect 13220 -4100 13300 -4020
rect 13360 -4100 13440 -4020
rect 13500 -4100 13580 -4020
rect 13220 -4220 13300 -4140
rect 13360 -4220 13440 -4140
rect 13500 -4220 13580 -4140
rect 13220 -4340 13300 -4260
rect 13360 -4340 13440 -4260
rect 13500 -4340 13580 -4260
rect 12420 -4500 12480 -4440
rect 12420 -4580 12480 -4520
rect 12420 -4660 12480 -4600
rect 13220 -4460 13300 -4380
rect 13360 -4460 13440 -4380
rect 13500 -4460 13580 -4380
rect 13220 -4580 13300 -4500
rect 13360 -4580 13440 -4500
rect 13500 -4580 13580 -4500
rect 13220 -4700 13300 -4620
rect 13360 -4700 13440 -4620
rect 13500 -4700 13580 -4620
rect 14300 -4500 14360 -4440
rect 14300 -4580 14360 -4520
rect 14300 -4660 14360 -4600
rect 13220 -4820 13300 -4740
rect 13360 -4820 13440 -4740
rect 13500 -4820 13580 -4740
rect 13220 -4940 13300 -4860
rect 13360 -4940 13440 -4860
rect 13500 -4940 13580 -4860
rect 13220 -5060 13300 -4980
rect 13360 -5060 13440 -4980
rect 13500 -5060 13580 -4980
rect 14620 -4500 14680 -4440
rect 14620 -4580 14680 -4520
rect 14620 -4660 14680 -4600
rect 16100 -4500 16160 -4440
rect 16100 -4580 16160 -4520
rect 16100 -4660 16160 -4600
rect 17960 -4020 18020 -3960
rect 17960 -4200 18020 -4140
rect 18420 -4020 18480 -3960
rect 18420 -4200 18480 -4140
rect 16420 -4500 16480 -4440
rect 16420 -4580 16480 -4520
rect 16420 -4660 16480 -4600
rect 18140 -4500 18200 -4440
rect 18140 -4600 18200 -4540
rect 10380 -5180 10440 -5120
rect 10540 -5180 10600 -5120
rect 12180 -5180 12240 -5120
rect 12340 -5180 12400 -5120
rect 13220 -5180 13300 -5100
rect 13360 -5180 13440 -5100
rect 13500 -5180 13580 -5100
rect 13220 -5300 13300 -5220
rect 13360 -5300 13440 -5220
rect 13500 -5300 13580 -5220
rect 14380 -5180 14440 -5120
rect 14540 -5180 14600 -5120
rect 16180 -5180 16240 -5120
rect 16340 -5180 16400 -5120
rect 13220 -5420 13300 -5340
rect 13360 -5420 13440 -5340
rect 13500 -5420 13580 -5340
rect 13220 -5540 13300 -5460
rect 13360 -5540 13440 -5460
rect 13500 -5540 13580 -5460
rect 10380 -5780 10440 -5720
rect 10540 -5780 10600 -5720
rect 12180 -5780 12240 -5720
rect 12340 -5780 12400 -5720
rect 13220 -5660 13300 -5580
rect 13360 -5660 13440 -5580
rect 13500 -5660 13580 -5580
rect 13220 -5780 13300 -5700
rect 13360 -5780 13440 -5700
rect 13500 -5780 13580 -5700
rect 7920 -6020 7980 -5960
rect 7920 -6200 7980 -6140
rect 8540 -6020 8600 -5960
rect 8540 -6200 8600 -6140
rect 9140 -6020 9200 -5960
rect 9140 -6200 9200 -6140
rect 10300 -6000 10360 -5940
rect 10300 -6080 10360 -6020
rect 10300 -6160 10360 -6100
rect 14380 -5780 14440 -5720
rect 14540 -5780 14600 -5720
rect 10620 -6000 10680 -5940
rect 10620 -6080 10680 -6020
rect 10620 -6160 10680 -6100
rect 12100 -6600 12160 -6540
rect 12100 -6680 12160 -6620
rect 12100 -6760 12160 -6700
rect 13220 -5900 13300 -5820
rect 13360 -5900 13440 -5820
rect 13500 -5900 13580 -5820
rect 16180 -5780 16240 -5720
rect 16340 -5780 16400 -5720
rect 13220 -6020 13300 -5940
rect 13360 -6020 13440 -5940
rect 13500 -6020 13580 -5940
rect 13220 -6140 13300 -6060
rect 13360 -6140 13440 -6060
rect 13500 -6140 13580 -6060
rect 13220 -6260 13300 -6180
rect 13360 -6260 13440 -6180
rect 13500 -6260 13580 -6180
rect 13220 -6380 13300 -6300
rect 13360 -6380 13440 -6300
rect 13500 -6380 13580 -6300
rect 13220 -6500 13300 -6420
rect 13360 -6500 13440 -6420
rect 13500 -6500 13580 -6420
rect 12420 -6600 12480 -6540
rect 12420 -6680 12480 -6620
rect 12420 -6760 12480 -6700
rect 13220 -6620 13300 -6540
rect 13360 -6620 13440 -6540
rect 13500 -6620 13580 -6540
rect 13220 -6740 13300 -6660
rect 13360 -6740 13440 -6660
rect 13500 -6740 13580 -6660
rect 14300 -6600 14360 -6540
rect 14300 -6680 14360 -6620
rect 14300 -6760 14360 -6700
rect 13220 -6860 13300 -6780
rect 13360 -6860 13440 -6780
rect 13500 -6860 13580 -6780
rect 13220 -6980 13300 -6900
rect 13360 -6980 13440 -6900
rect 13500 -6980 13580 -6900
rect 16100 -6000 16160 -5940
rect 16100 -6080 16160 -6020
rect 16100 -6160 16160 -6100
rect 14620 -6600 14680 -6540
rect 14620 -6680 14680 -6620
rect 14620 -6760 14680 -6700
rect 16420 -6000 16480 -5940
rect 16420 -6080 16480 -6020
rect 16420 -6160 16480 -6100
rect 17580 -6020 17640 -5960
rect 17580 -6200 17640 -6140
rect 18200 -6020 18260 -5960
rect 18200 -6200 18260 -6140
rect 18800 -6020 18860 -5960
rect 18800 -6200 18860 -6140
rect 8000 -7540 8060 -7480
rect 8080 -7540 8140 -7480
rect 8160 -7540 8220 -7480
rect 8240 -7540 8300 -7480
rect 8320 -7540 8380 -7480
rect 8400 -7540 8460 -7480
rect 8480 -7540 8540 -7480
rect 8560 -7540 8620 -7480
rect 8640 -7540 8700 -7480
rect 8720 -7540 8780 -7480
rect 8800 -7540 8860 -7480
rect 8880 -7540 8940 -7480
rect 8960 -7540 9060 -7480
rect 9080 -7540 9140 -7480
rect 8000 -7640 8060 -7580
rect 8080 -7640 8140 -7580
rect 8160 -7640 8220 -7580
rect 8240 -7640 8300 -7580
rect 8320 -7640 8380 -7580
rect 8400 -7640 8460 -7580
rect 8480 -7640 8540 -7580
rect 8560 -7640 8620 -7580
rect 8640 -7640 8700 -7580
rect 8720 -7640 8780 -7580
rect 8800 -7640 8860 -7580
rect 8880 -7640 8940 -7580
rect 8960 -7640 9060 -7580
rect 9080 -7640 9140 -7580
rect 10880 -7540 10940 -7480
rect 10980 -7540 11040 -7480
rect 10880 -7620 10940 -7560
rect 10980 -7620 11040 -7560
rect 10880 -7800 10940 -7740
rect 10980 -7800 11040 -7740
rect 10880 -7880 10940 -7820
rect 10980 -7880 11040 -7820
rect 11460 -7560 11520 -7500
rect 11540 -7560 11600 -7500
rect 11460 -7640 11520 -7580
rect 11540 -7640 11600 -7580
rect 11460 -7720 11520 -7660
rect 11540 -7720 11600 -7660
rect 11460 -7800 11520 -7740
rect 11540 -7800 11600 -7740
rect 11460 -7880 11520 -7820
rect 11540 -7880 11600 -7820
rect 12680 -7560 12740 -7500
rect 12760 -7560 12820 -7500
rect 12680 -7640 12740 -7580
rect 12760 -7640 12820 -7580
rect 12680 -7720 12740 -7660
rect 12760 -7720 12820 -7660
rect 12680 -7800 12740 -7740
rect 12760 -7800 12820 -7740
rect 12680 -7880 12740 -7820
rect 12760 -7880 12820 -7820
rect 13920 -7560 13980 -7500
rect 14000 -7560 14060 -7500
rect 13920 -7640 13980 -7580
rect 14000 -7640 14060 -7580
rect 13920 -7720 13980 -7660
rect 14000 -7720 14060 -7660
rect 13920 -7800 13980 -7740
rect 14000 -7800 14060 -7740
rect 13920 -7880 13980 -7820
rect 14000 -7880 14060 -7820
rect 15140 -7560 15200 -7500
rect 15220 -7560 15280 -7500
rect 15140 -7640 15200 -7580
rect 15220 -7640 15280 -7580
rect 15140 -7720 15200 -7660
rect 15220 -7720 15280 -7660
rect 15140 -7800 15200 -7740
rect 15220 -7800 15280 -7740
rect 15140 -7880 15200 -7820
rect 15220 -7880 15280 -7820
rect 15720 -7540 15780 -7480
rect 15820 -7540 15880 -7480
rect 15720 -7620 15780 -7560
rect 15820 -7620 15880 -7560
rect 17660 -7540 17720 -7480
rect 17740 -7540 17840 -7480
rect 17860 -7540 17920 -7480
rect 17940 -7540 18000 -7480
rect 18020 -7540 18080 -7480
rect 18100 -7540 18160 -7480
rect 18180 -7540 18240 -7480
rect 18260 -7540 18320 -7480
rect 18340 -7540 18400 -7480
rect 18420 -7540 18480 -7480
rect 18500 -7540 18560 -7480
rect 18580 -7540 18640 -7480
rect 18660 -7540 18720 -7480
rect 18740 -7540 18800 -7480
rect 17660 -7640 17720 -7580
rect 17740 -7640 17840 -7580
rect 17860 -7640 17920 -7580
rect 17940 -7640 18000 -7580
rect 18020 -7640 18080 -7580
rect 18100 -7640 18160 -7580
rect 18180 -7640 18240 -7580
rect 18260 -7640 18320 -7580
rect 18340 -7640 18400 -7580
rect 18420 -7640 18480 -7580
rect 18500 -7640 18560 -7580
rect 18580 -7640 18640 -7580
rect 18660 -7640 18720 -7580
rect 18740 -7640 18800 -7580
rect 15720 -7800 15780 -7740
rect 15820 -7800 15880 -7740
rect 15720 -7880 15780 -7820
rect 15820 -7880 15880 -7820
rect 10880 -8160 10940 -8100
rect 10980 -8160 11040 -8100
rect 10880 -8240 10940 -8180
rect 10980 -8240 11040 -8180
rect 10880 -8380 10940 -8320
rect 10980 -8380 11040 -8320
rect 10880 -8460 10940 -8400
rect 10980 -8460 11040 -8400
rect 12060 -8160 12120 -8100
rect 12160 -8160 12220 -8100
rect 12060 -8240 12120 -8180
rect 12160 -8240 12220 -8180
rect 12060 -8380 12120 -8320
rect 12160 -8380 12220 -8320
rect 12060 -8460 12120 -8400
rect 12160 -8460 12220 -8400
rect 13300 -8160 13360 -8100
rect 13400 -8160 13460 -8100
rect 13300 -8240 13360 -8180
rect 13400 -8240 13460 -8180
rect 13300 -8380 13360 -8320
rect 13400 -8380 13460 -8320
rect 13300 -8460 13360 -8400
rect 13400 -8460 13460 -8400
rect 14520 -8160 14580 -8100
rect 14620 -8160 14680 -8100
rect 14520 -8240 14580 -8180
rect 14620 -8240 14680 -8180
rect 14520 -8380 14580 -8320
rect 14620 -8380 14680 -8320
rect 14520 -8460 14580 -8400
rect 14620 -8460 14680 -8400
rect 15720 -8160 15780 -8100
rect 15820 -8160 15880 -8100
rect 15720 -8240 15780 -8180
rect 15820 -8240 15880 -8180
rect 15720 -8380 15780 -8320
rect 15820 -8380 15880 -8320
rect 15720 -8460 15780 -8400
rect 15820 -8460 15880 -8400
rect 9320 -10100 9400 -10020
rect 9460 -10100 9540 -10020
rect 9600 -10100 9680 -10020
rect 17120 -10100 17200 -10020
rect 17260 -10100 17340 -10020
rect 17400 -10100 17480 -10020
rect 9320 -10240 9400 -10160
rect 9460 -10240 9540 -10160
rect 9600 -10240 9680 -10160
rect 9320 -10380 9400 -10300
rect 9460 -10380 9540 -10300
rect 9600 -10380 9680 -10300
rect 17120 -10240 17200 -10160
rect 17260 -10240 17340 -10160
rect 17400 -10240 17480 -10160
rect 17120 -10380 17200 -10300
rect 17260 -10380 17340 -10300
rect 17400 -10380 17480 -10300
rect 13220 -10680 13280 -10620
rect 13320 -10680 13380 -10620
rect 13420 -10680 13480 -10620
rect 13520 -10680 13580 -10620
rect 13220 -10780 13280 -10720
rect 13320 -10780 13380 -10720
rect 13420 -10780 13480 -10720
rect 13520 -10780 13580 -10720
rect 13220 -10880 13280 -10820
rect 13320 -10880 13380 -10820
rect 13420 -10880 13480 -10820
rect 13520 -10880 13580 -10820
rect 13220 -10980 13280 -10920
rect 13320 -10980 13380 -10920
rect 13420 -10980 13480 -10920
rect 13520 -10980 13580 -10920
rect 8260 -11480 8320 -11420
rect 8360 -11480 8420 -11420
rect 8460 -11480 8520 -11420
rect 8560 -11480 8620 -11420
rect 8260 -11560 8320 -11500
rect 8360 -11560 8420 -11500
rect 8460 -11560 8520 -11500
rect 8560 -11560 8620 -11500
rect 8260 -11660 8320 -11600
rect 8360 -11660 8420 -11600
rect 8460 -11660 8520 -11600
rect 8560 -11660 8620 -11600
rect 8260 -11760 8320 -11700
rect 8360 -11760 8420 -11700
rect 8460 -11760 8520 -11700
rect 8560 -11760 8620 -11700
rect 18180 -11480 18240 -11420
rect 18280 -11480 18340 -11420
rect 18380 -11480 18440 -11420
rect 18480 -11480 18540 -11420
rect 18180 -11560 18240 -11500
rect 18280 -11560 18340 -11500
rect 18380 -11560 18440 -11500
rect 18480 -11560 18540 -11500
rect 18180 -11660 18240 -11600
rect 18280 -11660 18340 -11600
rect 18380 -11660 18440 -11600
rect 18480 -11660 18540 -11600
rect 18180 -11760 18240 -11700
rect 18280 -11760 18340 -11700
rect 18380 -11760 18440 -11700
rect 18480 -11760 18540 -11700
<< metal2 >>
rect 11320 -1980 15340 -1960
rect 11320 -2040 11400 -1980
rect 11460 -2040 11500 -1980
rect 11560 -2040 12640 -1980
rect 12700 -2040 12740 -1980
rect 12800 -2040 13220 -1980
rect 11320 -2060 13220 -2040
rect 13300 -2060 13360 -1980
rect 13440 -2060 13500 -1980
rect 13580 -2040 13860 -1980
rect 13920 -2040 13960 -1980
rect 14020 -2040 15100 -1980
rect 15160 -2040 15200 -1980
rect 15260 -2040 15340 -1980
rect 13580 -2060 15340 -2040
rect 11320 -2120 11400 -2060
rect 11460 -2120 11500 -2060
rect 11560 -2120 12640 -2060
rect 12700 -2120 12740 -2060
rect 12800 -2100 13860 -2060
rect 12800 -2120 13220 -2100
rect 11320 -2180 13220 -2120
rect 13300 -2180 13360 -2100
rect 13440 -2180 13500 -2100
rect 13580 -2120 13860 -2100
rect 13920 -2120 13960 -2060
rect 14020 -2120 15100 -2060
rect 15160 -2120 15200 -2060
rect 15260 -2120 15340 -2060
rect 13580 -2180 15340 -2120
rect 11320 -2240 11400 -2180
rect 11460 -2240 11500 -2180
rect 11560 -2240 12640 -2180
rect 12700 -2240 12740 -2180
rect 12800 -2240 13860 -2180
rect 13920 -2240 13960 -2180
rect 14020 -2240 15100 -2180
rect 15160 -2240 15200 -2180
rect 15260 -2240 15340 -2180
rect 11320 -2260 13220 -2240
rect 11320 -2320 11400 -2260
rect 11460 -2320 11500 -2260
rect 11560 -2320 12640 -2260
rect 12700 -2320 12740 -2260
rect 12800 -2320 13220 -2260
rect 13300 -2320 13360 -2240
rect 13440 -2320 13500 -2240
rect 13580 -2260 15340 -2240
rect 13580 -2320 13860 -2260
rect 13920 -2320 13960 -2260
rect 14020 -2320 15100 -2260
rect 15160 -2320 15200 -2260
rect 15260 -2320 15340 -2260
rect 11320 -2340 15340 -2320
rect 7360 -2880 10140 -2860
rect 7360 -2940 7400 -2880
rect 7460 -2940 8000 -2880
rect 8060 -2940 8280 -2880
rect 8340 -2940 8400 -2880
rect 8480 -2940 8540 -2880
rect 8600 -2940 8640 -2880
rect 8700 -2940 9240 -2880
rect 9300 -2940 9880 -2880
rect 9940 -2940 10140 -2880
rect 16640 -2880 19420 -2860
rect 7360 -3060 10140 -2940
rect 7360 -3120 7400 -3060
rect 7460 -3120 8000 -3060
rect 8060 -3120 8280 -3060
rect 8340 -3120 8400 -3060
rect 8480 -3120 8540 -3060
rect 8600 -3120 8640 -3060
rect 8700 -3120 9240 -3060
rect 9300 -3120 9880 -3060
rect 9940 -3120 10140 -3060
rect 7360 -3140 10140 -3120
rect 10320 -2940 16460 -2920
rect 10320 -3020 10740 -2940
rect 10820 -3020 10880 -2940
rect 10960 -3020 11020 -2940
rect 11100 -3020 11140 -2940
rect 11220 -3020 11260 -2940
rect 11340 -3020 11380 -2940
rect 11460 -3020 11500 -2940
rect 11580 -3020 11620 -2940
rect 11700 -3020 11740 -2940
rect 11820 -3020 11860 -2940
rect 11940 -3020 11980 -2940
rect 12060 -3020 12100 -2940
rect 12180 -3020 12220 -2940
rect 12300 -3020 12340 -2940
rect 12420 -3020 12460 -2940
rect 12540 -3020 12580 -2940
rect 12660 -3020 12700 -2940
rect 12780 -3020 12820 -2940
rect 12900 -3020 12940 -2940
rect 13020 -3020 13060 -2940
rect 13140 -3020 13180 -2940
rect 13260 -3020 13300 -2940
rect 13380 -3020 13420 -2940
rect 13500 -3020 13540 -2940
rect 13620 -3020 13660 -2940
rect 13740 -3020 13780 -2940
rect 13860 -3020 13900 -2940
rect 13980 -3020 14020 -2940
rect 14100 -3020 14140 -2940
rect 14220 -3020 14260 -2940
rect 14340 -3020 14380 -2940
rect 14460 -3020 14500 -2940
rect 14580 -3020 14620 -2940
rect 14700 -3020 14740 -2940
rect 14820 -3020 14860 -2940
rect 14940 -3020 14980 -2940
rect 15060 -3020 15100 -2940
rect 15180 -3020 15220 -2940
rect 15300 -3020 15340 -2940
rect 15420 -3020 15460 -2940
rect 15540 -3020 15580 -2940
rect 15660 -3020 15700 -2940
rect 15780 -3020 15840 -2940
rect 15920 -3020 15980 -2940
rect 16060 -3020 16460 -2940
rect 10320 -3080 16460 -3020
rect 10320 -3160 10740 -3080
rect 10820 -3160 10880 -3080
rect 10960 -3160 11020 -3080
rect 11100 -3160 11140 -3080
rect 11220 -3160 11260 -3080
rect 11340 -3160 11380 -3080
rect 11460 -3160 11500 -3080
rect 11580 -3160 11620 -3080
rect 11700 -3160 11740 -3080
rect 11820 -3160 11860 -3080
rect 11940 -3160 11980 -3080
rect 12060 -3160 12100 -3080
rect 12180 -3160 12220 -3080
rect 12300 -3160 12340 -3080
rect 12420 -3160 12460 -3080
rect 12540 -3160 12580 -3080
rect 12660 -3160 12700 -3080
rect 12780 -3160 12820 -3080
rect 12900 -3160 12940 -3080
rect 13020 -3160 13060 -3080
rect 13140 -3160 13180 -3080
rect 13260 -3160 13300 -3080
rect 13380 -3160 13420 -3080
rect 13500 -3160 13540 -3080
rect 13620 -3160 13660 -3080
rect 13740 -3160 13780 -3080
rect 13860 -3160 13900 -3080
rect 13980 -3160 14020 -3080
rect 14100 -3160 14140 -3080
rect 14220 -3160 14260 -3080
rect 14340 -3160 14380 -3080
rect 14460 -3160 14500 -3080
rect 14580 -3160 14620 -3080
rect 14700 -3160 14740 -3080
rect 14820 -3160 14860 -3080
rect 14940 -3160 14980 -3080
rect 15060 -3160 15100 -3080
rect 15180 -3160 15220 -3080
rect 15300 -3160 15340 -3080
rect 15420 -3160 15460 -3080
rect 15540 -3160 15580 -3080
rect 15660 -3160 15700 -3080
rect 15780 -3160 15840 -3080
rect 15920 -3160 15980 -3080
rect 16060 -3160 16460 -3080
rect 16640 -2940 16840 -2880
rect 16900 -2940 17440 -2880
rect 17500 -2940 18080 -2880
rect 18140 -2940 18200 -2880
rect 18260 -2940 18320 -2880
rect 18400 -2940 18460 -2880
rect 18520 -2940 18680 -2880
rect 18740 -2940 19300 -2880
rect 19360 -2940 19420 -2880
rect 16640 -3060 19420 -2940
rect 16640 -3120 16840 -3060
rect 16900 -3120 17440 -3060
rect 17500 -3120 18080 -3060
rect 18140 -3120 18200 -3060
rect 18260 -3120 18320 -3060
rect 18400 -3120 18460 -3060
rect 18520 -3120 18680 -3060
rect 18740 -3120 19300 -3060
rect 19360 -3120 19420 -3060
rect 16640 -3140 19420 -3120
rect 10320 -3220 16460 -3160
rect 10320 -3300 10740 -3220
rect 10820 -3300 10880 -3220
rect 10960 -3300 11020 -3220
rect 11100 -3300 11140 -3220
rect 11220 -3300 11260 -3220
rect 11340 -3300 11380 -3220
rect 11460 -3300 11500 -3220
rect 11580 -3300 11620 -3220
rect 11700 -3300 11740 -3220
rect 11820 -3300 11860 -3220
rect 11940 -3300 11980 -3220
rect 12060 -3300 12100 -3220
rect 12180 -3300 12220 -3220
rect 12300 -3300 12340 -3220
rect 12420 -3300 12460 -3220
rect 12540 -3300 12580 -3220
rect 12660 -3300 12700 -3220
rect 12780 -3300 12820 -3220
rect 12900 -3300 12940 -3220
rect 13020 -3300 13060 -3220
rect 13140 -3300 13180 -3220
rect 13260 -3300 13300 -3220
rect 13380 -3300 13420 -3220
rect 13500 -3300 13540 -3220
rect 13620 -3300 13660 -3220
rect 13740 -3300 13780 -3220
rect 13860 -3300 13900 -3220
rect 13980 -3300 14020 -3220
rect 14100 -3300 14140 -3220
rect 14220 -3300 14260 -3220
rect 14340 -3300 14380 -3220
rect 14460 -3300 14500 -3220
rect 14580 -3300 14620 -3220
rect 14700 -3300 14740 -3220
rect 14820 -3300 14860 -3220
rect 14940 -3300 14980 -3220
rect 15060 -3300 15100 -3220
rect 15180 -3300 15220 -3220
rect 15300 -3300 15340 -3220
rect 15420 -3300 15460 -3220
rect 15540 -3300 15580 -3220
rect 15660 -3300 15700 -3220
rect 15780 -3300 15840 -3220
rect 15920 -3300 15980 -3220
rect 16060 -3300 16460 -3220
rect 10320 -3320 16460 -3300
rect 7460 -3420 19320 -3400
rect 7460 -3500 7480 -3420
rect 7560 -3500 7580 -3420
rect 7660 -3500 7680 -3420
rect 7760 -3500 7780 -3420
rect 7860 -3500 7880 -3420
rect 7960 -3500 7980 -3420
rect 8060 -3500 8080 -3420
rect 8160 -3500 8180 -3420
rect 8260 -3500 8280 -3420
rect 8360 -3500 8380 -3420
rect 8460 -3500 8480 -3420
rect 8560 -3500 8580 -3420
rect 8660 -3500 8680 -3420
rect 8760 -3500 8780 -3420
rect 8860 -3500 8880 -3420
rect 8960 -3500 8980 -3420
rect 9060 -3500 9080 -3420
rect 9160 -3500 9180 -3420
rect 9260 -3500 9280 -3420
rect 9360 -3500 9380 -3420
rect 9460 -3500 9480 -3420
rect 9560 -3500 9580 -3420
rect 9660 -3500 9680 -3420
rect 9760 -3500 9780 -3420
rect 9860 -3480 10020 -3420
rect 10080 -3480 10120 -3420
rect 10180 -3480 10260 -3420
rect 10340 -3480 10420 -3420
rect 10480 -3480 10520 -3420
rect 10580 -3480 11720 -3420
rect 9860 -3500 11720 -3480
rect 11800 -3500 11860 -3420
rect 11940 -3500 12000 -3420
rect 12080 -3500 13220 -3420
rect 13300 -3500 13360 -3420
rect 13440 -3500 13500 -3420
rect 13580 -3500 14720 -3420
rect 14800 -3500 14860 -3420
rect 14940 -3500 15000 -3420
rect 15080 -3480 16220 -3420
rect 16280 -3480 16320 -3420
rect 16380 -3480 16460 -3420
rect 16540 -3480 16620 -3420
rect 16680 -3480 16720 -3420
rect 16780 -3480 16920 -3420
rect 15080 -3500 16920 -3480
rect 17000 -3500 17020 -3420
rect 17100 -3500 17120 -3420
rect 17200 -3500 17220 -3420
rect 17300 -3500 17320 -3420
rect 17400 -3500 17420 -3420
rect 17500 -3500 17520 -3420
rect 17600 -3500 17620 -3420
rect 17700 -3500 17720 -3420
rect 17800 -3500 17820 -3420
rect 17900 -3500 17920 -3420
rect 18000 -3500 18020 -3420
rect 18100 -3500 18120 -3420
rect 18200 -3500 18220 -3420
rect 18300 -3500 18320 -3420
rect 18400 -3500 18420 -3420
rect 18500 -3500 18520 -3420
rect 18600 -3500 18620 -3420
rect 18700 -3500 18720 -3420
rect 18800 -3500 18820 -3420
rect 18900 -3500 18920 -3420
rect 19000 -3500 19020 -3420
rect 19100 -3500 19120 -3420
rect 19200 -3500 19220 -3420
rect 19300 -3500 19320 -3420
rect 7460 -3560 19320 -3500
rect 7460 -3640 7480 -3560
rect 7560 -3640 7580 -3560
rect 7660 -3640 7680 -3560
rect 7760 -3640 7780 -3560
rect 7860 -3640 7880 -3560
rect 7960 -3640 7980 -3560
rect 8060 -3640 8080 -3560
rect 8160 -3640 8180 -3560
rect 8260 -3640 8280 -3560
rect 8360 -3640 8380 -3560
rect 8460 -3640 8480 -3560
rect 8560 -3640 8580 -3560
rect 8660 -3640 8680 -3560
rect 8760 -3640 8780 -3560
rect 8860 -3640 8880 -3560
rect 8960 -3640 8980 -3560
rect 9060 -3640 9080 -3560
rect 9160 -3640 9180 -3560
rect 9260 -3640 9280 -3560
rect 9360 -3640 9380 -3560
rect 9460 -3640 9480 -3560
rect 9560 -3640 9580 -3560
rect 9660 -3640 9680 -3560
rect 9760 -3640 9780 -3560
rect 9860 -3640 10020 -3560
rect 10100 -3640 10140 -3560
rect 10200 -3640 10260 -3560
rect 10340 -3640 10400 -3560
rect 10460 -3640 10500 -3560
rect 10580 -3640 11720 -3560
rect 11800 -3640 11860 -3560
rect 11940 -3640 12000 -3560
rect 12080 -3640 13220 -3560
rect 13300 -3640 13360 -3560
rect 13440 -3640 13500 -3560
rect 13580 -3640 14720 -3560
rect 14800 -3640 14860 -3560
rect 14940 -3640 15000 -3560
rect 15080 -3640 16220 -3560
rect 16300 -3640 16340 -3560
rect 16400 -3640 16460 -3560
rect 16540 -3640 16600 -3560
rect 16660 -3640 16700 -3560
rect 16780 -3640 16920 -3560
rect 17000 -3640 17020 -3560
rect 17100 -3640 17120 -3560
rect 17200 -3640 17220 -3560
rect 17300 -3640 17320 -3560
rect 17400 -3640 17420 -3560
rect 17500 -3640 17520 -3560
rect 17600 -3640 17620 -3560
rect 17700 -3640 17720 -3560
rect 17800 -3640 17820 -3560
rect 17900 -3640 17920 -3560
rect 18000 -3640 18020 -3560
rect 18100 -3640 18120 -3560
rect 18200 -3640 18220 -3560
rect 18300 -3640 18320 -3560
rect 18400 -3640 18420 -3560
rect 18500 -3640 18520 -3560
rect 18600 -3640 18620 -3560
rect 18700 -3640 18720 -3560
rect 18800 -3640 18820 -3560
rect 18900 -3640 18920 -3560
rect 19000 -3640 19020 -3560
rect 19100 -3640 19120 -3560
rect 19200 -3640 19220 -3560
rect 19300 -3640 19320 -3560
rect 7460 -3700 19320 -3640
rect 7460 -3780 7480 -3700
rect 7560 -3780 7580 -3700
rect 7660 -3780 7680 -3700
rect 7760 -3780 7780 -3700
rect 7860 -3780 7880 -3700
rect 7960 -3780 7980 -3700
rect 8060 -3780 8080 -3700
rect 8160 -3780 8180 -3700
rect 8260 -3780 8280 -3700
rect 8360 -3780 8380 -3700
rect 8460 -3780 8480 -3700
rect 8560 -3780 8580 -3700
rect 8660 -3780 8680 -3700
rect 8760 -3780 8780 -3700
rect 8860 -3780 8880 -3700
rect 8960 -3780 8980 -3700
rect 9060 -3780 9080 -3700
rect 9160 -3780 9180 -3700
rect 9260 -3780 9280 -3700
rect 9360 -3780 9380 -3700
rect 9460 -3780 9480 -3700
rect 9560 -3780 9580 -3700
rect 9660 -3780 9680 -3700
rect 9760 -3780 9780 -3700
rect 9860 -3720 11720 -3700
rect 9860 -3780 10020 -3720
rect 10080 -3780 10120 -3720
rect 10180 -3780 10260 -3720
rect 10340 -3780 10420 -3720
rect 10480 -3780 10520 -3720
rect 10580 -3780 11720 -3720
rect 11800 -3780 11860 -3700
rect 11940 -3780 12000 -3700
rect 12080 -3780 13220 -3700
rect 13300 -3780 13360 -3700
rect 13440 -3780 13500 -3700
rect 13580 -3780 14720 -3700
rect 14800 -3780 14860 -3700
rect 14940 -3780 15000 -3700
rect 15080 -3720 16920 -3700
rect 15080 -3780 16220 -3720
rect 16280 -3780 16320 -3720
rect 16380 -3780 16460 -3720
rect 16540 -3780 16620 -3720
rect 16680 -3780 16720 -3720
rect 16780 -3780 16920 -3720
rect 17000 -3780 17020 -3700
rect 17100 -3780 17120 -3700
rect 17200 -3780 17220 -3700
rect 17300 -3780 17320 -3700
rect 17400 -3780 17420 -3700
rect 17500 -3780 17520 -3700
rect 17600 -3780 17620 -3700
rect 17700 -3780 17720 -3700
rect 17800 -3780 17820 -3700
rect 17900 -3780 17920 -3700
rect 18000 -3780 18020 -3700
rect 18100 -3780 18120 -3700
rect 18200 -3780 18220 -3700
rect 18300 -3780 18320 -3700
rect 18400 -3780 18420 -3700
rect 18500 -3780 18520 -3700
rect 18600 -3780 18620 -3700
rect 18700 -3780 18720 -3700
rect 18800 -3780 18820 -3700
rect 18900 -3780 18920 -3700
rect 19000 -3780 19020 -3700
rect 19100 -3780 19120 -3700
rect 19200 -3780 19220 -3700
rect 19300 -3780 19320 -3700
rect 7460 -3800 19320 -3780
rect 13200 -3900 13600 -3880
rect 7180 -3960 8920 -3940
rect 7180 -4020 8360 -3960
rect 8420 -4020 8820 -3960
rect 8880 -4020 8920 -3960
rect 7180 -4040 7340 -4020
rect 7180 -4100 7220 -4040
rect 7300 -4080 7340 -4040
rect 7400 -4040 7600 -4020
rect 7400 -4080 7460 -4040
rect 7300 -4100 7460 -4080
rect 7540 -4080 7600 -4040
rect 7660 -4040 8920 -4020
rect 7660 -4080 7700 -4040
rect 7540 -4100 7700 -4080
rect 7780 -4100 8920 -4040
rect 7180 -4140 8920 -4100
rect 7180 -4200 7220 -4140
rect 7300 -4200 7340 -4140
rect 7400 -4200 7460 -4140
rect 7540 -4200 7600 -4140
rect 7660 -4200 7700 -4140
rect 7780 -4200 8360 -4140
rect 8420 -4200 8820 -4140
rect 8880 -4200 8920 -4140
rect 7180 -4220 8920 -4200
rect 13200 -3980 13220 -3900
rect 13300 -3980 13360 -3900
rect 13440 -3980 13500 -3900
rect 13580 -3980 13600 -3900
rect 13200 -4020 13600 -3980
rect 13200 -4100 13220 -4020
rect 13300 -4100 13360 -4020
rect 13440 -4100 13500 -4020
rect 13580 -4100 13600 -4020
rect 13200 -4140 13600 -4100
rect 13200 -4220 13220 -4140
rect 13300 -4220 13360 -4140
rect 13440 -4220 13500 -4140
rect 13580 -4220 13600 -4140
rect 17940 -3960 19680 -3940
rect 17940 -4020 17960 -3960
rect 18020 -4020 18420 -3960
rect 18480 -4020 19680 -3960
rect 17940 -4040 19140 -4020
rect 17940 -4100 19020 -4040
rect 19100 -4080 19140 -4040
rect 19200 -4040 19400 -4020
rect 19200 -4080 19260 -4040
rect 19100 -4100 19260 -4080
rect 19340 -4080 19400 -4040
rect 19460 -4040 19680 -4020
rect 19460 -4080 19500 -4040
rect 19340 -4100 19500 -4080
rect 19580 -4100 19680 -4040
rect 17940 -4140 19680 -4100
rect 17940 -4200 17960 -4140
rect 18020 -4200 18420 -4140
rect 18480 -4200 19020 -4140
rect 19100 -4200 19140 -4140
rect 19200 -4200 19260 -4140
rect 19340 -4200 19400 -4140
rect 19460 -4200 19500 -4140
rect 19580 -4200 19680 -4140
rect 17940 -4220 19680 -4200
rect 13200 -4260 13600 -4220
rect 13200 -4340 13220 -4260
rect 13300 -4340 13360 -4260
rect 13440 -4340 13500 -4260
rect 13580 -4340 13600 -4260
rect 13200 -4380 13600 -4340
rect 10300 -4420 11100 -4400
rect 8240 -4440 8740 -4420
rect 8240 -4500 8420 -4440
rect 8480 -4500 8520 -4440
rect 8580 -4500 8620 -4440
rect 8680 -4500 8740 -4440
rect 8240 -4540 8740 -4500
rect 8240 -4600 8420 -4540
rect 8480 -4600 8520 -4540
rect 8580 -4600 8620 -4540
rect 8680 -4600 8740 -4540
rect 8240 -4620 8740 -4600
rect 10280 -4440 10740 -4420
rect 10280 -4500 10300 -4440
rect 10360 -4500 10620 -4440
rect 10680 -4500 10740 -4440
rect 10820 -4500 10860 -4420
rect 10960 -4500 11000 -4420
rect 11080 -4500 11100 -4420
rect 10280 -4520 11100 -4500
rect 10280 -4580 10300 -4520
rect 10360 -4580 10620 -4520
rect 10680 -4580 11100 -4520
rect 10280 -4600 11100 -4580
rect 10280 -4660 10300 -4600
rect 10360 -4660 10620 -4600
rect 10680 -4660 10740 -4600
rect 10280 -4680 10740 -4660
rect 10820 -4680 10860 -4600
rect 10960 -4680 11000 -4600
rect 11080 -4680 11100 -4600
rect 10300 -4700 11100 -4680
rect 11700 -4420 12480 -4400
rect 11700 -4500 11720 -4420
rect 11800 -4500 11840 -4420
rect 11960 -4500 12000 -4420
rect 12080 -4440 12500 -4420
rect 12080 -4500 12100 -4440
rect 12160 -4500 12420 -4440
rect 12480 -4500 12500 -4440
rect 11700 -4520 12500 -4500
rect 11700 -4580 12100 -4520
rect 12160 -4580 12420 -4520
rect 12480 -4580 12500 -4520
rect 11700 -4600 12500 -4580
rect 11700 -4680 11720 -4600
rect 11800 -4680 11840 -4600
rect 11960 -4680 12000 -4600
rect 12080 -4660 12100 -4600
rect 12160 -4660 12420 -4600
rect 12480 -4660 12500 -4600
rect 12080 -4680 12500 -4660
rect 13200 -4460 13220 -4380
rect 13300 -4460 13360 -4380
rect 13440 -4460 13500 -4380
rect 13580 -4460 13600 -4380
rect 14300 -4420 15100 -4400
rect 13200 -4500 13600 -4460
rect 13200 -4580 13220 -4500
rect 13300 -4580 13360 -4500
rect 13440 -4580 13500 -4500
rect 13580 -4580 13600 -4500
rect 13200 -4620 13600 -4580
rect 11700 -4700 12480 -4680
rect 13200 -4700 13220 -4620
rect 13300 -4700 13360 -4620
rect 13440 -4700 13500 -4620
rect 13580 -4700 13600 -4620
rect 14280 -4440 14720 -4420
rect 14280 -4500 14300 -4440
rect 14360 -4500 14620 -4440
rect 14680 -4500 14720 -4440
rect 14800 -4500 14840 -4420
rect 14960 -4500 15000 -4420
rect 15080 -4500 15100 -4420
rect 14280 -4520 15100 -4500
rect 14280 -4580 14300 -4520
rect 14360 -4580 14620 -4520
rect 14680 -4580 15100 -4520
rect 14280 -4600 15100 -4580
rect 14280 -4660 14300 -4600
rect 14360 -4660 14620 -4600
rect 14680 -4660 14720 -4600
rect 14280 -4680 14720 -4660
rect 14800 -4680 14840 -4600
rect 14960 -4680 15000 -4600
rect 15080 -4680 15100 -4600
rect 14300 -4700 15100 -4680
rect 15700 -4420 16480 -4400
rect 15700 -4500 15720 -4420
rect 15800 -4500 15840 -4420
rect 15940 -4500 15980 -4420
rect 16060 -4440 16500 -4420
rect 16060 -4500 16100 -4440
rect 16160 -4500 16420 -4440
rect 16480 -4500 16500 -4440
rect 15700 -4520 16500 -4500
rect 15700 -4580 16100 -4520
rect 16160 -4580 16420 -4520
rect 16480 -4580 16500 -4520
rect 15700 -4600 16500 -4580
rect 15700 -4680 15720 -4600
rect 15800 -4680 15840 -4600
rect 15940 -4680 15980 -4600
rect 16060 -4660 16100 -4600
rect 16160 -4660 16420 -4600
rect 16480 -4660 16500 -4600
rect 18060 -4440 18560 -4420
rect 18060 -4500 18140 -4440
rect 18200 -4500 18260 -4440
rect 18320 -4500 18360 -4440
rect 18420 -4500 18560 -4440
rect 18060 -4540 18560 -4500
rect 18060 -4600 18140 -4540
rect 18200 -4600 18260 -4540
rect 18320 -4600 18360 -4540
rect 18420 -4600 18560 -4540
rect 18060 -4620 18560 -4600
rect 16060 -4680 16500 -4660
rect 15700 -4700 16480 -4680
rect 13200 -4740 13600 -4700
rect 13200 -4820 13220 -4740
rect 13300 -4820 13360 -4740
rect 13440 -4820 13500 -4740
rect 13580 -4820 13600 -4740
rect 13200 -4860 13600 -4820
rect 12920 -4920 13100 -4900
rect 12920 -5060 12940 -4920
rect 13080 -5060 13100 -4920
rect 9300 -5100 9660 -5080
rect 9300 -5180 9320 -5100
rect 9400 -5180 9440 -5100
rect 9520 -5180 9560 -5100
rect 9640 -5180 9660 -5100
rect 9300 -5220 9660 -5180
rect 9300 -5280 9320 -5220
rect 9380 -5280 9440 -5220
rect 9520 -5280 9580 -5220
rect 9640 -5240 9660 -5220
rect 10360 -5120 10620 -5100
rect 10360 -5180 10380 -5120
rect 10440 -5180 10540 -5120
rect 10600 -5180 10620 -5120
rect 10360 -5240 10620 -5180
rect 11440 -5120 12420 -5100
rect 11500 -5180 11540 -5120
rect 11600 -5180 12180 -5120
rect 12240 -5180 12340 -5120
rect 12400 -5180 12420 -5120
rect 11440 -5200 12420 -5180
rect 12920 -5240 13100 -5060
rect 9640 -5260 13100 -5240
rect 9640 -5280 11200 -5260
rect 9300 -5320 11200 -5280
rect 11260 -5320 13100 -5260
rect 9300 -5400 9320 -5320
rect 9400 -5400 9440 -5320
rect 9520 -5400 9560 -5320
rect 9640 -5340 13100 -5320
rect 9640 -5400 11280 -5340
rect 11340 -5400 13100 -5340
rect 9300 -5420 13100 -5400
rect 13200 -4940 13220 -4860
rect 13300 -4940 13360 -4860
rect 13440 -4940 13500 -4860
rect 13580 -4940 13600 -4860
rect 13200 -4980 13600 -4940
rect 13200 -5060 13220 -4980
rect 13300 -5060 13360 -4980
rect 13440 -5060 13500 -4980
rect 13580 -5060 13600 -4980
rect 13200 -5100 13600 -5060
rect 13200 -5180 13220 -5100
rect 13300 -5180 13360 -5100
rect 13440 -5180 13500 -5100
rect 13580 -5180 13600 -5100
rect 13200 -5220 13600 -5180
rect 13200 -5300 13220 -5220
rect 13300 -5300 13360 -5220
rect 13440 -5300 13500 -5220
rect 13580 -5300 13600 -5220
rect 13200 -5340 13600 -5300
rect 13200 -5420 13220 -5340
rect 13300 -5420 13360 -5340
rect 13440 -5420 13500 -5340
rect 13580 -5420 13600 -5340
rect 13700 -4920 13880 -4900
rect 13700 -5060 13720 -4920
rect 13860 -5060 13880 -4920
rect 13700 -5240 13880 -5060
rect 14360 -5120 15360 -5100
rect 14360 -5180 14380 -5120
rect 14440 -5180 14540 -5120
rect 14600 -5180 15200 -5120
rect 15260 -5180 15300 -5120
rect 14360 -5200 15360 -5180
rect 16160 -5120 16420 -5100
rect 16160 -5180 16180 -5120
rect 16240 -5180 16340 -5120
rect 16400 -5180 16420 -5120
rect 16160 -5240 16420 -5180
rect 17140 -5240 17500 -5080
rect 13700 -5260 17500 -5240
rect 13700 -5320 15540 -5260
rect 15600 -5320 17500 -5260
rect 13700 -5340 17500 -5320
rect 13700 -5400 15460 -5340
rect 15520 -5400 17500 -5340
rect 13700 -5420 17500 -5400
rect 13200 -5460 13600 -5420
rect 9300 -5500 13100 -5480
rect 9300 -5560 11540 -5500
rect 11600 -5560 13100 -5500
rect 9300 -5580 13100 -5560
rect 9300 -5640 11460 -5580
rect 11520 -5640 13100 -5580
rect 9300 -5660 13100 -5640
rect 9300 -5820 9660 -5660
rect 10360 -5720 10620 -5660
rect 10360 -5780 10380 -5720
rect 10440 -5780 10540 -5720
rect 10600 -5780 10620 -5720
rect 10360 -5800 10620 -5780
rect 11180 -5720 12420 -5700
rect 11180 -5780 11200 -5720
rect 11260 -5780 11300 -5720
rect 11360 -5780 12180 -5720
rect 12240 -5780 12340 -5720
rect 12400 -5780 12420 -5720
rect 11180 -5800 12420 -5780
rect 12920 -5840 13100 -5660
rect 10300 -5920 12100 -5900
rect 10280 -5940 11720 -5920
rect 7720 -5960 9420 -5940
rect 7720 -6020 7920 -5960
rect 7980 -6020 8280 -5960
rect 8340 -6020 8400 -5960
rect 8460 -6020 8540 -5960
rect 8600 -6020 9140 -5960
rect 9200 -6020 9420 -5960
rect 7720 -6140 9420 -6020
rect 7720 -6200 7920 -6140
rect 7980 -6200 8280 -6140
rect 8340 -6200 8400 -6140
rect 8460 -6200 8540 -6140
rect 8600 -6200 9140 -6140
rect 9200 -6200 9420 -6140
rect 10280 -6000 10300 -5940
rect 10360 -6000 10620 -5940
rect 10680 -6000 11720 -5940
rect 11800 -6000 11840 -5920
rect 11960 -6000 12000 -5920
rect 12080 -6000 12100 -5920
rect 12920 -5980 12940 -5840
rect 13080 -5980 13100 -5840
rect 12920 -6000 13100 -5980
rect 13200 -5540 13220 -5460
rect 13300 -5540 13360 -5460
rect 13440 -5540 13500 -5460
rect 13580 -5540 13600 -5460
rect 13200 -5580 13600 -5540
rect 13200 -5660 13220 -5580
rect 13300 -5660 13360 -5580
rect 13440 -5660 13500 -5580
rect 13580 -5660 13600 -5580
rect 13200 -5700 13600 -5660
rect 13200 -5780 13220 -5700
rect 13300 -5780 13360 -5700
rect 13440 -5780 13500 -5700
rect 13580 -5780 13600 -5700
rect 13200 -5820 13600 -5780
rect 13200 -5900 13220 -5820
rect 13300 -5900 13360 -5820
rect 13440 -5900 13500 -5820
rect 13580 -5900 13600 -5820
rect 13200 -5940 13600 -5900
rect 10280 -6020 12100 -6000
rect 10280 -6080 10300 -6020
rect 10360 -6080 10620 -6020
rect 10680 -6080 12100 -6020
rect 10280 -6100 12100 -6080
rect 10280 -6160 10300 -6100
rect 10360 -6160 10620 -6100
rect 10680 -6160 11720 -6100
rect 10280 -6180 11720 -6160
rect 11800 -6180 11840 -6100
rect 11960 -6180 12000 -6100
rect 12080 -6180 12100 -6100
rect 10300 -6200 12100 -6180
rect 13200 -6020 13220 -5940
rect 13300 -6020 13360 -5940
rect 13440 -6020 13500 -5940
rect 13580 -6020 13600 -5940
rect 13700 -5500 17500 -5480
rect 13700 -5560 15200 -5500
rect 15260 -5560 17160 -5500
rect 13700 -5580 17160 -5560
rect 17240 -5580 17280 -5500
rect 17360 -5580 17400 -5500
rect 17480 -5580 17500 -5500
rect 13700 -5640 15280 -5580
rect 15340 -5620 17500 -5580
rect 15340 -5640 17160 -5620
rect 13700 -5660 17160 -5640
rect 13700 -5840 13880 -5660
rect 14360 -5720 15620 -5700
rect 14360 -5780 14380 -5720
rect 14440 -5780 14540 -5720
rect 14600 -5780 15440 -5720
rect 15500 -5780 15540 -5720
rect 15600 -5780 15620 -5720
rect 14360 -5800 15620 -5780
rect 16160 -5720 16420 -5660
rect 16160 -5780 16180 -5720
rect 16240 -5780 16340 -5720
rect 16400 -5780 16420 -5720
rect 16160 -5800 16420 -5780
rect 17140 -5680 17160 -5660
rect 17240 -5680 17280 -5620
rect 17360 -5680 17400 -5620
rect 17480 -5680 17500 -5620
rect 17140 -5720 17500 -5680
rect 17140 -5800 17160 -5720
rect 17240 -5800 17280 -5720
rect 17360 -5800 17400 -5720
rect 17480 -5800 17500 -5720
rect 17140 -5820 17500 -5800
rect 13700 -5980 13720 -5840
rect 13860 -5980 13880 -5840
rect 13700 -6000 13880 -5980
rect 14700 -5920 16480 -5900
rect 14700 -6000 14720 -5920
rect 14800 -6000 14840 -5920
rect 14960 -6000 15000 -5920
rect 15080 -5940 16500 -5920
rect 15080 -6000 16100 -5940
rect 16160 -6000 16420 -5940
rect 16480 -6000 16500 -5940
rect 13200 -6060 13600 -6020
rect 13200 -6140 13220 -6060
rect 13300 -6140 13360 -6060
rect 13440 -6140 13500 -6060
rect 13580 -6140 13600 -6060
rect 13200 -6180 13600 -6140
rect 7720 -6220 9420 -6200
rect 13200 -6260 13220 -6180
rect 13300 -6260 13360 -6180
rect 13440 -6260 13500 -6180
rect 13580 -6260 13600 -6180
rect 14700 -6020 16500 -6000
rect 14700 -6080 16100 -6020
rect 16160 -6080 16420 -6020
rect 16480 -6080 16500 -6020
rect 14700 -6100 16500 -6080
rect 14700 -6180 14720 -6100
rect 14800 -6180 14840 -6100
rect 14960 -6180 15000 -6100
rect 15080 -6160 16100 -6100
rect 16160 -6160 16420 -6100
rect 16480 -6160 16500 -6100
rect 15080 -6180 16500 -6160
rect 17380 -5960 19080 -5940
rect 17380 -6020 17580 -5960
rect 17640 -6020 18200 -5960
rect 18260 -6020 18340 -5960
rect 18400 -6020 18460 -5960
rect 18520 -6020 18800 -5960
rect 18860 -6020 19080 -5960
rect 17380 -6140 19080 -6020
rect 14700 -6200 16480 -6180
rect 17380 -6200 17580 -6140
rect 17640 -6200 18200 -6140
rect 18260 -6200 18340 -6140
rect 18400 -6200 18460 -6140
rect 18520 -6200 18800 -6140
rect 18860 -6200 19080 -6140
rect 17380 -6220 19080 -6200
rect 13200 -6300 13600 -6260
rect 13200 -6380 13220 -6300
rect 13300 -6380 13360 -6300
rect 13440 -6380 13500 -6300
rect 13580 -6380 13600 -6300
rect 13200 -6420 13600 -6380
rect 13200 -6500 13220 -6420
rect 13300 -6500 13360 -6420
rect 13440 -6500 13500 -6420
rect 13580 -6500 13600 -6420
rect 10700 -6520 12480 -6500
rect 10700 -6600 10740 -6520
rect 10820 -6600 10860 -6520
rect 10980 -6600 11020 -6520
rect 11100 -6540 12500 -6520
rect 11100 -6600 12100 -6540
rect 12160 -6600 12420 -6540
rect 12480 -6600 12500 -6540
rect 10700 -6620 12500 -6600
rect 10700 -6680 12100 -6620
rect 12160 -6680 12420 -6620
rect 12480 -6680 12500 -6620
rect 10700 -6700 12500 -6680
rect 10700 -6780 10740 -6700
rect 10820 -6780 10860 -6700
rect 10980 -6780 11020 -6700
rect 11100 -6760 12100 -6700
rect 12160 -6760 12420 -6700
rect 12480 -6760 12500 -6700
rect 11100 -6780 12500 -6760
rect 13200 -6540 13600 -6500
rect 14300 -6520 16100 -6500
rect 13200 -6620 13220 -6540
rect 13300 -6620 13360 -6540
rect 13440 -6620 13500 -6540
rect 13580 -6620 13600 -6540
rect 13200 -6660 13600 -6620
rect 13200 -6740 13220 -6660
rect 13300 -6740 13360 -6660
rect 13440 -6740 13500 -6660
rect 13580 -6740 13600 -6660
rect 13200 -6780 13600 -6740
rect 14280 -6540 15700 -6520
rect 14280 -6600 14300 -6540
rect 14360 -6600 14620 -6540
rect 14680 -6600 15700 -6540
rect 15780 -6600 15820 -6520
rect 15940 -6600 15980 -6520
rect 16060 -6600 16100 -6520
rect 14280 -6620 16100 -6600
rect 14280 -6680 14300 -6620
rect 14360 -6680 14620 -6620
rect 14680 -6680 16100 -6620
rect 14280 -6700 16100 -6680
rect 14280 -6760 14300 -6700
rect 14360 -6760 14620 -6700
rect 14680 -6760 15700 -6700
rect 14280 -6780 15700 -6760
rect 15780 -6780 15820 -6700
rect 15940 -6780 15980 -6700
rect 16060 -6780 16100 -6700
rect 10700 -6800 12480 -6780
rect 13200 -6860 13220 -6780
rect 13300 -6860 13360 -6780
rect 13440 -6860 13500 -6780
rect 13580 -6860 13600 -6780
rect 14300 -6800 16100 -6780
rect 13200 -6900 13600 -6860
rect 13200 -6980 13220 -6900
rect 13300 -6980 13360 -6900
rect 13440 -6980 13500 -6900
rect 13580 -6980 13600 -6900
rect 13200 -7460 13600 -6980
rect 7900 -7480 11200 -7460
rect 7900 -7540 8000 -7480
rect 8060 -7540 8080 -7480
rect 8140 -7540 8160 -7480
rect 8220 -7540 8240 -7480
rect 8300 -7540 8320 -7480
rect 8380 -7540 8400 -7480
rect 8460 -7540 8480 -7480
rect 8540 -7540 8560 -7480
rect 8620 -7540 8640 -7480
rect 8700 -7540 8720 -7480
rect 8780 -7540 8800 -7480
rect 8860 -7540 8880 -7480
rect 8940 -7540 8960 -7480
rect 9060 -7540 9080 -7480
rect 9140 -7540 10880 -7480
rect 10940 -7540 10980 -7480
rect 11040 -7540 11200 -7480
rect 7900 -7560 11200 -7540
rect 7900 -7580 10880 -7560
rect 7900 -7640 8000 -7580
rect 8060 -7640 8080 -7580
rect 8140 -7640 8160 -7580
rect 8220 -7640 8240 -7580
rect 8300 -7640 8320 -7580
rect 8380 -7640 8400 -7580
rect 8460 -7640 8480 -7580
rect 8540 -7640 8560 -7580
rect 8620 -7640 8640 -7580
rect 8700 -7640 8720 -7580
rect 8780 -7640 8800 -7580
rect 8860 -7640 8880 -7580
rect 8940 -7640 8960 -7580
rect 9060 -7640 9080 -7580
rect 9140 -7620 10880 -7580
rect 10940 -7620 10980 -7560
rect 11040 -7620 11200 -7560
rect 9140 -7640 11200 -7620
rect 7900 -7740 11200 -7640
rect 7900 -7800 10880 -7740
rect 10940 -7800 10980 -7740
rect 11040 -7800 11200 -7740
rect 7900 -7820 11200 -7800
rect 7900 -7880 10880 -7820
rect 10940 -7880 10980 -7820
rect 11040 -7880 11200 -7820
rect 7900 -7900 11200 -7880
rect 11294 -7500 15434 -7460
rect 11294 -7560 11460 -7500
rect 11520 -7560 11540 -7500
rect 11600 -7560 12680 -7500
rect 12740 -7560 12760 -7500
rect 12820 -7560 13920 -7500
rect 13980 -7560 14000 -7500
rect 14060 -7560 15140 -7500
rect 15200 -7560 15220 -7500
rect 15280 -7560 15434 -7500
rect 11294 -7580 15434 -7560
rect 11294 -7640 11460 -7580
rect 11520 -7640 11540 -7580
rect 11600 -7640 12680 -7580
rect 12740 -7640 12760 -7580
rect 12820 -7640 13920 -7580
rect 13980 -7640 14000 -7580
rect 14060 -7640 15140 -7580
rect 15200 -7640 15220 -7580
rect 15280 -7640 15434 -7580
rect 11294 -7660 15434 -7640
rect 11294 -7720 11460 -7660
rect 11520 -7720 11540 -7660
rect 11600 -7720 12680 -7660
rect 12740 -7720 12760 -7660
rect 12820 -7720 13920 -7660
rect 13980 -7720 14000 -7660
rect 14060 -7720 15140 -7660
rect 15200 -7720 15220 -7660
rect 15280 -7720 15434 -7660
rect 11294 -7740 15434 -7720
rect 11294 -7800 11460 -7740
rect 11520 -7800 11540 -7740
rect 11600 -7800 12680 -7740
rect 12740 -7800 12760 -7740
rect 12820 -7800 13920 -7740
rect 13980 -7800 14000 -7740
rect 14060 -7800 15140 -7740
rect 15200 -7800 15220 -7740
rect 15280 -7800 15434 -7740
rect 11294 -7820 15434 -7800
rect 11294 -7880 11460 -7820
rect 11520 -7880 11540 -7820
rect 11600 -7880 12680 -7820
rect 12740 -7880 12760 -7820
rect 12820 -7880 13920 -7820
rect 13980 -7880 14000 -7820
rect 14060 -7880 15140 -7820
rect 15200 -7880 15220 -7820
rect 15280 -7880 15434 -7820
rect 11294 -7900 15434 -7880
rect 15560 -7480 18860 -7460
rect 15560 -7540 15720 -7480
rect 15780 -7540 15820 -7480
rect 15880 -7540 17660 -7480
rect 17720 -7540 17740 -7480
rect 17840 -7540 17860 -7480
rect 17920 -7540 17940 -7480
rect 18000 -7540 18020 -7480
rect 18080 -7540 18100 -7480
rect 18160 -7540 18180 -7480
rect 18240 -7540 18260 -7480
rect 18320 -7540 18340 -7480
rect 18400 -7540 18420 -7480
rect 18480 -7540 18500 -7480
rect 18560 -7540 18580 -7480
rect 18640 -7540 18660 -7480
rect 18720 -7540 18740 -7480
rect 18800 -7540 18860 -7480
rect 15560 -7560 18860 -7540
rect 15560 -7620 15720 -7560
rect 15780 -7620 15820 -7560
rect 15880 -7580 18860 -7560
rect 15880 -7620 17660 -7580
rect 15560 -7640 17660 -7620
rect 17720 -7640 17740 -7580
rect 17840 -7640 17860 -7580
rect 17920 -7640 17940 -7580
rect 18000 -7640 18020 -7580
rect 18080 -7640 18100 -7580
rect 18160 -7640 18180 -7580
rect 18240 -7640 18260 -7580
rect 18320 -7640 18340 -7580
rect 18400 -7640 18420 -7580
rect 18480 -7640 18500 -7580
rect 18560 -7640 18580 -7580
rect 18640 -7640 18660 -7580
rect 18720 -7640 18740 -7580
rect 18800 -7640 18860 -7580
rect 15560 -7740 18860 -7640
rect 15560 -7800 15720 -7740
rect 15780 -7800 15820 -7740
rect 15880 -7800 18860 -7740
rect 15560 -7820 18860 -7800
rect 15560 -7880 15720 -7820
rect 15780 -7880 15820 -7820
rect 15880 -7880 18860 -7820
rect 15560 -7900 18860 -7880
rect 10860 -8080 11200 -7900
rect 15560 -8080 15900 -7900
rect 10860 -8100 15900 -8080
rect 10860 -8160 10880 -8100
rect 10940 -8160 10980 -8100
rect 11040 -8160 12060 -8100
rect 12120 -8160 12160 -8100
rect 12220 -8160 13300 -8100
rect 13360 -8160 13400 -8100
rect 13460 -8160 14520 -8100
rect 14580 -8160 14620 -8100
rect 14680 -8160 15720 -8100
rect 15780 -8160 15820 -8100
rect 15880 -8160 15900 -8100
rect 10860 -8180 15900 -8160
rect 10860 -8240 10880 -8180
rect 10940 -8240 10980 -8180
rect 11040 -8240 12060 -8180
rect 12120 -8240 12160 -8180
rect 12220 -8240 13300 -8180
rect 13360 -8240 13400 -8180
rect 13460 -8240 14520 -8180
rect 14580 -8240 14620 -8180
rect 14680 -8240 15720 -8180
rect 15780 -8240 15820 -8180
rect 15880 -8240 15900 -8180
rect 10860 -8320 15900 -8240
rect 10860 -8380 10880 -8320
rect 10940 -8380 10980 -8320
rect 11040 -8380 12060 -8320
rect 12120 -8380 12160 -8320
rect 12220 -8380 13300 -8320
rect 13360 -8380 13400 -8320
rect 13460 -8380 14520 -8320
rect 14580 -8380 14620 -8320
rect 14680 -8380 15720 -8320
rect 15780 -8380 15820 -8320
rect 15880 -8380 15900 -8320
rect 10860 -8400 15900 -8380
rect 10860 -8460 10880 -8400
rect 10940 -8460 10980 -8400
rect 11040 -8460 12060 -8400
rect 12120 -8460 12160 -8400
rect 12220 -8460 13300 -8400
rect 13360 -8460 13400 -8400
rect 13460 -8460 14520 -8400
rect 14580 -8460 14620 -8400
rect 14680 -8460 15720 -8400
rect 15780 -8460 15820 -8400
rect 15880 -8460 15900 -8400
rect 10860 -8480 15900 -8460
rect 9300 -10020 9700 -10000
rect 9300 -10100 9320 -10020
rect 9400 -10100 9460 -10020
rect 9540 -10100 9600 -10020
rect 9680 -10100 9700 -10020
rect 9300 -10160 9700 -10100
rect 9300 -10240 9320 -10160
rect 9400 -10240 9460 -10160
rect 9540 -10240 9600 -10160
rect 9680 -10240 9700 -10160
rect 9300 -10300 9700 -10240
rect 9300 -10380 9320 -10300
rect 9400 -10380 9460 -10300
rect 9540 -10380 9600 -10300
rect 9680 -10380 9700 -10300
rect 9300 -10400 9700 -10380
rect 13200 -10620 13600 -8480
rect 17100 -10020 17500 -10000
rect 17100 -10100 17120 -10020
rect 17200 -10100 17260 -10020
rect 17340 -10100 17400 -10020
rect 17480 -10100 17500 -10020
rect 17100 -10160 17500 -10100
rect 17100 -10240 17120 -10160
rect 17200 -10240 17260 -10160
rect 17340 -10240 17400 -10160
rect 17480 -10240 17500 -10160
rect 17100 -10300 17500 -10240
rect 17100 -10380 17120 -10300
rect 17200 -10380 17260 -10300
rect 17340 -10380 17400 -10300
rect 17480 -10380 17500 -10300
rect 17100 -10400 17500 -10380
rect 13200 -10680 13220 -10620
rect 13280 -10680 13320 -10620
rect 13380 -10680 13420 -10620
rect 13480 -10680 13520 -10620
rect 13580 -10680 13600 -10620
rect 13200 -10720 13600 -10680
rect 13200 -10780 13220 -10720
rect 13280 -10780 13320 -10720
rect 13380 -10780 13420 -10720
rect 13480 -10780 13520 -10720
rect 13580 -10780 13600 -10720
rect 13200 -10820 13600 -10780
rect 13200 -10880 13220 -10820
rect 13280 -10880 13320 -10820
rect 13380 -10880 13420 -10820
rect 13480 -10880 13520 -10820
rect 13580 -10880 13600 -10820
rect 13200 -10920 13600 -10880
rect 13200 -10980 13220 -10920
rect 13280 -10980 13320 -10920
rect 13380 -10980 13420 -10920
rect 13480 -10980 13520 -10920
rect 13580 -10980 13600 -10920
rect 8240 -11420 8640 -11400
rect 8240 -11480 8260 -11420
rect 8320 -11480 8360 -11420
rect 8420 -11480 8460 -11420
rect 8520 -11480 8560 -11420
rect 8620 -11480 8640 -11420
rect 8240 -11500 8640 -11480
rect 8240 -11560 8260 -11500
rect 8320 -11560 8360 -11500
rect 8420 -11560 8460 -11500
rect 8520 -11560 8560 -11500
rect 8620 -11560 8640 -11500
rect 8240 -11600 8640 -11560
rect 8240 -11660 8260 -11600
rect 8320 -11660 8360 -11600
rect 8420 -11660 8460 -11600
rect 8520 -11660 8560 -11600
rect 8620 -11660 8640 -11600
rect 8240 -11700 8640 -11660
rect 8240 -11760 8260 -11700
rect 8320 -11760 8360 -11700
rect 8420 -11760 8460 -11700
rect 8520 -11760 8560 -11700
rect 8620 -11760 8640 -11700
rect 8240 -11780 8640 -11760
rect 18160 -11420 18560 -11400
rect 18160 -11480 18180 -11420
rect 18240 -11480 18280 -11420
rect 18340 -11480 18380 -11420
rect 18440 -11480 18480 -11420
rect 18540 -11480 18560 -11420
rect 18160 -11500 18560 -11480
rect 18160 -11560 18180 -11500
rect 18240 -11560 18280 -11500
rect 18340 -11560 18380 -11500
rect 18440 -11560 18480 -11500
rect 18540 -11560 18560 -11500
rect 18160 -11600 18560 -11560
rect 18160 -11660 18180 -11600
rect 18240 -11660 18280 -11600
rect 18340 -11660 18380 -11600
rect 18440 -11660 18480 -11600
rect 18540 -11660 18560 -11600
rect 18160 -11700 18560 -11660
rect 18160 -11760 18180 -11700
rect 18240 -11760 18280 -11700
rect 18340 -11760 18380 -11700
rect 18440 -11760 18480 -11700
rect 18540 -11760 18560 -11700
rect 18160 -11780 18560 -11760
<< via2 >>
rect 13220 -2060 13300 -1980
rect 13360 -2060 13440 -1980
rect 13500 -2060 13580 -1980
rect 13220 -2180 13300 -2100
rect 13360 -2180 13440 -2100
rect 13500 -2180 13580 -2100
rect 13220 -2320 13300 -2240
rect 13360 -2320 13440 -2240
rect 13500 -2320 13580 -2240
rect 8280 -2940 8340 -2880
rect 8400 -2940 8480 -2880
rect 8540 -2940 8600 -2880
rect 8280 -3120 8340 -3060
rect 8400 -3120 8480 -3060
rect 8540 -3120 8600 -3060
rect 10740 -3020 10820 -2940
rect 10880 -3020 10960 -2940
rect 11020 -3020 11100 -2940
rect 15700 -3020 15780 -2940
rect 15840 -3020 15920 -2940
rect 15980 -3020 16060 -2940
rect 10740 -3160 10820 -3080
rect 10880 -3160 10960 -3080
rect 11020 -3160 11100 -3080
rect 15700 -3160 15780 -3080
rect 15840 -3160 15920 -3080
rect 15980 -3160 16060 -3080
rect 18200 -2940 18260 -2880
rect 18320 -2940 18400 -2880
rect 18460 -2940 18520 -2880
rect 18200 -3120 18260 -3060
rect 18320 -3120 18400 -3060
rect 18460 -3120 18520 -3060
rect 10740 -3300 10820 -3220
rect 10880 -3300 10960 -3220
rect 11020 -3300 11100 -3220
rect 15700 -3300 15780 -3220
rect 15840 -3300 15920 -3220
rect 15980 -3300 16060 -3220
rect 10020 -3480 10080 -3420
rect 10120 -3480 10180 -3420
rect 10260 -3480 10340 -3420
rect 10420 -3480 10480 -3420
rect 10520 -3480 10580 -3420
rect 11720 -3500 11800 -3420
rect 11860 -3500 11940 -3420
rect 12000 -3500 12080 -3420
rect 13220 -3500 13300 -3420
rect 13360 -3500 13440 -3420
rect 13500 -3500 13580 -3420
rect 14720 -3500 14800 -3420
rect 14860 -3500 14940 -3420
rect 15000 -3500 15080 -3420
rect 16220 -3480 16280 -3420
rect 16320 -3480 16380 -3420
rect 16460 -3480 16540 -3420
rect 16620 -3480 16680 -3420
rect 16720 -3480 16780 -3420
rect 10020 -3640 10100 -3560
rect 10140 -3640 10200 -3560
rect 10260 -3640 10340 -3560
rect 10400 -3640 10460 -3560
rect 10500 -3640 10580 -3560
rect 11720 -3640 11800 -3560
rect 11860 -3640 11940 -3560
rect 12000 -3640 12080 -3560
rect 13220 -3640 13300 -3560
rect 13360 -3640 13440 -3560
rect 13500 -3640 13580 -3560
rect 14720 -3640 14800 -3560
rect 14860 -3640 14940 -3560
rect 15000 -3640 15080 -3560
rect 16220 -3640 16300 -3560
rect 16340 -3640 16400 -3560
rect 16460 -3640 16540 -3560
rect 16600 -3640 16660 -3560
rect 16700 -3640 16780 -3560
rect 10020 -3780 10080 -3720
rect 10120 -3780 10180 -3720
rect 10260 -3780 10340 -3720
rect 10420 -3780 10480 -3720
rect 10520 -3780 10580 -3720
rect 11720 -3780 11800 -3700
rect 11860 -3780 11940 -3700
rect 12000 -3780 12080 -3700
rect 13220 -3780 13300 -3700
rect 13360 -3780 13440 -3700
rect 13500 -3780 13580 -3700
rect 14720 -3780 14800 -3700
rect 14860 -3780 14940 -3700
rect 15000 -3780 15080 -3700
rect 16220 -3780 16280 -3720
rect 16320 -3780 16380 -3720
rect 16460 -3780 16540 -3720
rect 16620 -3780 16680 -3720
rect 16720 -3780 16780 -3720
rect 7220 -4100 7300 -4040
rect 7340 -4080 7400 -4020
rect 7460 -4100 7540 -4040
rect 7600 -4080 7660 -4020
rect 7700 -4100 7780 -4040
rect 7220 -4200 7300 -4140
rect 7340 -4200 7400 -4140
rect 7460 -4200 7540 -4140
rect 7600 -4200 7660 -4140
rect 7700 -4200 7780 -4140
rect 19020 -4100 19100 -4040
rect 19140 -4080 19200 -4020
rect 19260 -4100 19340 -4040
rect 19400 -4080 19460 -4020
rect 19500 -4100 19580 -4040
rect 19020 -4200 19100 -4140
rect 19140 -4200 19200 -4140
rect 19260 -4200 19340 -4140
rect 19400 -4200 19460 -4140
rect 19500 -4200 19580 -4140
rect 8420 -4500 8480 -4440
rect 8520 -4500 8580 -4440
rect 8420 -4600 8480 -4540
rect 8520 -4600 8580 -4540
rect 10740 -4500 10820 -4420
rect 10860 -4500 10960 -4420
rect 11000 -4500 11080 -4420
rect 10740 -4680 10820 -4600
rect 10860 -4680 10960 -4600
rect 11000 -4680 11080 -4600
rect 11720 -4500 11800 -4420
rect 11840 -4500 11960 -4420
rect 12000 -4500 12080 -4420
rect 11720 -4680 11800 -4600
rect 11840 -4680 11960 -4600
rect 12000 -4680 12080 -4600
rect 14720 -4500 14800 -4420
rect 14840 -4500 14960 -4420
rect 15000 -4500 15080 -4420
rect 14720 -4680 14800 -4600
rect 14840 -4680 14960 -4600
rect 15000 -4680 15080 -4600
rect 15720 -4500 15800 -4420
rect 15840 -4500 15940 -4420
rect 15980 -4500 16060 -4420
rect 15720 -4680 15800 -4600
rect 15840 -4680 15940 -4600
rect 15980 -4680 16060 -4600
rect 18260 -4500 18320 -4440
rect 18360 -4500 18420 -4440
rect 18260 -4600 18320 -4540
rect 18360 -4600 18420 -4540
rect 12940 -5060 13080 -4920
rect 9320 -5180 9400 -5100
rect 9440 -5180 9520 -5100
rect 9560 -5180 9640 -5100
rect 9320 -5280 9380 -5220
rect 9440 -5280 9520 -5220
rect 9580 -5280 9640 -5220
rect 11440 -5180 11500 -5120
rect 11540 -5180 11600 -5120
rect 11200 -5320 11260 -5260
rect 9320 -5400 9400 -5320
rect 9440 -5400 9520 -5320
rect 9560 -5400 9640 -5320
rect 11280 -5400 11340 -5340
rect 13720 -5060 13860 -4920
rect 15200 -5180 15260 -5120
rect 15300 -5180 15360 -5120
rect 15540 -5320 15600 -5260
rect 15460 -5400 15520 -5340
rect 11540 -5560 11600 -5500
rect 11460 -5640 11520 -5580
rect 11200 -5780 11260 -5720
rect 11300 -5780 11360 -5720
rect 8280 -6020 8340 -5960
rect 8400 -6020 8460 -5960
rect 8280 -6200 8340 -6140
rect 8400 -6200 8460 -6140
rect 11720 -6000 11800 -5920
rect 11840 -6000 11960 -5920
rect 12000 -6000 12080 -5920
rect 12940 -5980 13080 -5840
rect 11720 -6180 11800 -6100
rect 11840 -6180 11960 -6100
rect 12000 -6180 12080 -6100
rect 15200 -5560 15260 -5500
rect 17160 -5580 17240 -5500
rect 17280 -5580 17360 -5500
rect 17400 -5580 17480 -5500
rect 15280 -5640 15340 -5580
rect 15440 -5780 15500 -5720
rect 15540 -5780 15600 -5720
rect 17160 -5680 17240 -5620
rect 17280 -5680 17360 -5620
rect 17400 -5680 17480 -5620
rect 17160 -5800 17240 -5720
rect 17280 -5800 17360 -5720
rect 17400 -5800 17480 -5720
rect 13720 -5980 13860 -5840
rect 14720 -6000 14800 -5920
rect 14840 -6000 14960 -5920
rect 15000 -6000 15080 -5920
rect 14720 -6180 14800 -6100
rect 14840 -6180 14960 -6100
rect 15000 -6180 15080 -6100
rect 18340 -6020 18400 -5960
rect 18460 -6020 18520 -5960
rect 18340 -6200 18400 -6140
rect 18460 -6200 18520 -6140
rect 10740 -6600 10820 -6520
rect 10860 -6600 10980 -6520
rect 11020 -6600 11100 -6520
rect 10740 -6780 10820 -6700
rect 10860 -6780 10980 -6700
rect 11020 -6780 11100 -6700
rect 15700 -6600 15780 -6520
rect 15820 -6600 15940 -6520
rect 15980 -6600 16060 -6520
rect 15700 -6780 15780 -6700
rect 15820 -6780 15940 -6700
rect 15980 -6780 16060 -6700
rect 9320 -10100 9400 -10020
rect 9460 -10100 9540 -10020
rect 9600 -10100 9680 -10020
rect 9320 -10240 9400 -10160
rect 9460 -10240 9540 -10160
rect 9600 -10240 9680 -10160
rect 9320 -10380 9400 -10300
rect 9460 -10380 9540 -10300
rect 9600 -10380 9680 -10300
rect 17120 -10100 17200 -10020
rect 17260 -10100 17340 -10020
rect 17400 -10100 17480 -10020
rect 17120 -10240 17200 -10160
rect 17260 -10240 17340 -10160
rect 17400 -10240 17480 -10160
rect 17120 -10380 17200 -10300
rect 17260 -10380 17340 -10300
rect 17400 -10380 17480 -10300
rect 8260 -11480 8320 -11420
rect 8360 -11480 8420 -11420
rect 8460 -11480 8520 -11420
rect 8560 -11480 8620 -11420
rect 8260 -11760 8320 -11700
rect 8360 -11760 8420 -11700
rect 8460 -11760 8520 -11700
rect 8560 -11760 8620 -11700
rect 18180 -11480 18240 -11420
rect 18280 -11480 18340 -11420
rect 18380 -11480 18440 -11420
rect 18480 -11480 18540 -11420
rect 18180 -11760 18240 -11700
rect 18280 -11760 18340 -11700
rect 18380 -11760 18440 -11700
rect 18480 -11760 18540 -11700
<< metal3 >>
rect 13200 -1980 13600 -1960
rect 13200 -2060 13220 -1980
rect 13300 -2060 13360 -1980
rect 13440 -2060 13500 -1980
rect 13580 -2060 13600 -1980
rect 13200 -2100 13600 -2060
rect 13200 -2180 13220 -2100
rect 13300 -2180 13360 -2100
rect 13440 -2180 13500 -2100
rect 13580 -2180 13600 -2100
rect 13200 -2240 13600 -2180
rect 13200 -2320 13220 -2240
rect 13300 -2320 13360 -2240
rect 13440 -2320 13500 -2240
rect 13580 -2320 13600 -2240
rect 8240 -2880 8640 -2860
rect 8240 -2940 8280 -2880
rect 8340 -2940 8400 -2880
rect 8480 -2940 8540 -2880
rect 8600 -2940 8640 -2880
rect 8240 -3060 8640 -2940
rect 8240 -3120 8280 -3060
rect 8340 -3120 8400 -3060
rect 8480 -3120 8540 -3060
rect 8600 -3120 8640 -3060
rect 7200 -4020 7800 -4000
rect 7200 -4100 7220 -4020
rect 7300 -4100 7320 -4020
rect 7400 -4100 7460 -4020
rect 7540 -4100 7600 -4020
rect 7680 -4100 7700 -4020
rect 7780 -4100 7800 -4020
rect 7200 -4140 7800 -4100
rect 7200 -4220 7220 -4140
rect 7300 -4220 7320 -4140
rect 7400 -4220 7460 -4140
rect 7540 -4220 7600 -4140
rect 7680 -4220 7700 -4140
rect 7780 -4220 7800 -4140
rect 8240 -4440 8640 -3120
rect 10720 -2940 11120 -2920
rect 10720 -3020 10740 -2940
rect 10820 -3020 10880 -2940
rect 10960 -3020 11020 -2940
rect 11100 -3020 11120 -2940
rect 10720 -3080 11120 -3020
rect 10720 -3160 10740 -3080
rect 10820 -3160 10880 -3080
rect 10960 -3160 11020 -3080
rect 11100 -3160 11120 -3080
rect 10720 -3220 11120 -3160
rect 10720 -3300 10740 -3220
rect 10820 -3300 10880 -3220
rect 10960 -3300 11020 -3220
rect 11100 -3300 11120 -3220
rect 10000 -3420 10600 -3400
rect 10000 -3500 10020 -3420
rect 10100 -3500 10120 -3420
rect 10200 -3500 10260 -3420
rect 10340 -3500 10400 -3420
rect 10480 -3500 10500 -3420
rect 10580 -3500 10600 -3420
rect 10000 -3560 10600 -3500
rect 10000 -3640 10020 -3560
rect 10100 -3640 10120 -3560
rect 10200 -3640 10260 -3560
rect 10340 -3640 10400 -3560
rect 10480 -3640 10500 -3560
rect 10580 -3640 10600 -3560
rect 10000 -3700 10600 -3640
rect 10000 -3780 10020 -3700
rect 10100 -3780 10120 -3700
rect 10200 -3780 10260 -3700
rect 10340 -3780 10400 -3700
rect 10480 -3780 10500 -3700
rect 10580 -3780 10600 -3700
rect 10000 -3800 10600 -3780
rect 8240 -4500 8420 -4440
rect 8480 -4500 8520 -4440
rect 8580 -4500 8640 -4440
rect 8240 -4540 8640 -4500
rect 8240 -4600 8420 -4540
rect 8480 -4600 8520 -4540
rect 8580 -4600 8640 -4540
rect 8240 -5960 8640 -4600
rect 10720 -4420 11120 -3300
rect 10720 -4500 10740 -4420
rect 10820 -4500 10860 -4420
rect 10960 -4500 11000 -4420
rect 11080 -4500 11120 -4420
rect 10720 -4600 11120 -4500
rect 10720 -4680 10740 -4600
rect 10820 -4680 10860 -4600
rect 10960 -4680 11000 -4600
rect 11080 -4680 11120 -4600
rect 8240 -6020 8280 -5960
rect 8340 -6020 8400 -5960
rect 8460 -6020 8640 -5960
rect 8240 -6140 8640 -6020
rect 8240 -6200 8280 -6140
rect 8340 -6200 8400 -6140
rect 8460 -6200 8640 -6140
rect 8240 -11400 8640 -6200
rect 9300 -5100 9660 -5080
rect 9300 -5180 9320 -5100
rect 9400 -5180 9440 -5100
rect 9520 -5180 9560 -5100
rect 9640 -5180 9660 -5100
rect 9300 -5220 9660 -5180
rect 9300 -5280 9320 -5220
rect 9380 -5280 9440 -5220
rect 9520 -5280 9580 -5220
rect 9640 -5240 9660 -5220
rect 9640 -5280 9700 -5240
rect 9300 -5320 9700 -5280
rect 9300 -5400 9320 -5320
rect 9400 -5400 9440 -5320
rect 9520 -5400 9560 -5320
rect 9640 -5400 9700 -5320
rect 9300 -10020 9700 -5400
rect 10720 -6520 11120 -4680
rect 11700 -3420 12100 -3400
rect 11700 -3500 11720 -3420
rect 11800 -3500 11860 -3420
rect 11940 -3500 12000 -3420
rect 12080 -3500 12100 -3420
rect 11700 -3560 12100 -3500
rect 11700 -3640 11720 -3560
rect 11800 -3640 11860 -3560
rect 11940 -3640 12000 -3560
rect 12080 -3640 12100 -3560
rect 11700 -3700 12100 -3640
rect 11700 -3780 11720 -3700
rect 11800 -3780 11860 -3700
rect 11940 -3780 12000 -3700
rect 12080 -3780 12100 -3700
rect 11700 -4420 12100 -3780
rect 13200 -3420 13600 -2320
rect 18160 -2880 18560 -2860
rect 15680 -2940 16080 -2920
rect 15680 -3020 15700 -2940
rect 15780 -3020 15840 -2940
rect 15920 -3020 15980 -2940
rect 16060 -3020 16080 -2940
rect 15680 -3080 16080 -3020
rect 15680 -3160 15700 -3080
rect 15780 -3160 15840 -3080
rect 15920 -3160 15980 -3080
rect 16060 -3160 16080 -3080
rect 15680 -3220 16080 -3160
rect 15680 -3300 15700 -3220
rect 15780 -3300 15840 -3220
rect 15920 -3300 15980 -3220
rect 16060 -3300 16080 -3220
rect 13200 -3500 13220 -3420
rect 13300 -3500 13360 -3420
rect 13440 -3500 13500 -3420
rect 13580 -3500 13600 -3420
rect 13200 -3560 13600 -3500
rect 13200 -3640 13220 -3560
rect 13300 -3640 13360 -3560
rect 13440 -3640 13500 -3560
rect 13580 -3640 13600 -3560
rect 13200 -3700 13600 -3640
rect 13200 -3780 13220 -3700
rect 13300 -3780 13360 -3700
rect 13440 -3780 13500 -3700
rect 13580 -3780 13600 -3700
rect 13200 -3800 13600 -3780
rect 14700 -3420 15100 -3400
rect 14700 -3500 14720 -3420
rect 14800 -3500 14860 -3420
rect 14940 -3500 15000 -3420
rect 15080 -3500 15100 -3420
rect 14700 -3560 15100 -3500
rect 14700 -3640 14720 -3560
rect 14800 -3640 14860 -3560
rect 14940 -3640 15000 -3560
rect 15080 -3640 15100 -3560
rect 14700 -3700 15100 -3640
rect 14700 -3780 14720 -3700
rect 14800 -3780 14860 -3700
rect 14940 -3780 15000 -3700
rect 15080 -3780 15100 -3700
rect 11700 -4500 11720 -4420
rect 11800 -4500 11840 -4420
rect 11960 -4500 12000 -4420
rect 12080 -4500 12100 -4420
rect 11700 -4600 12100 -4500
rect 11700 -4680 11720 -4600
rect 11800 -4680 11840 -4600
rect 11960 -4680 12000 -4600
rect 12080 -4680 12100 -4600
rect 11420 -5120 11620 -5100
rect 11420 -5180 11440 -5120
rect 11500 -5180 11540 -5120
rect 11600 -5180 11620 -5120
rect 11420 -5200 11620 -5180
rect 11180 -5260 11360 -5240
rect 11180 -5320 11200 -5260
rect 11260 -5320 11360 -5260
rect 11180 -5340 11360 -5320
rect 11180 -5400 11280 -5340
rect 11340 -5400 11360 -5340
rect 11180 -5700 11360 -5400
rect 11440 -5500 11620 -5200
rect 11440 -5560 11540 -5500
rect 11600 -5560 11620 -5500
rect 11440 -5580 11620 -5560
rect 11440 -5640 11460 -5580
rect 11520 -5640 11620 -5580
rect 11440 -5660 11620 -5640
rect 11180 -5720 11380 -5700
rect 11180 -5780 11200 -5720
rect 11260 -5780 11300 -5720
rect 11360 -5780 11380 -5720
rect 11180 -5800 11380 -5780
rect 10720 -6600 10740 -6520
rect 10820 -6600 10860 -6520
rect 10980 -6600 11020 -6520
rect 11100 -6600 11120 -6520
rect 10720 -6700 11120 -6600
rect 10720 -6780 10740 -6700
rect 10820 -6780 10860 -6700
rect 10980 -6780 11020 -6700
rect 11100 -6780 11120 -6700
rect 10720 -7100 11120 -6780
rect 11700 -5920 12100 -4680
rect 14700 -4420 15100 -3780
rect 14700 -4500 14720 -4420
rect 14800 -4500 14840 -4420
rect 14960 -4500 15000 -4420
rect 15080 -4500 15100 -4420
rect 14700 -4600 15100 -4500
rect 14700 -4680 14720 -4600
rect 14800 -4680 14840 -4600
rect 14960 -4680 15000 -4600
rect 15080 -4680 15100 -4600
rect 12920 -4920 13880 -4900
rect 12920 -5060 12940 -4920
rect 13080 -5060 13720 -4920
rect 13860 -5060 13880 -4920
rect 12920 -5080 13880 -5060
rect 11700 -6000 11720 -5920
rect 11800 -6000 11840 -5920
rect 11960 -6000 12000 -5920
rect 12080 -6000 12100 -5920
rect 12920 -5840 13880 -5820
rect 12920 -5980 12940 -5840
rect 13080 -5980 13720 -5840
rect 13860 -5980 13880 -5840
rect 12920 -6000 13880 -5980
rect 14700 -5920 15100 -4680
rect 15680 -4420 16080 -3300
rect 18160 -2940 18200 -2880
rect 18260 -2940 18320 -2880
rect 18400 -2940 18460 -2880
rect 18520 -2940 18560 -2880
rect 18160 -3060 18560 -2940
rect 18160 -3120 18200 -3060
rect 18260 -3120 18320 -3060
rect 18400 -3120 18460 -3060
rect 18520 -3120 18560 -3060
rect 16200 -3420 16800 -3400
rect 16200 -3500 16220 -3420
rect 16300 -3500 16320 -3420
rect 16400 -3500 16460 -3420
rect 16540 -3500 16600 -3420
rect 16680 -3500 16700 -3420
rect 16780 -3500 16800 -3420
rect 16200 -3560 16800 -3500
rect 16200 -3640 16220 -3560
rect 16300 -3640 16320 -3560
rect 16400 -3640 16460 -3560
rect 16540 -3640 16600 -3560
rect 16680 -3640 16700 -3560
rect 16780 -3640 16800 -3560
rect 16200 -3700 16800 -3640
rect 16200 -3780 16220 -3700
rect 16300 -3780 16320 -3700
rect 16400 -3780 16460 -3700
rect 16540 -3780 16600 -3700
rect 16680 -3780 16700 -3700
rect 16780 -3780 16800 -3700
rect 16200 -3800 16800 -3780
rect 15680 -4500 15720 -4420
rect 15800 -4500 15840 -4420
rect 15940 -4500 15980 -4420
rect 16060 -4500 16080 -4420
rect 15680 -4600 16080 -4500
rect 15680 -4680 15720 -4600
rect 15800 -4680 15840 -4600
rect 15940 -4680 15980 -4600
rect 16060 -4680 16080 -4600
rect 15180 -5120 15380 -5100
rect 15180 -5180 15200 -5120
rect 15260 -5180 15300 -5120
rect 15360 -5180 15380 -5120
rect 15180 -5200 15380 -5180
rect 15180 -5500 15360 -5200
rect 15180 -5560 15200 -5500
rect 15260 -5560 15360 -5500
rect 15180 -5580 15360 -5560
rect 15180 -5640 15280 -5580
rect 15340 -5640 15360 -5580
rect 15180 -5660 15360 -5640
rect 15440 -5260 15620 -5240
rect 15440 -5320 15540 -5260
rect 15600 -5320 15620 -5260
rect 15440 -5340 15620 -5320
rect 15440 -5400 15460 -5340
rect 15520 -5400 15620 -5340
rect 15440 -5700 15620 -5400
rect 15420 -5720 15620 -5700
rect 15420 -5780 15440 -5720
rect 15500 -5780 15540 -5720
rect 15600 -5780 15620 -5720
rect 15420 -5800 15620 -5780
rect 14700 -6000 14720 -5920
rect 14800 -6000 14840 -5920
rect 14960 -6000 15000 -5920
rect 15080 -6000 15100 -5920
rect 11700 -6100 12100 -6000
rect 11700 -6180 11720 -6100
rect 11800 -6180 11840 -6100
rect 11960 -6180 12000 -6100
rect 12080 -6180 12100 -6100
rect 11700 -7100 12100 -6180
rect 14700 -6100 15100 -6000
rect 14700 -6180 14720 -6100
rect 14800 -6180 14840 -6100
rect 14960 -6180 15000 -6100
rect 15080 -6180 15100 -6100
rect 14700 -7100 15100 -6180
rect 15680 -6520 16080 -4680
rect 18160 -4440 18560 -3120
rect 19000 -4020 19600 -4000
rect 19000 -4100 19020 -4020
rect 19100 -4100 19120 -4020
rect 19200 -4100 19260 -4020
rect 19340 -4100 19400 -4020
rect 19480 -4100 19500 -4020
rect 19580 -4100 19600 -4020
rect 19000 -4140 19600 -4100
rect 19000 -4220 19020 -4140
rect 19100 -4220 19120 -4140
rect 19200 -4220 19260 -4140
rect 19340 -4220 19400 -4140
rect 19480 -4220 19500 -4140
rect 19580 -4220 19600 -4140
rect 18160 -4500 18260 -4440
rect 18320 -4500 18360 -4440
rect 18420 -4500 18560 -4440
rect 18160 -4540 18560 -4500
rect 18160 -4600 18260 -4540
rect 18320 -4600 18360 -4540
rect 18420 -4600 18560 -4540
rect 17140 -5240 17500 -5080
rect 15680 -6600 15700 -6520
rect 15780 -6600 15820 -6520
rect 15940 -6600 15980 -6520
rect 16060 -6600 16080 -6520
rect 15680 -6700 16080 -6600
rect 15680 -6780 15700 -6700
rect 15780 -6780 15820 -6700
rect 15940 -6780 15980 -6700
rect 16060 -6780 16080 -6700
rect 15680 -7100 16080 -6780
rect 17100 -5500 17500 -5240
rect 17100 -5580 17160 -5500
rect 17240 -5580 17280 -5500
rect 17360 -5580 17400 -5500
rect 17480 -5580 17500 -5500
rect 17100 -5620 17500 -5580
rect 17100 -5680 17160 -5620
rect 17240 -5680 17280 -5620
rect 17360 -5680 17400 -5620
rect 17480 -5680 17500 -5620
rect 17100 -5720 17500 -5680
rect 17100 -5800 17160 -5720
rect 17240 -5800 17280 -5720
rect 17360 -5800 17400 -5720
rect 17480 -5800 17500 -5720
rect 9300 -10100 9320 -10020
rect 9400 -10100 9460 -10020
rect 9540 -10100 9600 -10020
rect 9680 -10100 9700 -10020
rect 9300 -10160 9700 -10100
rect 9300 -10240 9320 -10160
rect 9400 -10240 9460 -10160
rect 9540 -10240 9600 -10160
rect 9680 -10240 9700 -10160
rect 9300 -10300 9700 -10240
rect 9300 -10380 9320 -10300
rect 9400 -10380 9460 -10300
rect 9540 -10380 9600 -10300
rect 9680 -10380 9700 -10300
rect 9300 -10400 9700 -10380
rect 17100 -10020 17500 -5800
rect 17100 -10100 17120 -10020
rect 17200 -10100 17260 -10020
rect 17340 -10100 17400 -10020
rect 17480 -10100 17500 -10020
rect 17100 -10160 17500 -10100
rect 17100 -10240 17120 -10160
rect 17200 -10240 17260 -10160
rect 17340 -10240 17400 -10160
rect 17480 -10240 17500 -10160
rect 17100 -10300 17500 -10240
rect 17100 -10380 17120 -10300
rect 17200 -10380 17260 -10300
rect 17340 -10380 17400 -10300
rect 17480 -10380 17500 -10300
rect 17100 -10400 17500 -10380
rect 18160 -5960 18560 -4600
rect 18160 -6020 18340 -5960
rect 18400 -6020 18460 -5960
rect 18520 -6020 18560 -5960
rect 18160 -6140 18560 -6020
rect 18160 -6200 18340 -6140
rect 18400 -6200 18460 -6140
rect 18520 -6200 18560 -6140
rect 18160 -11400 18560 -6200
rect 8240 -11420 18560 -11400
rect 8240 -11480 8260 -11420
rect 8320 -11480 8360 -11420
rect 8420 -11480 8460 -11420
rect 8520 -11480 8560 -11420
rect 8620 -11480 18180 -11420
rect 18240 -11480 18280 -11420
rect 18340 -11480 18380 -11420
rect 18440 -11480 18480 -11420
rect 18540 -11480 18560 -11420
rect 8240 -11700 18560 -11480
rect 8240 -11760 8260 -11700
rect 8320 -11760 8360 -11700
rect 8420 -11760 8460 -11700
rect 8520 -11760 8560 -11700
rect 8620 -11760 18180 -11700
rect 18240 -11760 18280 -11700
rect 18340 -11760 18380 -11700
rect 18440 -11760 18480 -11700
rect 18540 -11760 18560 -11700
rect 8240 -11780 18560 -11760
<< via3 >>
rect 7220 -4040 7300 -4020
rect 7220 -4100 7300 -4040
rect 7320 -4080 7340 -4020
rect 7340 -4080 7400 -4020
rect 7320 -4100 7400 -4080
rect 7460 -4040 7540 -4020
rect 7460 -4100 7540 -4040
rect 7600 -4080 7660 -4020
rect 7660 -4080 7680 -4020
rect 7600 -4100 7680 -4080
rect 7700 -4040 7780 -4020
rect 7700 -4100 7780 -4040
rect 7220 -4200 7300 -4140
rect 7220 -4220 7300 -4200
rect 7320 -4200 7340 -4140
rect 7340 -4200 7400 -4140
rect 7320 -4220 7400 -4200
rect 7460 -4200 7540 -4140
rect 7460 -4220 7540 -4200
rect 7600 -4200 7660 -4140
rect 7660 -4200 7680 -4140
rect 7600 -4220 7680 -4200
rect 7700 -4200 7780 -4140
rect 7700 -4220 7780 -4200
rect 10020 -3480 10080 -3420
rect 10080 -3480 10100 -3420
rect 10020 -3500 10100 -3480
rect 10120 -3480 10180 -3420
rect 10180 -3480 10200 -3420
rect 10120 -3500 10200 -3480
rect 10260 -3480 10340 -3420
rect 10260 -3500 10340 -3480
rect 10400 -3480 10420 -3420
rect 10420 -3480 10480 -3420
rect 10400 -3500 10480 -3480
rect 10500 -3480 10520 -3420
rect 10520 -3480 10580 -3420
rect 10500 -3500 10580 -3480
rect 10020 -3640 10100 -3560
rect 10120 -3640 10140 -3560
rect 10140 -3640 10200 -3560
rect 10260 -3640 10340 -3560
rect 10400 -3640 10460 -3560
rect 10460 -3640 10480 -3560
rect 10500 -3640 10580 -3560
rect 10020 -3720 10100 -3700
rect 10020 -3780 10080 -3720
rect 10080 -3780 10100 -3720
rect 10120 -3720 10200 -3700
rect 10120 -3780 10180 -3720
rect 10180 -3780 10200 -3720
rect 10260 -3720 10340 -3700
rect 10260 -3780 10340 -3720
rect 10400 -3720 10480 -3700
rect 10400 -3780 10420 -3720
rect 10420 -3780 10480 -3720
rect 10500 -3720 10580 -3700
rect 10500 -3780 10520 -3720
rect 10520 -3780 10580 -3720
rect 16220 -3480 16280 -3420
rect 16280 -3480 16300 -3420
rect 16220 -3500 16300 -3480
rect 16320 -3480 16380 -3420
rect 16380 -3480 16400 -3420
rect 16320 -3500 16400 -3480
rect 16460 -3480 16540 -3420
rect 16460 -3500 16540 -3480
rect 16600 -3480 16620 -3420
rect 16620 -3480 16680 -3420
rect 16600 -3500 16680 -3480
rect 16700 -3480 16720 -3420
rect 16720 -3480 16780 -3420
rect 16700 -3500 16780 -3480
rect 16220 -3640 16300 -3560
rect 16320 -3640 16340 -3560
rect 16340 -3640 16400 -3560
rect 16460 -3640 16540 -3560
rect 16600 -3640 16660 -3560
rect 16660 -3640 16680 -3560
rect 16700 -3640 16780 -3560
rect 16220 -3720 16300 -3700
rect 16220 -3780 16280 -3720
rect 16280 -3780 16300 -3720
rect 16320 -3720 16400 -3700
rect 16320 -3780 16380 -3720
rect 16380 -3780 16400 -3720
rect 16460 -3720 16540 -3700
rect 16460 -3780 16540 -3720
rect 16600 -3720 16680 -3700
rect 16600 -3780 16620 -3720
rect 16620 -3780 16680 -3720
rect 16700 -3720 16780 -3700
rect 16700 -3780 16720 -3720
rect 16720 -3780 16780 -3720
rect 19020 -4040 19100 -4020
rect 19020 -4100 19100 -4040
rect 19120 -4080 19140 -4020
rect 19140 -4080 19200 -4020
rect 19120 -4100 19200 -4080
rect 19260 -4040 19340 -4020
rect 19260 -4100 19340 -4040
rect 19400 -4080 19460 -4020
rect 19460 -4080 19480 -4020
rect 19400 -4100 19480 -4080
rect 19500 -4040 19580 -4020
rect 19500 -4100 19580 -4040
rect 19020 -4200 19100 -4140
rect 19020 -4220 19100 -4200
rect 19120 -4200 19140 -4140
rect 19140 -4200 19200 -4140
rect 19120 -4220 19200 -4200
rect 19260 -4200 19340 -4140
rect 19260 -4220 19340 -4200
rect 19400 -4200 19460 -4140
rect 19460 -4200 19480 -4140
rect 19400 -4220 19480 -4200
rect 19500 -4200 19580 -4140
rect 19500 -4220 19580 -4200
<< metal4 >>
rect 1200 400 25600 1000
rect 1200 200 1440 400
rect 6800 240 7040 400
rect 10000 -3420 10600 400
rect 10000 -3500 10020 -3420
rect 10100 -3500 10120 -3420
rect 10200 -3500 10260 -3420
rect 10340 -3500 10400 -3420
rect 10480 -3500 10500 -3420
rect 10580 -3500 10600 -3420
rect 10000 -3560 10600 -3500
rect 10000 -3640 10020 -3560
rect 10100 -3640 10120 -3560
rect 10200 -3640 10260 -3560
rect 10340 -3640 10400 -3560
rect 10480 -3640 10500 -3560
rect 10580 -3640 10600 -3560
rect 10000 -3700 10600 -3640
rect 10000 -3780 10020 -3700
rect 10100 -3780 10120 -3700
rect 10200 -3780 10260 -3700
rect 10340 -3780 10400 -3700
rect 10480 -3780 10500 -3700
rect 10580 -3780 10600 -3700
rect 10000 -3800 10600 -3780
rect 16200 -3420 16800 400
rect 19720 240 19960 400
rect 25360 240 25600 400
rect 16200 -3500 16220 -3420
rect 16300 -3500 16320 -3420
rect 16400 -3500 16460 -3420
rect 16540 -3500 16600 -3420
rect 16680 -3500 16700 -3420
rect 16780 -3500 16800 -3420
rect 16200 -3560 16800 -3500
rect 16200 -3640 16220 -3560
rect 16300 -3640 16320 -3560
rect 16400 -3640 16460 -3560
rect 16540 -3640 16600 -3560
rect 16680 -3640 16700 -3560
rect 16780 -3640 16800 -3560
rect 16200 -3700 16800 -3640
rect 16200 -3780 16220 -3700
rect 16300 -3780 16320 -3700
rect 16400 -3780 16460 -3700
rect 16540 -3780 16600 -3700
rect 16680 -3780 16700 -3700
rect 16780 -3780 16800 -3700
rect 16200 -3800 16800 -3780
rect 7200 -4020 7800 -4000
rect 7200 -4100 7220 -4020
rect 7300 -4100 7320 -4020
rect 7400 -4100 7460 -4020
rect 7540 -4100 7600 -4020
rect 7680 -4100 7700 -4020
rect 7780 -4100 7800 -4020
rect 7200 -4140 7800 -4100
rect 7200 -4220 7220 -4140
rect 7300 -4220 7320 -4140
rect 7400 -4220 7460 -4140
rect 7540 -4220 7600 -4140
rect 7680 -4220 7700 -4140
rect 7780 -4220 7800 -4140
rect -1600 -10600 -1320 -10400
rect 4020 -10600 4280 -10400
rect 7200 -10600 7800 -4220
rect 19000 -4020 19600 -4000
rect 19000 -4100 19020 -4020
rect 19100 -4100 19120 -4020
rect 19200 -4100 19260 -4020
rect 19340 -4100 19400 -4020
rect 19480 -4100 19500 -4020
rect 19580 -4100 19600 -4020
rect 19000 -4140 19600 -4100
rect 19000 -4220 19020 -4140
rect 19100 -4220 19120 -4140
rect 19200 -4220 19260 -4140
rect 19340 -4220 19400 -4140
rect 19480 -4220 19500 -4140
rect 19580 -4220 19600 -4140
rect 19000 -10600 19600 -4220
rect 22500 -10600 22760 -10380
rect 28120 -10600 28400 -10380
rect -1600 -11200 28400 -10600
use sky130_fd_pr__cap_mim_m3_1_RK594X  sky130_fd_pr__cap_mim_m3_1_RK594X_0
timestamp 1770370310
transform -1 0 25292 0 -1 -5080
box -5492 -5320 5492 5320
use sky130_fd_pr__cap_mim_m3_1_RK594X  sky130_fd_pr__cap_mim_m3_1_RK594X_1
timestamp 1770370310
transform 1 0 1492 0 1 -5080
box -5492 -5320 5492 5320
use sky130_fd_pr__nfet_g5v0d10v5_686LYQ  sky130_fd_pr__nfet_g5v0d10v5_686LYQ_0
timestamp 1770112220
transform 1 0 8565 0 1 -6513
box -645 -807 645 807
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_0
timestamp 1770105080
transform 1 0 11847 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_1
timestamp 1770105080
transform 1 0 10047 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_2
timestamp 1770105080
transform 1 0 10487 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_3
timestamp 1770105080
transform 1 0 10927 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_4
timestamp 1770105080
transform 1 0 12287 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_5
timestamp 1770105080
transform 1 0 12727 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_6
timestamp 1770105080
transform 1 0 14047 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_7
timestamp 1770105080
transform 1 0 14487 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_8
timestamp 1770105080
transform 1 0 14927 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_9
timestamp 1770105080
transform 1 0 15847 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_10
timestamp 1770105080
transform 1 0 16287 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_838SN6  sky130_fd_pr__nfet_g5v0d10v5_838SN6_11
timestamp 1770105080
transform 1 0 16727 0 1 -6268
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_DNNC3W  sky130_fd_pr__nfet_g5v0d10v5_DNNC3W_0
timestamp 1770112220
transform 1 0 16127 0 1 -8093
box -187 -807 187 807
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_0
timestamp 1770105080
transform 1 0 11847 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_1
timestamp 1770105080
transform 1 0 10047 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_2
timestamp 1770105080
transform 1 0 10487 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_3
timestamp 1770105080
transform 1 0 10927 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_4
timestamp 1770105080
transform 1 0 12287 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_5
timestamp 1770105080
transform 1 0 12727 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_6
timestamp 1770105080
transform 1 0 14047 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_7
timestamp 1770105080
transform 1 0 14487 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_8
timestamp 1770105080
transform 1 0 14927 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_9
timestamp 1770105080
transform 1 0 15847 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_10
timestamp 1770105080
transform 1 0 16287 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7  sky130_fd_pr__nfet_g5v0d10v5_QN6TJ7_11
timestamp 1770105080
transform 1 0 16727 0 1 -4628
box -187 -532 187 532
use sky130_fd_pr__pfet_g5v0d10v5_AXYYHE  sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_0
timestamp 1770181000
transform 1 0 8633 0 1 -4436
box -333 -564 333 602
use sky130_fd_pr__pfet_g5v0d10v5_AXYYHE  sky130_fd_pr__pfet_g5v0d10v5_AXYYHE_1
timestamp 1770181000
transform 1 0 18213 0 1 -4416
box -333 -564 333 602
use sky130_fd_pr__pfet_g5v0d10v5_DETAA8  sky130_fd_pr__pfet_g5v0d10v5_DETAA8_0
timestamp 1770112220
transform 1 0 8667 0 1 -2236
box -1327 -1064 1327 1102
use sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y  sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y_0
timestamp 1770112220
transform 1 0 16133 0 1 -1816
box -253 -1004 253 1042
use sky130_fd_pr__pfet_g5v0d10v5_Y7F49Y  XM2
timestamp 1770196220
transform 1 0 13334 0 1 -1821
box -2559 -1004 2559 1042
use sky130_fd_pr__pfet_g5v0d10v5_DU7D3Y  XM4
timestamp 1770112220
transform 1 0 10593 0 1 -1816
box -253 -1004 253 1042
use sky130_fd_pr__nfet_g5v0d10v5_DQUD5W  XM24
timestamp 1770112220
transform 1 0 13373 0 1 -8093
box -2493 -807 2493 807
use sky130_fd_pr__nfet_g5v0d10v5_DNNC3W  XM25
timestamp 1770112220
transform 1 0 10627 0 1 -8093
box -187 -807 187 807
use sky130_fd_pr__pfet_g5v0d10v5_DETAA8  XM27
timestamp 1770112220
transform 1 0 18107 0 1 -2236
box -1327 -1064 1327 1102
use sky130_fd_pr__nfet_g5v0d10v5_686LYQ  XM28
timestamp 1770112220
transform 1 0 18225 0 1 -6533
box -645 -807 645 807
<< labels >>
flabel metal1 12920 -180 13120 20 0 FreeSans 800 0 0 0 VDD
port 17 nsew
flabel metal1 14400 -9700 14600 -9500 0 FreeSans 256 0 0 0 VSS
port 11 nsew
flabel metal1 9400 -10300 9600 -10100 0 FreeSans 256 0 0 0 VP
port 3 nsew
flabel metal1 17200 -10300 17400 -10100 0 FreeSans 256 0 0 0 VN
port 4 nsew
flabel metal1 13300 -10900 13500 -10700 0 FreeSans 256 0 0 0 IBIAS
port 9 nsew
flabel metal1 8340 -11680 8540 -11480 0 FreeSans 800 0 0 0 OUT
port 14 nsew
<< end >>
