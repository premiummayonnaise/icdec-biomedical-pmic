magic
tech sky130A
magscale 1 2
timestamp 1769076474
<< error_p >>
rect -511 473 511 477
rect -511 -405 -481 473
rect -445 407 445 411
rect -445 -339 -415 407
rect 415 -339 445 407
rect 481 -405 511 473
<< nwell >>
rect -481 -439 481 473
<< mvpmos >>
rect -387 -339 -237 411
rect -179 -339 -29 411
rect 29 -339 179 411
rect 237 -339 387 411
<< mvpdiff >>
rect -445 399 -387 411
rect -445 -327 -433 399
rect -399 -327 -387 399
rect -445 -339 -387 -327
rect -237 399 -179 411
rect -237 -327 -225 399
rect -191 -327 -179 399
rect -237 -339 -179 -327
rect -29 399 29 411
rect -29 -327 -17 399
rect 17 -327 29 399
rect -29 -339 29 -327
rect 179 399 237 411
rect 179 -327 191 399
rect 225 -327 237 399
rect 179 -339 237 -327
rect 387 399 445 411
rect 387 -327 399 399
rect 433 -327 445 399
rect 387 -339 445 -327
<< mvpdiffc >>
rect -433 -327 -399 399
rect -225 -327 -191 399
rect -17 -327 17 399
rect 191 -327 225 399
rect 399 -327 433 399
<< poly >>
rect -387 411 -237 437
rect -179 411 -29 437
rect 29 411 179 437
rect 237 411 387 437
rect -387 -386 -237 -339
rect -387 -420 -371 -386
rect -253 -420 -237 -386
rect -387 -436 -237 -420
rect -179 -386 -29 -339
rect -179 -420 -163 -386
rect -45 -420 -29 -386
rect -179 -436 -29 -420
rect 29 -386 179 -339
rect 29 -420 45 -386
rect 163 -420 179 -386
rect 29 -436 179 -420
rect 237 -386 387 -339
rect 237 -420 253 -386
rect 371 -420 387 -386
rect 237 -436 387 -420
<< polycont >>
rect -371 -420 -253 -386
rect -163 -420 -45 -386
rect 45 -420 163 -386
rect 253 -420 371 -386
<< locali >>
rect -433 399 -399 415
rect -433 -343 -399 -327
rect -225 399 -191 415
rect -225 -343 -191 -327
rect -17 399 17 415
rect -17 -343 17 -327
rect 191 399 225 415
rect 191 -343 225 -327
rect 399 399 433 415
rect 399 -343 433 -327
rect -387 -420 -371 -386
rect -253 -420 -237 -386
rect -179 -420 -163 -386
rect -45 -420 -29 -386
rect 29 -420 45 -386
rect 163 -420 179 -386
rect 237 -420 253 -386
rect 371 -420 387 -386
<< viali >>
rect -433 -327 -399 399
rect -225 -327 -191 399
rect -17 -327 17 399
rect 191 -327 225 399
rect 399 -327 433 399
rect -371 -420 -253 -386
rect -163 -420 -45 -386
rect 45 -420 163 -386
rect 253 -420 371 -386
<< metal1 >>
rect -439 399 -393 411
rect -439 -327 -433 399
rect -399 -327 -393 399
rect -439 -339 -393 -327
rect -231 399 -185 411
rect -231 -327 -225 399
rect -191 -327 -185 399
rect -231 -339 -185 -327
rect -23 399 23 411
rect -23 -327 -17 399
rect 17 -327 23 399
rect -23 -339 23 -327
rect 185 399 231 411
rect 185 -327 191 399
rect 225 -327 231 399
rect 185 -339 231 -327
rect 393 399 439 411
rect 393 -327 399 399
rect 433 -327 439 399
rect 393 -339 439 -327
rect -383 -386 -241 -380
rect -383 -420 -371 -386
rect -253 -420 -241 -386
rect -383 -426 -241 -420
rect -175 -386 -33 -380
rect -175 -420 -163 -386
rect -45 -420 -33 -386
rect -175 -426 -33 -420
rect 33 -386 175 -380
rect 33 -420 45 -386
rect 163 -420 175 -386
rect 33 -426 175 -420
rect 241 -386 383 -380
rect 241 -420 253 -386
rect 371 -420 383 -386
rect 241 -426 383 -420
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3.75 l 0.75 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
