magic
tech sky130A
magscale 1 2
timestamp 1768990256
<< error_p >>
rect -3459 1098 3459 1102
rect -3459 -1030 -3429 1098
rect -3393 1032 -3027 1036
rect -2965 1032 -2599 1036
rect -2537 1032 -2171 1036
rect -2109 1032 -1743 1036
rect -1681 1032 -1315 1036
rect -1253 1032 -887 1036
rect -825 1032 -459 1036
rect -397 1032 -31 1036
rect 31 1032 397 1036
rect 459 1032 825 1036
rect 887 1032 1253 1036
rect 1315 1032 1681 1036
rect 1743 1032 2109 1036
rect 2171 1032 2537 1036
rect 2599 1032 2965 1036
rect 3027 1032 3393 1036
rect -3393 -964 -3363 1032
rect 3363 -964 3393 1032
rect 3429 -1030 3459 1098
<< nwell >>
rect -3429 -1064 3429 1098
<< mvpmos >>
rect -3335 -964 -3085 1036
rect -2907 -964 -2657 1036
rect -2479 -964 -2229 1036
rect -2051 -964 -1801 1036
rect -1623 -964 -1373 1036
rect -1195 -964 -945 1036
rect -767 -964 -517 1036
rect -339 -964 -89 1036
rect 89 -964 339 1036
rect 517 -964 767 1036
rect 945 -964 1195 1036
rect 1373 -964 1623 1036
rect 1801 -964 2051 1036
rect 2229 -964 2479 1036
rect 2657 -964 2907 1036
rect 3085 -964 3335 1036
<< mvpdiff >>
rect -3393 1024 -3335 1036
rect -3393 -952 -3381 1024
rect -3347 -952 -3335 1024
rect -3393 -964 -3335 -952
rect -3085 1024 -3027 1036
rect -3085 -952 -3073 1024
rect -3039 -952 -3027 1024
rect -3085 -964 -3027 -952
rect -2965 1024 -2907 1036
rect -2965 -952 -2953 1024
rect -2919 -952 -2907 1024
rect -2965 -964 -2907 -952
rect -2657 1024 -2599 1036
rect -2657 -952 -2645 1024
rect -2611 -952 -2599 1024
rect -2657 -964 -2599 -952
rect -2537 1024 -2479 1036
rect -2537 -952 -2525 1024
rect -2491 -952 -2479 1024
rect -2537 -964 -2479 -952
rect -2229 1024 -2171 1036
rect -2229 -952 -2217 1024
rect -2183 -952 -2171 1024
rect -2229 -964 -2171 -952
rect -2109 1024 -2051 1036
rect -2109 -952 -2097 1024
rect -2063 -952 -2051 1024
rect -2109 -964 -2051 -952
rect -1801 1024 -1743 1036
rect -1801 -952 -1789 1024
rect -1755 -952 -1743 1024
rect -1801 -964 -1743 -952
rect -1681 1024 -1623 1036
rect -1681 -952 -1669 1024
rect -1635 -952 -1623 1024
rect -1681 -964 -1623 -952
rect -1373 1024 -1315 1036
rect -1373 -952 -1361 1024
rect -1327 -952 -1315 1024
rect -1373 -964 -1315 -952
rect -1253 1024 -1195 1036
rect -1253 -952 -1241 1024
rect -1207 -952 -1195 1024
rect -1253 -964 -1195 -952
rect -945 1024 -887 1036
rect -945 -952 -933 1024
rect -899 -952 -887 1024
rect -945 -964 -887 -952
rect -825 1024 -767 1036
rect -825 -952 -813 1024
rect -779 -952 -767 1024
rect -825 -964 -767 -952
rect -517 1024 -459 1036
rect -517 -952 -505 1024
rect -471 -952 -459 1024
rect -517 -964 -459 -952
rect -397 1024 -339 1036
rect -397 -952 -385 1024
rect -351 -952 -339 1024
rect -397 -964 -339 -952
rect -89 1024 -31 1036
rect -89 -952 -77 1024
rect -43 -952 -31 1024
rect -89 -964 -31 -952
rect 31 1024 89 1036
rect 31 -952 43 1024
rect 77 -952 89 1024
rect 31 -964 89 -952
rect 339 1024 397 1036
rect 339 -952 351 1024
rect 385 -952 397 1024
rect 339 -964 397 -952
rect 459 1024 517 1036
rect 459 -952 471 1024
rect 505 -952 517 1024
rect 459 -964 517 -952
rect 767 1024 825 1036
rect 767 -952 779 1024
rect 813 -952 825 1024
rect 767 -964 825 -952
rect 887 1024 945 1036
rect 887 -952 899 1024
rect 933 -952 945 1024
rect 887 -964 945 -952
rect 1195 1024 1253 1036
rect 1195 -952 1207 1024
rect 1241 -952 1253 1024
rect 1195 -964 1253 -952
rect 1315 1024 1373 1036
rect 1315 -952 1327 1024
rect 1361 -952 1373 1024
rect 1315 -964 1373 -952
rect 1623 1024 1681 1036
rect 1623 -952 1635 1024
rect 1669 -952 1681 1024
rect 1623 -964 1681 -952
rect 1743 1024 1801 1036
rect 1743 -952 1755 1024
rect 1789 -952 1801 1024
rect 1743 -964 1801 -952
rect 2051 1024 2109 1036
rect 2051 -952 2063 1024
rect 2097 -952 2109 1024
rect 2051 -964 2109 -952
rect 2171 1024 2229 1036
rect 2171 -952 2183 1024
rect 2217 -952 2229 1024
rect 2171 -964 2229 -952
rect 2479 1024 2537 1036
rect 2479 -952 2491 1024
rect 2525 -952 2537 1024
rect 2479 -964 2537 -952
rect 2599 1024 2657 1036
rect 2599 -952 2611 1024
rect 2645 -952 2657 1024
rect 2599 -964 2657 -952
rect 2907 1024 2965 1036
rect 2907 -952 2919 1024
rect 2953 -952 2965 1024
rect 2907 -964 2965 -952
rect 3027 1024 3085 1036
rect 3027 -952 3039 1024
rect 3073 -952 3085 1024
rect 3027 -964 3085 -952
rect 3335 1024 3393 1036
rect 3335 -952 3347 1024
rect 3381 -952 3393 1024
rect 3335 -964 3393 -952
<< mvpdiffc >>
rect -3381 -952 -3347 1024
rect -3073 -952 -3039 1024
rect -2953 -952 -2919 1024
rect -2645 -952 -2611 1024
rect -2525 -952 -2491 1024
rect -2217 -952 -2183 1024
rect -2097 -952 -2063 1024
rect -1789 -952 -1755 1024
rect -1669 -952 -1635 1024
rect -1361 -952 -1327 1024
rect -1241 -952 -1207 1024
rect -933 -952 -899 1024
rect -813 -952 -779 1024
rect -505 -952 -471 1024
rect -385 -952 -351 1024
rect -77 -952 -43 1024
rect 43 -952 77 1024
rect 351 -952 385 1024
rect 471 -952 505 1024
rect 779 -952 813 1024
rect 899 -952 933 1024
rect 1207 -952 1241 1024
rect 1327 -952 1361 1024
rect 1635 -952 1669 1024
rect 1755 -952 1789 1024
rect 2063 -952 2097 1024
rect 2183 -952 2217 1024
rect 2491 -952 2525 1024
rect 2611 -952 2645 1024
rect 2919 -952 2953 1024
rect 3039 -952 3073 1024
rect 3347 -952 3381 1024
<< poly >>
rect -3335 1036 -3085 1062
rect -2907 1036 -2657 1062
rect -2479 1036 -2229 1062
rect -2051 1036 -1801 1062
rect -1623 1036 -1373 1062
rect -1195 1036 -945 1062
rect -767 1036 -517 1062
rect -339 1036 -89 1062
rect 89 1036 339 1062
rect 517 1036 767 1062
rect 945 1036 1195 1062
rect 1373 1036 1623 1062
rect 1801 1036 2051 1062
rect 2229 1036 2479 1062
rect 2657 1036 2907 1062
rect 3085 1036 3335 1062
rect -3335 -1011 -3085 -964
rect -3335 -1045 -3319 -1011
rect -3101 -1045 -3085 -1011
rect -3335 -1061 -3085 -1045
rect -2907 -1011 -2657 -964
rect -2907 -1045 -2891 -1011
rect -2673 -1045 -2657 -1011
rect -2907 -1061 -2657 -1045
rect -2479 -1011 -2229 -964
rect -2479 -1045 -2463 -1011
rect -2245 -1045 -2229 -1011
rect -2479 -1061 -2229 -1045
rect -2051 -1011 -1801 -964
rect -2051 -1045 -2035 -1011
rect -1817 -1045 -1801 -1011
rect -2051 -1061 -1801 -1045
rect -1623 -1011 -1373 -964
rect -1623 -1045 -1607 -1011
rect -1389 -1045 -1373 -1011
rect -1623 -1061 -1373 -1045
rect -1195 -1011 -945 -964
rect -1195 -1045 -1179 -1011
rect -961 -1045 -945 -1011
rect -1195 -1061 -945 -1045
rect -767 -1011 -517 -964
rect -767 -1045 -751 -1011
rect -533 -1045 -517 -1011
rect -767 -1061 -517 -1045
rect -339 -1011 -89 -964
rect -339 -1045 -323 -1011
rect -105 -1045 -89 -1011
rect -339 -1061 -89 -1045
rect 89 -1011 339 -964
rect 89 -1045 105 -1011
rect 323 -1045 339 -1011
rect 89 -1061 339 -1045
rect 517 -1011 767 -964
rect 517 -1045 533 -1011
rect 751 -1045 767 -1011
rect 517 -1061 767 -1045
rect 945 -1011 1195 -964
rect 945 -1045 961 -1011
rect 1179 -1045 1195 -1011
rect 945 -1061 1195 -1045
rect 1373 -1011 1623 -964
rect 1373 -1045 1389 -1011
rect 1607 -1045 1623 -1011
rect 1373 -1061 1623 -1045
rect 1801 -1011 2051 -964
rect 1801 -1045 1817 -1011
rect 2035 -1045 2051 -1011
rect 1801 -1061 2051 -1045
rect 2229 -1011 2479 -964
rect 2229 -1045 2245 -1011
rect 2463 -1045 2479 -1011
rect 2229 -1061 2479 -1045
rect 2657 -1011 2907 -964
rect 2657 -1045 2673 -1011
rect 2891 -1045 2907 -1011
rect 2657 -1061 2907 -1045
rect 3085 -1011 3335 -964
rect 3085 -1045 3101 -1011
rect 3319 -1045 3335 -1011
rect 3085 -1061 3335 -1045
<< polycont >>
rect -3319 -1045 -3101 -1011
rect -2891 -1045 -2673 -1011
rect -2463 -1045 -2245 -1011
rect -2035 -1045 -1817 -1011
rect -1607 -1045 -1389 -1011
rect -1179 -1045 -961 -1011
rect -751 -1045 -533 -1011
rect -323 -1045 -105 -1011
rect 105 -1045 323 -1011
rect 533 -1045 751 -1011
rect 961 -1045 1179 -1011
rect 1389 -1045 1607 -1011
rect 1817 -1045 2035 -1011
rect 2245 -1045 2463 -1011
rect 2673 -1045 2891 -1011
rect 3101 -1045 3319 -1011
<< locali >>
rect -3381 1024 -3347 1040
rect -3381 -968 -3347 -952
rect -3073 1024 -3039 1040
rect -3073 -968 -3039 -952
rect -2953 1024 -2919 1040
rect -2953 -968 -2919 -952
rect -2645 1024 -2611 1040
rect -2645 -968 -2611 -952
rect -2525 1024 -2491 1040
rect -2525 -968 -2491 -952
rect -2217 1024 -2183 1040
rect -2217 -968 -2183 -952
rect -2097 1024 -2063 1040
rect -2097 -968 -2063 -952
rect -1789 1024 -1755 1040
rect -1789 -968 -1755 -952
rect -1669 1024 -1635 1040
rect -1669 -968 -1635 -952
rect -1361 1024 -1327 1040
rect -1361 -968 -1327 -952
rect -1241 1024 -1207 1040
rect -1241 -968 -1207 -952
rect -933 1024 -899 1040
rect -933 -968 -899 -952
rect -813 1024 -779 1040
rect -813 -968 -779 -952
rect -505 1024 -471 1040
rect -505 -968 -471 -952
rect -385 1024 -351 1040
rect -385 -968 -351 -952
rect -77 1024 -43 1040
rect -77 -968 -43 -952
rect 43 1024 77 1040
rect 43 -968 77 -952
rect 351 1024 385 1040
rect 351 -968 385 -952
rect 471 1024 505 1040
rect 471 -968 505 -952
rect 779 1024 813 1040
rect 779 -968 813 -952
rect 899 1024 933 1040
rect 899 -968 933 -952
rect 1207 1024 1241 1040
rect 1207 -968 1241 -952
rect 1327 1024 1361 1040
rect 1327 -968 1361 -952
rect 1635 1024 1669 1040
rect 1635 -968 1669 -952
rect 1755 1024 1789 1040
rect 1755 -968 1789 -952
rect 2063 1024 2097 1040
rect 2063 -968 2097 -952
rect 2183 1024 2217 1040
rect 2183 -968 2217 -952
rect 2491 1024 2525 1040
rect 2491 -968 2525 -952
rect 2611 1024 2645 1040
rect 2611 -968 2645 -952
rect 2919 1024 2953 1040
rect 2919 -968 2953 -952
rect 3039 1024 3073 1040
rect 3039 -968 3073 -952
rect 3347 1024 3381 1040
rect 3347 -968 3381 -952
rect -3335 -1045 -3319 -1011
rect -3101 -1045 -3085 -1011
rect -2907 -1045 -2891 -1011
rect -2673 -1045 -2657 -1011
rect -2479 -1045 -2463 -1011
rect -2245 -1045 -2229 -1011
rect -2051 -1045 -2035 -1011
rect -1817 -1045 -1801 -1011
rect -1623 -1045 -1607 -1011
rect -1389 -1045 -1373 -1011
rect -1195 -1045 -1179 -1011
rect -961 -1045 -945 -1011
rect -767 -1045 -751 -1011
rect -533 -1045 -517 -1011
rect -339 -1045 -323 -1011
rect -105 -1045 -89 -1011
rect 89 -1045 105 -1011
rect 323 -1045 339 -1011
rect 517 -1045 533 -1011
rect 751 -1045 767 -1011
rect 945 -1045 961 -1011
rect 1179 -1045 1195 -1011
rect 1373 -1045 1389 -1011
rect 1607 -1045 1623 -1011
rect 1801 -1045 1817 -1011
rect 2035 -1045 2051 -1011
rect 2229 -1045 2245 -1011
rect 2463 -1045 2479 -1011
rect 2657 -1045 2673 -1011
rect 2891 -1045 2907 -1011
rect 3085 -1045 3101 -1011
rect 3319 -1045 3335 -1011
<< viali >>
rect -3381 -952 -3347 1024
rect -3073 -952 -3039 1024
rect -2953 -952 -2919 1024
rect -2645 -952 -2611 1024
rect -2525 -952 -2491 1024
rect -2217 -952 -2183 1024
rect -2097 -952 -2063 1024
rect -1789 -952 -1755 1024
rect -1669 -952 -1635 1024
rect -1361 -952 -1327 1024
rect -1241 -952 -1207 1024
rect -933 -952 -899 1024
rect -813 -952 -779 1024
rect -505 -952 -471 1024
rect -385 -952 -351 1024
rect -77 -952 -43 1024
rect 43 -952 77 1024
rect 351 -952 385 1024
rect 471 -952 505 1024
rect 779 -952 813 1024
rect 899 -952 933 1024
rect 1207 -952 1241 1024
rect 1327 -952 1361 1024
rect 1635 -952 1669 1024
rect 1755 -952 1789 1024
rect 2063 -952 2097 1024
rect 2183 -952 2217 1024
rect 2491 -952 2525 1024
rect 2611 -952 2645 1024
rect 2919 -952 2953 1024
rect 3039 -952 3073 1024
rect 3347 -952 3381 1024
rect -3319 -1045 -3101 -1011
rect -2891 -1045 -2673 -1011
rect -2463 -1045 -2245 -1011
rect -2035 -1045 -1817 -1011
rect -1607 -1045 -1389 -1011
rect -1179 -1045 -961 -1011
rect -751 -1045 -533 -1011
rect -323 -1045 -105 -1011
rect 105 -1045 323 -1011
rect 533 -1045 751 -1011
rect 961 -1045 1179 -1011
rect 1389 -1045 1607 -1011
rect 1817 -1045 2035 -1011
rect 2245 -1045 2463 -1011
rect 2673 -1045 2891 -1011
rect 3101 -1045 3319 -1011
<< metal1 >>
rect -3387 1024 -3341 1036
rect -3387 -952 -3381 1024
rect -3347 -952 -3341 1024
rect -3387 -964 -3341 -952
rect -3079 1024 -3033 1036
rect -3079 -952 -3073 1024
rect -3039 -952 -3033 1024
rect -3079 -964 -3033 -952
rect -2959 1024 -2913 1036
rect -2959 -952 -2953 1024
rect -2919 -952 -2913 1024
rect -2959 -964 -2913 -952
rect -2651 1024 -2605 1036
rect -2651 -952 -2645 1024
rect -2611 -952 -2605 1024
rect -2651 -964 -2605 -952
rect -2531 1024 -2485 1036
rect -2531 -952 -2525 1024
rect -2491 -952 -2485 1024
rect -2531 -964 -2485 -952
rect -2223 1024 -2177 1036
rect -2223 -952 -2217 1024
rect -2183 -952 -2177 1024
rect -2223 -964 -2177 -952
rect -2103 1024 -2057 1036
rect -2103 -952 -2097 1024
rect -2063 -952 -2057 1024
rect -2103 -964 -2057 -952
rect -1795 1024 -1749 1036
rect -1795 -952 -1789 1024
rect -1755 -952 -1749 1024
rect -1795 -964 -1749 -952
rect -1675 1024 -1629 1036
rect -1675 -952 -1669 1024
rect -1635 -952 -1629 1024
rect -1675 -964 -1629 -952
rect -1367 1024 -1321 1036
rect -1367 -952 -1361 1024
rect -1327 -952 -1321 1024
rect -1367 -964 -1321 -952
rect -1247 1024 -1201 1036
rect -1247 -952 -1241 1024
rect -1207 -952 -1201 1024
rect -1247 -964 -1201 -952
rect -939 1024 -893 1036
rect -939 -952 -933 1024
rect -899 -952 -893 1024
rect -939 -964 -893 -952
rect -819 1024 -773 1036
rect -819 -952 -813 1024
rect -779 -952 -773 1024
rect -819 -964 -773 -952
rect -511 1024 -465 1036
rect -511 -952 -505 1024
rect -471 -952 -465 1024
rect -511 -964 -465 -952
rect -391 1024 -345 1036
rect -391 -952 -385 1024
rect -351 -952 -345 1024
rect -391 -964 -345 -952
rect -83 1024 -37 1036
rect -83 -952 -77 1024
rect -43 -952 -37 1024
rect -83 -964 -37 -952
rect 37 1024 83 1036
rect 37 -952 43 1024
rect 77 -952 83 1024
rect 37 -964 83 -952
rect 345 1024 391 1036
rect 345 -952 351 1024
rect 385 -952 391 1024
rect 345 -964 391 -952
rect 465 1024 511 1036
rect 465 -952 471 1024
rect 505 -952 511 1024
rect 465 -964 511 -952
rect 773 1024 819 1036
rect 773 -952 779 1024
rect 813 -952 819 1024
rect 773 -964 819 -952
rect 893 1024 939 1036
rect 893 -952 899 1024
rect 933 -952 939 1024
rect 893 -964 939 -952
rect 1201 1024 1247 1036
rect 1201 -952 1207 1024
rect 1241 -952 1247 1024
rect 1201 -964 1247 -952
rect 1321 1024 1367 1036
rect 1321 -952 1327 1024
rect 1361 -952 1367 1024
rect 1321 -964 1367 -952
rect 1629 1024 1675 1036
rect 1629 -952 1635 1024
rect 1669 -952 1675 1024
rect 1629 -964 1675 -952
rect 1749 1024 1795 1036
rect 1749 -952 1755 1024
rect 1789 -952 1795 1024
rect 1749 -964 1795 -952
rect 2057 1024 2103 1036
rect 2057 -952 2063 1024
rect 2097 -952 2103 1024
rect 2057 -964 2103 -952
rect 2177 1024 2223 1036
rect 2177 -952 2183 1024
rect 2217 -952 2223 1024
rect 2177 -964 2223 -952
rect 2485 1024 2531 1036
rect 2485 -952 2491 1024
rect 2525 -952 2531 1024
rect 2485 -964 2531 -952
rect 2605 1024 2651 1036
rect 2605 -952 2611 1024
rect 2645 -952 2651 1024
rect 2605 -964 2651 -952
rect 2913 1024 2959 1036
rect 2913 -952 2919 1024
rect 2953 -952 2959 1024
rect 2913 -964 2959 -952
rect 3033 1024 3079 1036
rect 3033 -952 3039 1024
rect 3073 -952 3079 1024
rect 3033 -964 3079 -952
rect 3341 1024 3387 1036
rect 3341 -952 3347 1024
rect 3381 -952 3387 1024
rect 3341 -964 3387 -952
rect -3331 -1011 -3089 -1005
rect -3331 -1045 -3319 -1011
rect -3101 -1045 -3089 -1011
rect -3331 -1051 -3089 -1045
rect -2903 -1011 -2661 -1005
rect -2903 -1045 -2891 -1011
rect -2673 -1045 -2661 -1011
rect -2903 -1051 -2661 -1045
rect -2475 -1011 -2233 -1005
rect -2475 -1045 -2463 -1011
rect -2245 -1045 -2233 -1011
rect -2475 -1051 -2233 -1045
rect -2047 -1011 -1805 -1005
rect -2047 -1045 -2035 -1011
rect -1817 -1045 -1805 -1011
rect -2047 -1051 -1805 -1045
rect -1619 -1011 -1377 -1005
rect -1619 -1045 -1607 -1011
rect -1389 -1045 -1377 -1011
rect -1619 -1051 -1377 -1045
rect -1191 -1011 -949 -1005
rect -1191 -1045 -1179 -1011
rect -961 -1045 -949 -1011
rect -1191 -1051 -949 -1045
rect -763 -1011 -521 -1005
rect -763 -1045 -751 -1011
rect -533 -1045 -521 -1011
rect -763 -1051 -521 -1045
rect -335 -1011 -93 -1005
rect -335 -1045 -323 -1011
rect -105 -1045 -93 -1011
rect -335 -1051 -93 -1045
rect 93 -1011 335 -1005
rect 93 -1045 105 -1011
rect 323 -1045 335 -1011
rect 93 -1051 335 -1045
rect 521 -1011 763 -1005
rect 521 -1045 533 -1011
rect 751 -1045 763 -1011
rect 521 -1051 763 -1045
rect 949 -1011 1191 -1005
rect 949 -1045 961 -1011
rect 1179 -1045 1191 -1011
rect 949 -1051 1191 -1045
rect 1377 -1011 1619 -1005
rect 1377 -1045 1389 -1011
rect 1607 -1045 1619 -1011
rect 1377 -1051 1619 -1045
rect 1805 -1011 2047 -1005
rect 1805 -1045 1817 -1011
rect 2035 -1045 2047 -1011
rect 1805 -1051 2047 -1045
rect 2233 -1011 2475 -1005
rect 2233 -1045 2245 -1011
rect 2463 -1045 2475 -1011
rect 2233 -1051 2475 -1045
rect 2661 -1011 2903 -1005
rect 2661 -1045 2673 -1011
rect 2891 -1045 2903 -1011
rect 2661 -1051 2903 -1045
rect 3089 -1011 3331 -1005
rect 3089 -1045 3101 -1011
rect 3319 -1045 3331 -1011
rect 3089 -1051 3331 -1045
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 1.25 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
