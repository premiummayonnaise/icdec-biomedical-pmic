magic
tech sky130A
magscale 1 2
timestamp 1770023980
<< nwell >>
rect -2693 -1297 2693 1297
<< mvpmos >>
rect -2435 -1000 -2185 1000
rect -2127 -1000 -1877 1000
rect -1819 -1000 -1569 1000
rect -1511 -1000 -1261 1000
rect -1203 -1000 -953 1000
rect -895 -1000 -645 1000
rect -587 -1000 -337 1000
rect -279 -1000 -29 1000
rect 29 -1000 279 1000
rect 337 -1000 587 1000
rect 645 -1000 895 1000
rect 953 -1000 1203 1000
rect 1261 -1000 1511 1000
rect 1569 -1000 1819 1000
rect 1877 -1000 2127 1000
rect 2185 -1000 2435 1000
<< mvpdiff >>
rect -2493 988 -2435 1000
rect -2493 -988 -2481 988
rect -2447 -988 -2435 988
rect -2493 -1000 -2435 -988
rect -2185 988 -2127 1000
rect -2185 -988 -2173 988
rect -2139 -988 -2127 988
rect -2185 -1000 -2127 -988
rect -1877 988 -1819 1000
rect -1877 -988 -1865 988
rect -1831 -988 -1819 988
rect -1877 -1000 -1819 -988
rect -1569 988 -1511 1000
rect -1569 -988 -1557 988
rect -1523 -988 -1511 988
rect -1569 -1000 -1511 -988
rect -1261 988 -1203 1000
rect -1261 -988 -1249 988
rect -1215 -988 -1203 988
rect -1261 -1000 -1203 -988
rect -953 988 -895 1000
rect -953 -988 -941 988
rect -907 -988 -895 988
rect -953 -1000 -895 -988
rect -645 988 -587 1000
rect -645 -988 -633 988
rect -599 -988 -587 988
rect -645 -1000 -587 -988
rect -337 988 -279 1000
rect -337 -988 -325 988
rect -291 -988 -279 988
rect -337 -1000 -279 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 279 988 337 1000
rect 279 -988 291 988
rect 325 -988 337 988
rect 279 -1000 337 -988
rect 587 988 645 1000
rect 587 -988 599 988
rect 633 -988 645 988
rect 587 -1000 645 -988
rect 895 988 953 1000
rect 895 -988 907 988
rect 941 -988 953 988
rect 895 -1000 953 -988
rect 1203 988 1261 1000
rect 1203 -988 1215 988
rect 1249 -988 1261 988
rect 1203 -1000 1261 -988
rect 1511 988 1569 1000
rect 1511 -988 1523 988
rect 1557 -988 1569 988
rect 1511 -1000 1569 -988
rect 1819 988 1877 1000
rect 1819 -988 1831 988
rect 1865 -988 1877 988
rect 1819 -1000 1877 -988
rect 2127 988 2185 1000
rect 2127 -988 2139 988
rect 2173 -988 2185 988
rect 2127 -1000 2185 -988
rect 2435 988 2493 1000
rect 2435 -988 2447 988
rect 2481 -988 2493 988
rect 2435 -1000 2493 -988
<< mvpdiffc >>
rect -2481 -988 -2447 988
rect -2173 -988 -2139 988
rect -1865 -988 -1831 988
rect -1557 -988 -1523 988
rect -1249 -988 -1215 988
rect -941 -988 -907 988
rect -633 -988 -599 988
rect -325 -988 -291 988
rect -17 -988 17 988
rect 291 -988 325 988
rect 599 -988 633 988
rect 907 -988 941 988
rect 1215 -988 1249 988
rect 1523 -988 1557 988
rect 1831 -988 1865 988
rect 2139 -988 2173 988
rect 2447 -988 2481 988
<< mvnsubdiff >>
rect -2627 1219 2627 1231
rect -2627 1185 -2519 1219
rect 2519 1185 2627 1219
rect -2627 1173 2627 1185
rect -2627 1123 -2569 1173
rect -2627 -1123 -2615 1123
rect -2581 -1123 -2569 1123
rect 2569 1123 2627 1173
rect -2627 -1173 -2569 -1123
rect 2569 -1123 2581 1123
rect 2615 -1123 2627 1123
rect 2569 -1173 2627 -1123
rect -2627 -1185 2627 -1173
rect -2627 -1219 -2519 -1185
rect 2519 -1219 2627 -1185
rect -2627 -1231 2627 -1219
<< mvnsubdiffcont >>
rect -2519 1185 2519 1219
rect -2615 -1123 -2581 1123
rect 2581 -1123 2615 1123
rect -2519 -1219 2519 -1185
<< poly >>
rect -2435 1081 -2185 1097
rect -2435 1047 -2419 1081
rect -2201 1047 -2185 1081
rect -2435 1000 -2185 1047
rect -2127 1081 -1877 1097
rect -2127 1047 -2111 1081
rect -1893 1047 -1877 1081
rect -2127 1000 -1877 1047
rect -1819 1081 -1569 1097
rect -1819 1047 -1803 1081
rect -1585 1047 -1569 1081
rect -1819 1000 -1569 1047
rect -1511 1081 -1261 1097
rect -1511 1047 -1495 1081
rect -1277 1047 -1261 1081
rect -1511 1000 -1261 1047
rect -1203 1081 -953 1097
rect -1203 1047 -1187 1081
rect -969 1047 -953 1081
rect -1203 1000 -953 1047
rect -895 1081 -645 1097
rect -895 1047 -879 1081
rect -661 1047 -645 1081
rect -895 1000 -645 1047
rect -587 1081 -337 1097
rect -587 1047 -571 1081
rect -353 1047 -337 1081
rect -587 1000 -337 1047
rect -279 1081 -29 1097
rect -279 1047 -263 1081
rect -45 1047 -29 1081
rect -279 1000 -29 1047
rect 29 1081 279 1097
rect 29 1047 45 1081
rect 263 1047 279 1081
rect 29 1000 279 1047
rect 337 1081 587 1097
rect 337 1047 353 1081
rect 571 1047 587 1081
rect 337 1000 587 1047
rect 645 1081 895 1097
rect 645 1047 661 1081
rect 879 1047 895 1081
rect 645 1000 895 1047
rect 953 1081 1203 1097
rect 953 1047 969 1081
rect 1187 1047 1203 1081
rect 953 1000 1203 1047
rect 1261 1081 1511 1097
rect 1261 1047 1277 1081
rect 1495 1047 1511 1081
rect 1261 1000 1511 1047
rect 1569 1081 1819 1097
rect 1569 1047 1585 1081
rect 1803 1047 1819 1081
rect 1569 1000 1819 1047
rect 1877 1081 2127 1097
rect 1877 1047 1893 1081
rect 2111 1047 2127 1081
rect 1877 1000 2127 1047
rect 2185 1081 2435 1097
rect 2185 1047 2201 1081
rect 2419 1047 2435 1081
rect 2185 1000 2435 1047
rect -2435 -1047 -2185 -1000
rect -2435 -1081 -2419 -1047
rect -2201 -1081 -2185 -1047
rect -2435 -1097 -2185 -1081
rect -2127 -1047 -1877 -1000
rect -2127 -1081 -2111 -1047
rect -1893 -1081 -1877 -1047
rect -2127 -1097 -1877 -1081
rect -1819 -1047 -1569 -1000
rect -1819 -1081 -1803 -1047
rect -1585 -1081 -1569 -1047
rect -1819 -1097 -1569 -1081
rect -1511 -1047 -1261 -1000
rect -1511 -1081 -1495 -1047
rect -1277 -1081 -1261 -1047
rect -1511 -1097 -1261 -1081
rect -1203 -1047 -953 -1000
rect -1203 -1081 -1187 -1047
rect -969 -1081 -953 -1047
rect -1203 -1097 -953 -1081
rect -895 -1047 -645 -1000
rect -895 -1081 -879 -1047
rect -661 -1081 -645 -1047
rect -895 -1097 -645 -1081
rect -587 -1047 -337 -1000
rect -587 -1081 -571 -1047
rect -353 -1081 -337 -1047
rect -587 -1097 -337 -1081
rect -279 -1047 -29 -1000
rect -279 -1081 -263 -1047
rect -45 -1081 -29 -1047
rect -279 -1097 -29 -1081
rect 29 -1047 279 -1000
rect 29 -1081 45 -1047
rect 263 -1081 279 -1047
rect 29 -1097 279 -1081
rect 337 -1047 587 -1000
rect 337 -1081 353 -1047
rect 571 -1081 587 -1047
rect 337 -1097 587 -1081
rect 645 -1047 895 -1000
rect 645 -1081 661 -1047
rect 879 -1081 895 -1047
rect 645 -1097 895 -1081
rect 953 -1047 1203 -1000
rect 953 -1081 969 -1047
rect 1187 -1081 1203 -1047
rect 953 -1097 1203 -1081
rect 1261 -1047 1511 -1000
rect 1261 -1081 1277 -1047
rect 1495 -1081 1511 -1047
rect 1261 -1097 1511 -1081
rect 1569 -1047 1819 -1000
rect 1569 -1081 1585 -1047
rect 1803 -1081 1819 -1047
rect 1569 -1097 1819 -1081
rect 1877 -1047 2127 -1000
rect 1877 -1081 1893 -1047
rect 2111 -1081 2127 -1047
rect 1877 -1097 2127 -1081
rect 2185 -1047 2435 -1000
rect 2185 -1081 2201 -1047
rect 2419 -1081 2435 -1047
rect 2185 -1097 2435 -1081
<< polycont >>
rect -2419 1047 -2201 1081
rect -2111 1047 -1893 1081
rect -1803 1047 -1585 1081
rect -1495 1047 -1277 1081
rect -1187 1047 -969 1081
rect -879 1047 -661 1081
rect -571 1047 -353 1081
rect -263 1047 -45 1081
rect 45 1047 263 1081
rect 353 1047 571 1081
rect 661 1047 879 1081
rect 969 1047 1187 1081
rect 1277 1047 1495 1081
rect 1585 1047 1803 1081
rect 1893 1047 2111 1081
rect 2201 1047 2419 1081
rect -2419 -1081 -2201 -1047
rect -2111 -1081 -1893 -1047
rect -1803 -1081 -1585 -1047
rect -1495 -1081 -1277 -1047
rect -1187 -1081 -969 -1047
rect -879 -1081 -661 -1047
rect -571 -1081 -353 -1047
rect -263 -1081 -45 -1047
rect 45 -1081 263 -1047
rect 353 -1081 571 -1047
rect 661 -1081 879 -1047
rect 969 -1081 1187 -1047
rect 1277 -1081 1495 -1047
rect 1585 -1081 1803 -1047
rect 1893 -1081 2111 -1047
rect 2201 -1081 2419 -1047
<< locali >>
rect -2615 1185 -2519 1219
rect 2519 1185 2615 1219
rect -2615 1123 -2581 1185
rect 2581 1123 2615 1185
rect -2435 1047 -2419 1081
rect -2201 1047 -2185 1081
rect -2127 1047 -2111 1081
rect -1893 1047 -1877 1081
rect -1819 1047 -1803 1081
rect -1585 1047 -1569 1081
rect -1511 1047 -1495 1081
rect -1277 1047 -1261 1081
rect -1203 1047 -1187 1081
rect -969 1047 -953 1081
rect -895 1047 -879 1081
rect -661 1047 -645 1081
rect -587 1047 -571 1081
rect -353 1047 -337 1081
rect -279 1047 -263 1081
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect 263 1047 279 1081
rect 337 1047 353 1081
rect 571 1047 587 1081
rect 645 1047 661 1081
rect 879 1047 895 1081
rect 953 1047 969 1081
rect 1187 1047 1203 1081
rect 1261 1047 1277 1081
rect 1495 1047 1511 1081
rect 1569 1047 1585 1081
rect 1803 1047 1819 1081
rect 1877 1047 1893 1081
rect 2111 1047 2127 1081
rect 2185 1047 2201 1081
rect 2419 1047 2435 1081
rect -2481 988 -2447 1004
rect -2481 -1004 -2447 -988
rect -2173 988 -2139 1004
rect -2173 -1004 -2139 -988
rect -1865 988 -1831 1004
rect -1865 -1004 -1831 -988
rect -1557 988 -1523 1004
rect -1557 -1004 -1523 -988
rect -1249 988 -1215 1004
rect -1249 -1004 -1215 -988
rect -941 988 -907 1004
rect -941 -1004 -907 -988
rect -633 988 -599 1004
rect -633 -1004 -599 -988
rect -325 988 -291 1004
rect -325 -1004 -291 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 291 988 325 1004
rect 291 -1004 325 -988
rect 599 988 633 1004
rect 599 -1004 633 -988
rect 907 988 941 1004
rect 907 -1004 941 -988
rect 1215 988 1249 1004
rect 1215 -1004 1249 -988
rect 1523 988 1557 1004
rect 1523 -1004 1557 -988
rect 1831 988 1865 1004
rect 1831 -1004 1865 -988
rect 2139 988 2173 1004
rect 2139 -1004 2173 -988
rect 2447 988 2481 1004
rect 2447 -1004 2481 -988
rect -2435 -1081 -2419 -1047
rect -2201 -1081 -2185 -1047
rect -2127 -1081 -2111 -1047
rect -1893 -1081 -1877 -1047
rect -1819 -1081 -1803 -1047
rect -1585 -1081 -1569 -1047
rect -1511 -1081 -1495 -1047
rect -1277 -1081 -1261 -1047
rect -1203 -1081 -1187 -1047
rect -969 -1081 -953 -1047
rect -895 -1081 -879 -1047
rect -661 -1081 -645 -1047
rect -587 -1081 -571 -1047
rect -353 -1081 -337 -1047
rect -279 -1081 -263 -1047
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect 263 -1081 279 -1047
rect 337 -1081 353 -1047
rect 571 -1081 587 -1047
rect 645 -1081 661 -1047
rect 879 -1081 895 -1047
rect 953 -1081 969 -1047
rect 1187 -1081 1203 -1047
rect 1261 -1081 1277 -1047
rect 1495 -1081 1511 -1047
rect 1569 -1081 1585 -1047
rect 1803 -1081 1819 -1047
rect 1877 -1081 1893 -1047
rect 2111 -1081 2127 -1047
rect 2185 -1081 2201 -1047
rect 2419 -1081 2435 -1047
rect -2615 -1185 -2581 -1123
rect 2581 -1185 2615 -1123
rect -2615 -1219 -2519 -1185
rect 2519 -1219 2615 -1185
<< viali >>
rect -2419 1047 -2201 1081
rect -2111 1047 -1893 1081
rect -1803 1047 -1585 1081
rect -1495 1047 -1277 1081
rect -1187 1047 -969 1081
rect -879 1047 -661 1081
rect -571 1047 -353 1081
rect -263 1047 -45 1081
rect 45 1047 263 1081
rect 353 1047 571 1081
rect 661 1047 879 1081
rect 969 1047 1187 1081
rect 1277 1047 1495 1081
rect 1585 1047 1803 1081
rect 1893 1047 2111 1081
rect 2201 1047 2419 1081
rect -2481 -988 -2447 988
rect -2173 -988 -2139 988
rect -1865 -988 -1831 988
rect -1557 -988 -1523 988
rect -1249 -988 -1215 988
rect -941 -988 -907 988
rect -633 -988 -599 988
rect -325 -988 -291 988
rect -17 -988 17 988
rect 291 -988 325 988
rect 599 -988 633 988
rect 907 -988 941 988
rect 1215 -988 1249 988
rect 1523 -988 1557 988
rect 1831 -988 1865 988
rect 2139 -988 2173 988
rect 2447 -988 2481 988
rect -2419 -1081 -2201 -1047
rect -2111 -1081 -1893 -1047
rect -1803 -1081 -1585 -1047
rect -1495 -1081 -1277 -1047
rect -1187 -1081 -969 -1047
rect -879 -1081 -661 -1047
rect -571 -1081 -353 -1047
rect -263 -1081 -45 -1047
rect 45 -1081 263 -1047
rect 353 -1081 571 -1047
rect 661 -1081 879 -1047
rect 969 -1081 1187 -1047
rect 1277 -1081 1495 -1047
rect 1585 -1081 1803 -1047
rect 1893 -1081 2111 -1047
rect 2201 -1081 2419 -1047
<< metal1 >>
rect -2431 1081 -2189 1087
rect -2431 1047 -2419 1081
rect -2201 1047 -2189 1081
rect -2431 1041 -2189 1047
rect -2123 1081 -1881 1087
rect -2123 1047 -2111 1081
rect -1893 1047 -1881 1081
rect -2123 1041 -1881 1047
rect -1815 1081 -1573 1087
rect -1815 1047 -1803 1081
rect -1585 1047 -1573 1081
rect -1815 1041 -1573 1047
rect -1507 1081 -1265 1087
rect -1507 1047 -1495 1081
rect -1277 1047 -1265 1081
rect -1507 1041 -1265 1047
rect -1199 1081 -957 1087
rect -1199 1047 -1187 1081
rect -969 1047 -957 1081
rect -1199 1041 -957 1047
rect -891 1081 -649 1087
rect -891 1047 -879 1081
rect -661 1047 -649 1081
rect -891 1041 -649 1047
rect -583 1081 -341 1087
rect -583 1047 -571 1081
rect -353 1047 -341 1081
rect -583 1041 -341 1047
rect -275 1081 -33 1087
rect -275 1047 -263 1081
rect -45 1047 -33 1081
rect -275 1041 -33 1047
rect 33 1081 275 1087
rect 33 1047 45 1081
rect 263 1047 275 1081
rect 33 1041 275 1047
rect 341 1081 583 1087
rect 341 1047 353 1081
rect 571 1047 583 1081
rect 341 1041 583 1047
rect 649 1081 891 1087
rect 649 1047 661 1081
rect 879 1047 891 1081
rect 649 1041 891 1047
rect 957 1081 1199 1087
rect 957 1047 969 1081
rect 1187 1047 1199 1081
rect 957 1041 1199 1047
rect 1265 1081 1507 1087
rect 1265 1047 1277 1081
rect 1495 1047 1507 1081
rect 1265 1041 1507 1047
rect 1573 1081 1815 1087
rect 1573 1047 1585 1081
rect 1803 1047 1815 1081
rect 1573 1041 1815 1047
rect 1881 1081 2123 1087
rect 1881 1047 1893 1081
rect 2111 1047 2123 1081
rect 1881 1041 2123 1047
rect 2189 1081 2431 1087
rect 2189 1047 2201 1081
rect 2419 1047 2431 1081
rect 2189 1041 2431 1047
rect -2487 988 -2441 1000
rect -2487 -988 -2481 988
rect -2447 -988 -2441 988
rect -2487 -1000 -2441 -988
rect -2179 988 -2133 1000
rect -2179 -988 -2173 988
rect -2139 -988 -2133 988
rect -2179 -1000 -2133 -988
rect -1871 988 -1825 1000
rect -1871 -988 -1865 988
rect -1831 -988 -1825 988
rect -1871 -1000 -1825 -988
rect -1563 988 -1517 1000
rect -1563 -988 -1557 988
rect -1523 -988 -1517 988
rect -1563 -1000 -1517 -988
rect -1255 988 -1209 1000
rect -1255 -988 -1249 988
rect -1215 -988 -1209 988
rect -1255 -1000 -1209 -988
rect -947 988 -901 1000
rect -947 -988 -941 988
rect -907 -988 -901 988
rect -947 -1000 -901 -988
rect -639 988 -593 1000
rect -639 -988 -633 988
rect -599 -988 -593 988
rect -639 -1000 -593 -988
rect -331 988 -285 1000
rect -331 -988 -325 988
rect -291 -988 -285 988
rect -331 -1000 -285 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 285 988 331 1000
rect 285 -988 291 988
rect 325 -988 331 988
rect 285 -1000 331 -988
rect 593 988 639 1000
rect 593 -988 599 988
rect 633 -988 639 988
rect 593 -1000 639 -988
rect 901 988 947 1000
rect 901 -988 907 988
rect 941 -988 947 988
rect 901 -1000 947 -988
rect 1209 988 1255 1000
rect 1209 -988 1215 988
rect 1249 -988 1255 988
rect 1209 -1000 1255 -988
rect 1517 988 1563 1000
rect 1517 -988 1523 988
rect 1557 -988 1563 988
rect 1517 -1000 1563 -988
rect 1825 988 1871 1000
rect 1825 -988 1831 988
rect 1865 -988 1871 988
rect 1825 -1000 1871 -988
rect 2133 988 2179 1000
rect 2133 -988 2139 988
rect 2173 -988 2179 988
rect 2133 -1000 2179 -988
rect 2441 988 2487 1000
rect 2441 -988 2447 988
rect 2481 -988 2487 988
rect 2441 -1000 2487 -988
rect -2431 -1047 -2189 -1041
rect -2431 -1081 -2419 -1047
rect -2201 -1081 -2189 -1047
rect -2431 -1087 -2189 -1081
rect -2123 -1047 -1881 -1041
rect -2123 -1081 -2111 -1047
rect -1893 -1081 -1881 -1047
rect -2123 -1087 -1881 -1081
rect -1815 -1047 -1573 -1041
rect -1815 -1081 -1803 -1047
rect -1585 -1081 -1573 -1047
rect -1815 -1087 -1573 -1081
rect -1507 -1047 -1265 -1041
rect -1507 -1081 -1495 -1047
rect -1277 -1081 -1265 -1047
rect -1507 -1087 -1265 -1081
rect -1199 -1047 -957 -1041
rect -1199 -1081 -1187 -1047
rect -969 -1081 -957 -1047
rect -1199 -1087 -957 -1081
rect -891 -1047 -649 -1041
rect -891 -1081 -879 -1047
rect -661 -1081 -649 -1047
rect -891 -1087 -649 -1081
rect -583 -1047 -341 -1041
rect -583 -1081 -571 -1047
rect -353 -1081 -341 -1047
rect -583 -1087 -341 -1081
rect -275 -1047 -33 -1041
rect -275 -1081 -263 -1047
rect -45 -1081 -33 -1047
rect -275 -1087 -33 -1081
rect 33 -1047 275 -1041
rect 33 -1081 45 -1047
rect 263 -1081 275 -1047
rect 33 -1087 275 -1081
rect 341 -1047 583 -1041
rect 341 -1081 353 -1047
rect 571 -1081 583 -1047
rect 341 -1087 583 -1081
rect 649 -1047 891 -1041
rect 649 -1081 661 -1047
rect 879 -1081 891 -1047
rect 649 -1087 891 -1081
rect 957 -1047 1199 -1041
rect 957 -1081 969 -1047
rect 1187 -1081 1199 -1047
rect 957 -1087 1199 -1081
rect 1265 -1047 1507 -1041
rect 1265 -1081 1277 -1047
rect 1495 -1081 1507 -1047
rect 1265 -1087 1507 -1081
rect 1573 -1047 1815 -1041
rect 1573 -1081 1585 -1047
rect 1803 -1081 1815 -1047
rect 1573 -1087 1815 -1081
rect 1881 -1047 2123 -1041
rect 1881 -1081 1893 -1047
rect 2111 -1081 2123 -1047
rect 1881 -1087 2123 -1081
rect 2189 -1047 2431 -1041
rect 2189 -1081 2201 -1047
rect 2419 -1081 2431 -1047
rect 2189 -1087 2431 -1081
<< properties >>
string FIXED_BBOX -2598 -1202 2598 1202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 1.25 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
