magic
tech sky130A
magscale 1 2
timestamp 1770026962
<< nwell >>
rect -34200 -50400 -18400 -50100
rect -34200 -55100 -29800 -50400
rect -22400 -50700 -18400 -50400
rect -22400 -52800 -21700 -50700
rect -18800 -52800 -18400 -50700
rect -34200 -56080 -30200 -55100
rect -34200 -59800 -33800 -56080
rect -30900 -59800 -30200 -56080
rect -34200 -60100 -30200 -59800
rect -22400 -56080 -18400 -52800
rect -22400 -59800 -21700 -56080
rect -18800 -59800 -18400 -56080
rect -22400 -60100 -18400 -59800
rect -34200 -60200 -18400 -60100
<< pwell >>
rect -33800 -59800 -30900 -56080
rect -21700 -59800 -18800 -56100
<< mvpdiff >>
rect -32380 -54620 -32340 -54580
<< nsubdiff >>
rect -34100 -50240 -18500 -50200
rect -34100 -50360 -33900 -50240
rect -18700 -50360 -18500 -50240
rect -34100 -50400 -18500 -50360
rect -34100 -50440 -33900 -50400
rect -34100 -59820 -34060 -50440
rect -33940 -59820 -33900 -50440
rect -30800 -50440 -30600 -50400
rect -34100 -59900 -33900 -59820
rect -30800 -59820 -30760 -50440
rect -30640 -59820 -30600 -50440
rect -30300 -50500 -22300 -50400
rect -22000 -50460 -21800 -50400
rect -30800 -59900 -30600 -59820
rect -22000 -59840 -21960 -50460
rect -21840 -59840 -21800 -50460
rect -22000 -59900 -21800 -59840
rect -18700 -50460 -18500 -50400
rect -18700 -59840 -18660 -50460
rect -18540 -59840 -18500 -50460
rect -18700 -59900 -18500 -59840
rect -34100 -59920 -18500 -59900
rect -34100 -59940 -22580 -59920
rect -34100 -60060 -33900 -59940
rect -30820 -60060 -30600 -59940
rect -30060 -60040 -22580 -59940
rect -22040 -60040 -21800 -59920
rect -18700 -60040 -18500 -59920
rect -30060 -60060 -18500 -60040
rect -34100 -60100 -18500 -60060
<< nsubdiffcont >>
rect -33900 -50360 -18700 -50240
rect -34060 -59820 -33940 -50440
rect -30760 -59820 -30640 -50440
rect -21960 -59840 -21840 -50460
rect -18660 -59840 -18540 -50460
rect -33900 -60060 -30820 -59940
rect -30600 -60060 -30060 -59940
rect -22580 -60040 -22040 -59920
rect -21800 -60040 -18700 -59920
<< locali >>
rect -34100 -50240 -18500 -50200
rect -34100 -50360 -33900 -50240
rect -18700 -50360 -18500 -50240
rect -34100 -50400 -18500 -50360
rect -34100 -50440 -30600 -50400
rect -34100 -59820 -34060 -50440
rect -33940 -50700 -30760 -50440
rect -33940 -53000 -33700 -50700
rect -33320 -52800 -33200 -50700
rect -32700 -52800 -32580 -50700
rect -32100 -52800 -31980 -50700
rect -31480 -52800 -31360 -50700
rect -31000 -53000 -30760 -50700
rect -33940 -53660 -30760 -53000
rect -33940 -55000 -32740 -53660
rect -31980 -55000 -30760 -53660
rect -33940 -55600 -30760 -55000
rect -33940 -59820 -33900 -55600
rect -33800 -56120 -30900 -56100
rect -33800 -56220 -32560 -56120
rect -32460 -56220 -32400 -56120
rect -32300 -56220 -32240 -56120
rect -32140 -56220 -30900 -56120
rect -33800 -57120 -30900 -56220
rect -33800 -58924 -33139 -57120
rect -32760 -58740 -32620 -57120
rect -32140 -58740 -32000 -57120
rect -31640 -58924 -30900 -57120
rect -33800 -59320 -30900 -58924
rect -33800 -59420 -33780 -59320
rect -33680 -59420 -33640 -59320
rect -33540 -59420 -33500 -59320
rect -33400 -59420 -33360 -59320
rect -33260 -59420 -33220 -59320
rect -33120 -59420 -33080 -59320
rect -32980 -59420 -32940 -59320
rect -32840 -59420 -32800 -59320
rect -32700 -59420 -32660 -59320
rect -32560 -59420 -32520 -59320
rect -32420 -59420 -32380 -59320
rect -32280 -59420 -32240 -59320
rect -32140 -59420 -32100 -59320
rect -32000 -59420 -31960 -59320
rect -31860 -59420 -31820 -59320
rect -31720 -59420 -31680 -59320
rect -31580 -59420 -31540 -59320
rect -31440 -59420 -31400 -59320
rect -31300 -59420 -31260 -59320
rect -31160 -59420 -31120 -59320
rect -31020 -59420 -30900 -59320
rect -33800 -59500 -30900 -59420
rect -33800 -59600 -33780 -59500
rect -33680 -59600 -33640 -59500
rect -33540 -59600 -33500 -59500
rect -33400 -59600 -33360 -59500
rect -33260 -59600 -33220 -59500
rect -33120 -59600 -33080 -59500
rect -32980 -59600 -32940 -59500
rect -32840 -59600 -32800 -59500
rect -32700 -59600 -32660 -59500
rect -32560 -59600 -32520 -59500
rect -32420 -59600 -32380 -59500
rect -32280 -59600 -32240 -59500
rect -32140 -59600 -32100 -59500
rect -32000 -59600 -31960 -59500
rect -31860 -59600 -31820 -59500
rect -31720 -59600 -31680 -59500
rect -31580 -59600 -31540 -59500
rect -31440 -59600 -31400 -59500
rect -31300 -59600 -31260 -59500
rect -31160 -59600 -31120 -59500
rect -31020 -59600 -30900 -59500
rect -33800 -59680 -30900 -59600
rect -33800 -59780 -33780 -59680
rect -33680 -59780 -33640 -59680
rect -33540 -59780 -33500 -59680
rect -33400 -59780 -33360 -59680
rect -33260 -59780 -33220 -59680
rect -33120 -59780 -33080 -59680
rect -32980 -59780 -32940 -59680
rect -32840 -59780 -32800 -59680
rect -32700 -59780 -32660 -59680
rect -32560 -59780 -32520 -59680
rect -32420 -59780 -32380 -59680
rect -32280 -59780 -32240 -59680
rect -32140 -59780 -32100 -59680
rect -32000 -59780 -31960 -59680
rect -31860 -59780 -31820 -59680
rect -31720 -59780 -31680 -59680
rect -31580 -59780 -31540 -59680
rect -31440 -59780 -31400 -59680
rect -31300 -59780 -31260 -59680
rect -31160 -59780 -31120 -59680
rect -31020 -59780 -30900 -59680
rect -33800 -59800 -30900 -59780
rect -34100 -59900 -33900 -59820
rect -30800 -59820 -30760 -55600
rect -30640 -59820 -30600 -50440
rect -30320 -50500 -22300 -50400
rect -22000 -50460 -18500 -50400
rect -29960 -59300 -29480 -53540
rect -23160 -59300 -22680 -53540
rect -29960 -59320 -29240 -59300
rect -29960 -59420 -29940 -59320
rect -29840 -59420 -29800 -59320
rect -29700 -59420 -29660 -59320
rect -29560 -59420 -29520 -59320
rect -29420 -59420 -29380 -59320
rect -29280 -59420 -29240 -59320
rect -29960 -59500 -29240 -59420
rect -29960 -59600 -29940 -59500
rect -29840 -59600 -29800 -59500
rect -29700 -59600 -29660 -59500
rect -29560 -59600 -29520 -59500
rect -29420 -59600 -29240 -59500
rect -29960 -59680 -29240 -59600
rect -23400 -59320 -22680 -59300
rect -23400 -59420 -23360 -59320
rect -23260 -59420 -23220 -59320
rect -23120 -59420 -23080 -59320
rect -22980 -59420 -22940 -59320
rect -22840 -59420 -22800 -59320
rect -22700 -59420 -22680 -59320
rect -23400 -59500 -22680 -59420
rect -23400 -59600 -23360 -59500
rect -23260 -59600 -23220 -59500
rect -23120 -59600 -23080 -59500
rect -22980 -59600 -22940 -59500
rect -22840 -59600 -22800 -59500
rect -22700 -59600 -22680 -59500
rect -23400 -59680 -22680 -59600
rect -29960 -59780 -29940 -59680
rect -29840 -59780 -29800 -59680
rect -29700 -59780 -29660 -59680
rect -29560 -59780 -29520 -59680
rect -29420 -59780 -23360 -59680
rect -23260 -59780 -23220 -59680
rect -23120 -59780 -23080 -59680
rect -22980 -59780 -22940 -59680
rect -22840 -59780 -22800 -59680
rect -22700 -59780 -22680 -59680
rect -29960 -59800 -22680 -59780
rect -30800 -59900 -30600 -59820
rect -22000 -59840 -21960 -50460
rect -21840 -50700 -18660 -50460
rect -21840 -53000 -21600 -50700
rect -21220 -52800 -21100 -50700
rect -20620 -52800 -20500 -50700
rect -19980 -52800 -19860 -50700
rect -19380 -52800 -19260 -50700
rect -18900 -53000 -18660 -50700
rect -21840 -53680 -18660 -53000
rect -21840 -55000 -20700 -53680
rect -19970 -55000 -18660 -53680
rect -21840 -55591 -18660 -55000
rect -21840 -59840 -21800 -55591
rect -21700 -56120 -18800 -56100
rect -21700 -56220 -20540 -56120
rect -20440 -56220 -20380 -56120
rect -20280 -56220 -20220 -56120
rect -20120 -56220 -18800 -56120
rect -21700 -57120 -18800 -56220
rect -21700 -58928 -21036 -57120
rect -20660 -58740 -20520 -57120
rect -20040 -58740 -19900 -57120
rect -19537 -58928 -18800 -57120
rect -21700 -59320 -18800 -58928
rect -21700 -59420 -21580 -59320
rect -21480 -59420 -21440 -59320
rect -21340 -59420 -21300 -59320
rect -21200 -59420 -21160 -59320
rect -21060 -59420 -21020 -59320
rect -20920 -59420 -20880 -59320
rect -20780 -59420 -20740 -59320
rect -20640 -59420 -20600 -59320
rect -20500 -59420 -20460 -59320
rect -20360 -59420 -20320 -59320
rect -20220 -59420 -20180 -59320
rect -20080 -59420 -20040 -59320
rect -19940 -59420 -19900 -59320
rect -19800 -59420 -19760 -59320
rect -19660 -59420 -19620 -59320
rect -19520 -59420 -19480 -59320
rect -19380 -59420 -19340 -59320
rect -19240 -59420 -19200 -59320
rect -19100 -59420 -19060 -59320
rect -18960 -59420 -18920 -59320
rect -18820 -59420 -18800 -59320
rect -21700 -59500 -18800 -59420
rect -21700 -59600 -21580 -59500
rect -21480 -59600 -21440 -59500
rect -21340 -59600 -21300 -59500
rect -21200 -59600 -21160 -59500
rect -21060 -59600 -21020 -59500
rect -20920 -59600 -20880 -59500
rect -20780 -59600 -20740 -59500
rect -20640 -59600 -20600 -59500
rect -20500 -59600 -20460 -59500
rect -20360 -59600 -20320 -59500
rect -20220 -59600 -20180 -59500
rect -20080 -59600 -20040 -59500
rect -19940 -59600 -19900 -59500
rect -19800 -59600 -19760 -59500
rect -19660 -59600 -19620 -59500
rect -19520 -59600 -19480 -59500
rect -19380 -59600 -19340 -59500
rect -19240 -59600 -19200 -59500
rect -19100 -59600 -19060 -59500
rect -18960 -59600 -18920 -59500
rect -18820 -59600 -18800 -59500
rect -21700 -59680 -18800 -59600
rect -21700 -59780 -21580 -59680
rect -21480 -59780 -21440 -59680
rect -21340 -59780 -21300 -59680
rect -21200 -59780 -21160 -59680
rect -21060 -59780 -21020 -59680
rect -20920 -59780 -20880 -59680
rect -20780 -59780 -20740 -59680
rect -20640 -59780 -20600 -59680
rect -20500 -59780 -20460 -59680
rect -20360 -59780 -20320 -59680
rect -20220 -59780 -20180 -59680
rect -20080 -59780 -20040 -59680
rect -19940 -59780 -19900 -59680
rect -19800 -59780 -19760 -59680
rect -19660 -59780 -19620 -59680
rect -19520 -59780 -19480 -59680
rect -19380 -59780 -19340 -59680
rect -19240 -59780 -19200 -59680
rect -19100 -59780 -19060 -59680
rect -18960 -59780 -18920 -59680
rect -18820 -59780 -18800 -59680
rect -21700 -59800 -18800 -59780
rect -22000 -59900 -21800 -59840
rect -18700 -59840 -18660 -55591
rect -18540 -59840 -18500 -50460
rect -18700 -59900 -18500 -59840
rect -34100 -59920 -18500 -59900
rect -34100 -59940 -22580 -59920
rect -34100 -60060 -33900 -59940
rect -30820 -60060 -30600 -59940
rect -30060 -60040 -22580 -59940
rect -22040 -60040 -21800 -59920
rect -18700 -60040 -18500 -59920
rect -30060 -60060 -18500 -60040
rect -34100 -60100 -18500 -60060
<< viali >>
rect -32560 -56220 -32460 -56120
rect -32400 -56220 -32300 -56120
rect -32240 -56220 -32140 -56120
rect -33780 -59420 -33680 -59320
rect -33640 -59420 -33540 -59320
rect -33500 -59420 -33400 -59320
rect -33360 -59420 -33260 -59320
rect -33220 -59420 -33120 -59320
rect -33080 -59420 -32980 -59320
rect -32940 -59420 -32840 -59320
rect -32800 -59420 -32700 -59320
rect -32660 -59420 -32560 -59320
rect -32520 -59420 -32420 -59320
rect -32380 -59420 -32280 -59320
rect -32240 -59420 -32140 -59320
rect -32100 -59420 -32000 -59320
rect -31960 -59420 -31860 -59320
rect -31820 -59420 -31720 -59320
rect -31680 -59420 -31580 -59320
rect -31540 -59420 -31440 -59320
rect -31400 -59420 -31300 -59320
rect -31260 -59420 -31160 -59320
rect -31120 -59420 -31020 -59320
rect -33780 -59600 -33680 -59500
rect -33640 -59600 -33540 -59500
rect -33500 -59600 -33400 -59500
rect -33360 -59600 -33260 -59500
rect -33220 -59600 -33120 -59500
rect -33080 -59600 -32980 -59500
rect -32940 -59600 -32840 -59500
rect -32800 -59600 -32700 -59500
rect -32660 -59600 -32560 -59500
rect -32520 -59600 -32420 -59500
rect -32380 -59600 -32280 -59500
rect -32240 -59600 -32140 -59500
rect -32100 -59600 -32000 -59500
rect -31960 -59600 -31860 -59500
rect -31820 -59600 -31720 -59500
rect -31680 -59600 -31580 -59500
rect -31540 -59600 -31440 -59500
rect -31400 -59600 -31300 -59500
rect -31260 -59600 -31160 -59500
rect -31120 -59600 -31020 -59500
rect -33780 -59780 -33680 -59680
rect -33640 -59780 -33540 -59680
rect -33500 -59780 -33400 -59680
rect -33360 -59780 -33260 -59680
rect -33220 -59780 -33120 -59680
rect -33080 -59780 -32980 -59680
rect -32940 -59780 -32840 -59680
rect -32800 -59780 -32700 -59680
rect -32660 -59780 -32560 -59680
rect -32520 -59780 -32420 -59680
rect -32380 -59780 -32280 -59680
rect -32240 -59780 -32140 -59680
rect -32100 -59780 -32000 -59680
rect -31960 -59780 -31860 -59680
rect -31820 -59780 -31720 -59680
rect -31680 -59780 -31580 -59680
rect -31540 -59780 -31440 -59680
rect -31400 -59780 -31300 -59680
rect -31260 -59780 -31160 -59680
rect -31120 -59780 -31020 -59680
rect -29940 -59420 -29840 -59320
rect -29800 -59420 -29700 -59320
rect -29660 -59420 -29560 -59320
rect -29520 -59420 -29420 -59320
rect -29380 -59420 -29280 -59320
rect -29940 -59600 -29840 -59500
rect -29800 -59600 -29700 -59500
rect -29660 -59600 -29560 -59500
rect -29520 -59600 -29420 -59500
rect -23360 -59420 -23260 -59320
rect -23220 -59420 -23120 -59320
rect -23080 -59420 -22980 -59320
rect -22940 -59420 -22840 -59320
rect -22800 -59420 -22700 -59320
rect -23360 -59600 -23260 -59500
rect -23220 -59600 -23120 -59500
rect -23080 -59600 -22980 -59500
rect -22940 -59600 -22840 -59500
rect -22800 -59600 -22700 -59500
rect -29940 -59780 -29840 -59680
rect -29800 -59780 -29700 -59680
rect -29660 -59780 -29560 -59680
rect -29520 -59780 -29420 -59680
rect -23360 -59780 -23260 -59680
rect -23220 -59780 -23120 -59680
rect -23080 -59780 -22980 -59680
rect -22940 -59780 -22840 -59680
rect -22800 -59780 -22700 -59680
rect -20540 -56220 -20440 -56120
rect -20380 -56220 -20280 -56120
rect -20220 -56220 -20120 -56120
rect -21580 -59420 -21480 -59320
rect -21440 -59420 -21340 -59320
rect -21300 -59420 -21200 -59320
rect -21160 -59420 -21060 -59320
rect -21020 -59420 -20920 -59320
rect -20880 -59420 -20780 -59320
rect -20740 -59420 -20640 -59320
rect -20600 -59420 -20500 -59320
rect -20460 -59420 -20360 -59320
rect -20320 -59420 -20220 -59320
rect -20180 -59420 -20080 -59320
rect -20040 -59420 -19940 -59320
rect -19900 -59420 -19800 -59320
rect -19760 -59420 -19660 -59320
rect -19620 -59420 -19520 -59320
rect -19480 -59420 -19380 -59320
rect -19340 -59420 -19240 -59320
rect -19200 -59420 -19100 -59320
rect -19060 -59420 -18960 -59320
rect -18920 -59420 -18820 -59320
rect -21580 -59600 -21480 -59500
rect -21440 -59600 -21340 -59500
rect -21300 -59600 -21200 -59500
rect -21160 -59600 -21060 -59500
rect -21020 -59600 -20920 -59500
rect -20880 -59600 -20780 -59500
rect -20740 -59600 -20640 -59500
rect -20600 -59600 -20500 -59500
rect -20460 -59600 -20360 -59500
rect -20320 -59600 -20220 -59500
rect -20180 -59600 -20080 -59500
rect -20040 -59600 -19940 -59500
rect -19900 -59600 -19800 -59500
rect -19760 -59600 -19660 -59500
rect -19620 -59600 -19520 -59500
rect -19480 -59600 -19380 -59500
rect -19340 -59600 -19240 -59500
rect -19200 -59600 -19100 -59500
rect -19060 -59600 -18960 -59500
rect -18920 -59600 -18820 -59500
rect -21580 -59780 -21480 -59680
rect -21440 -59780 -21340 -59680
rect -21300 -59780 -21200 -59680
rect -21160 -59780 -21060 -59680
rect -21020 -59780 -20920 -59680
rect -20880 -59780 -20780 -59680
rect -20740 -59780 -20640 -59680
rect -20600 -59780 -20500 -59680
rect -20460 -59780 -20360 -59680
rect -20320 -59780 -20220 -59680
rect -20180 -59780 -20080 -59680
rect -20040 -59780 -19940 -59680
rect -19900 -59780 -19800 -59680
rect -19760 -59780 -19660 -59680
rect -19620 -59780 -19520 -59680
rect -19480 -59780 -19380 -59680
rect -19340 -59780 -19240 -59680
rect -19200 -59780 -19100 -59680
rect -19060 -59780 -18960 -59680
rect -18920 -59780 -18820 -59680
<< metal1 >>
rect -33620 -51720 -33500 -51700
rect -33620 -51800 -33600 -51720
rect -33520 -51800 -33500 -51720
rect -33620 -51940 -33500 -51800
rect -33620 -52020 -33600 -51940
rect -33520 -52020 -33500 -51940
rect -33620 -52040 -33500 -52020
rect -33020 -51720 -32900 -51700
rect -33020 -51800 -33000 -51720
rect -32920 -51800 -32900 -51720
rect -33020 -51940 -32900 -51800
rect -33020 -52020 -33000 -51940
rect -32920 -52020 -32900 -51940
rect -33020 -52040 -32900 -52020
rect -32400 -51720 -32280 -51700
rect -32400 -51800 -32380 -51720
rect -32300 -51800 -32280 -51720
rect -32400 -51940 -32280 -51800
rect -32400 -52020 -32380 -51940
rect -32300 -52020 -32280 -51940
rect -32400 -52040 -32280 -52020
rect -31780 -51720 -31660 -51700
rect -31780 -51800 -31760 -51720
rect -31680 -51800 -31660 -51720
rect -31780 -51940 -31660 -51800
rect -31780 -52020 -31760 -51940
rect -31680 -52020 -31660 -51940
rect -31780 -52040 -31660 -52020
rect -31180 -51720 -31060 -51700
rect -31180 -51800 -31160 -51720
rect -31080 -51800 -31060 -51720
rect -31180 -51940 -31060 -51800
rect -31180 -52020 -31160 -51940
rect -31080 -52020 -31060 -51940
rect -31180 -52040 -31060 -52020
rect -21540 -51720 -21420 -51700
rect -21540 -51800 -21520 -51720
rect -21440 -51800 -21420 -51720
rect -21540 -51940 -21420 -51800
rect -21540 -52020 -21520 -51940
rect -21440 -52020 -21420 -51940
rect -21540 -52040 -21420 -52020
rect -20920 -51720 -20800 -51700
rect -20920 -51800 -20900 -51720
rect -20820 -51800 -20800 -51720
rect -20920 -51940 -20800 -51800
rect -20920 -52020 -20900 -51940
rect -20820 -52020 -20800 -51940
rect -20920 -52040 -20800 -52020
rect -20300 -51720 -20180 -51700
rect -20300 -51800 -20280 -51720
rect -20200 -51800 -20180 -51720
rect -20300 -51940 -20180 -51800
rect -20300 -52020 -20280 -51940
rect -20200 -52020 -20180 -51940
rect -20300 -52040 -20180 -52020
rect -19680 -51720 -19560 -51700
rect -19680 -51800 -19660 -51720
rect -19580 -51800 -19560 -51720
rect -19680 -51940 -19560 -51800
rect -19680 -52020 -19660 -51940
rect -19580 -52020 -19560 -51940
rect -19680 -52040 -19560 -52020
rect -19080 -51720 -18960 -51700
rect -19080 -51800 -19060 -51720
rect -18980 -51800 -18960 -51720
rect -19080 -51940 -18960 -51800
rect -19080 -52020 -19060 -51940
rect -18980 -52020 -18960 -51940
rect -19080 -52040 -18960 -52020
rect -33540 -52900 -31140 -52880
rect -21440 -52900 -19040 -52860
rect -33600 -52920 -30500 -52900
rect -33600 -52980 -30680 -52920
rect -30620 -52980 -30580 -52920
rect -30520 -52980 -30500 -52920
rect -33600 -53020 -30500 -52980
rect -33600 -53080 -30680 -53020
rect -30620 -53080 -30580 -53020
rect -30520 -53080 -30500 -53020
rect -33600 -53100 -30500 -53080
rect -22100 -52920 -19000 -52900
rect -22100 -52980 -22080 -52920
rect -22020 -52980 -21980 -52920
rect -21920 -52980 -19000 -52920
rect -22100 -53020 -19000 -52980
rect -22100 -53080 -22080 -53020
rect -22020 -53080 -21980 -53020
rect -21920 -53080 -19000 -53020
rect -22100 -53100 -19000 -53080
rect -32660 -53920 -32520 -53900
rect -32660 -53980 -32620 -53920
rect -32560 -53980 -32520 -53920
rect -32660 -54020 -32520 -53980
rect -32660 -54080 -32620 -54020
rect -32560 -54080 -32520 -54020
rect -32660 -54100 -32520 -54080
rect -32180 -53920 -32040 -53900
rect -32180 -53980 -32140 -53920
rect -32080 -53980 -32040 -53920
rect -32180 -54020 -32040 -53980
rect -32180 -54080 -32140 -54020
rect -32080 -54080 -32040 -54020
rect -32180 -54100 -32040 -54080
rect -20620 -53920 -20520 -53900
rect -20620 -53980 -20600 -53920
rect -20540 -53980 -20520 -53920
rect -20620 -54020 -20520 -53980
rect -20620 -54080 -20600 -54020
rect -20540 -54080 -20520 -54020
rect -20620 -54100 -20520 -54080
rect -20140 -53920 -20040 -53900
rect -20140 -53980 -20120 -53920
rect -20060 -53980 -20040 -53920
rect -20140 -54020 -20040 -53980
rect -20140 -54080 -20120 -54020
rect -20060 -54080 -20040 -54020
rect -20140 -54100 -20040 -54080
rect -33900 -54320 -33600 -54300
rect -33900 -54380 -33880 -54320
rect -33820 -54380 -33680 -54320
rect -33620 -54380 -33600 -54320
rect -33900 -54480 -33600 -54380
rect -33900 -54540 -33880 -54480
rect -33820 -54500 -33600 -54480
rect -33820 -54540 -33680 -54500
rect -33900 -54560 -33680 -54540
rect -33620 -54560 -33600 -54500
rect -33900 -54640 -33600 -54560
rect -33900 -54700 -33880 -54640
rect -33820 -54700 -33780 -54640
rect -33720 -54700 -33680 -54640
rect -33620 -54700 -33600 -54640
rect -33900 -54720 -33600 -54700
rect -32500 -54320 -32200 -54300
rect -32500 -54380 -32480 -54320
rect -32420 -54380 -32280 -54320
rect -32220 -54380 -32200 -54320
rect -32500 -54420 -32200 -54380
rect -32500 -54480 -32480 -54420
rect -32420 -54480 -32280 -54420
rect -32220 -54480 -32200 -54420
rect -32500 -54540 -32200 -54480
rect -32500 -54600 -32480 -54540
rect -32420 -54600 -32280 -54540
rect -32220 -54600 -32200 -54540
rect -32500 -54640 -32200 -54600
rect -32500 -54700 -32480 -54640
rect -32420 -54700 -32280 -54640
rect -32220 -54700 -32200 -54640
rect -32500 -54720 -32200 -54700
rect -20480 -54320 -20180 -54300
rect -20480 -54380 -20460 -54320
rect -20400 -54380 -20260 -54320
rect -20200 -54380 -20180 -54320
rect -20480 -54420 -20180 -54380
rect -20480 -54480 -20460 -54420
rect -20400 -54480 -20260 -54420
rect -20200 -54480 -20180 -54420
rect -20480 -54540 -20180 -54480
rect -20480 -54600 -20460 -54540
rect -20400 -54600 -20260 -54540
rect -20200 -54600 -20180 -54540
rect -20480 -54640 -20180 -54600
rect -20480 -54700 -20460 -54640
rect -20400 -54700 -20260 -54640
rect -20200 -54700 -20180 -54640
rect -20480 -54720 -20180 -54700
rect -19000 -54320 -18700 -54300
rect -19000 -54380 -18980 -54320
rect -18920 -54380 -18880 -54320
rect -18820 -54380 -18780 -54320
rect -18720 -54380 -18700 -54320
rect -19000 -54500 -18700 -54380
rect -19000 -54560 -18980 -54500
rect -18920 -54560 -18880 -54500
rect -18820 -54560 -18780 -54500
rect -18720 -54560 -18700 -54500
rect -19000 -54640 -18700 -54560
rect -19000 -54700 -18980 -54640
rect -18920 -54700 -18880 -54640
rect -18820 -54700 -18780 -54640
rect -18720 -54700 -18700 -54640
rect -19000 -54720 -18700 -54700
rect -32580 -56120 -32120 -54840
rect -23300 -55160 -23100 -55140
rect -23300 -55220 -23280 -55160
rect -23220 -55220 -23180 -55160
rect -23120 -55220 -23100 -55160
rect -23300 -55260 -23100 -55220
rect -23300 -55320 -23280 -55260
rect -23220 -55320 -23180 -55260
rect -23120 -55320 -23100 -55260
rect -23300 -55340 -23100 -55320
rect -29500 -55660 -29300 -55640
rect -29500 -55720 -29480 -55660
rect -29420 -55720 -29380 -55660
rect -29320 -55720 -29300 -55660
rect -29500 -55760 -29300 -55720
rect -29500 -55820 -29480 -55760
rect -29420 -55820 -29380 -55760
rect -29320 -55820 -29300 -55760
rect -29500 -55840 -29300 -55820
rect -32580 -56220 -32560 -56120
rect -32460 -56220 -32400 -56120
rect -32300 -56220 -32240 -56120
rect -32140 -56220 -32120 -56120
rect -32580 -56240 -32120 -56220
rect -20560 -56120 -20100 -54860
rect -20560 -56220 -20540 -56120
rect -20440 -56220 -20380 -56120
rect -20280 -56220 -20220 -56120
rect -20120 -56220 -20100 -56120
rect -20560 -56240 -20100 -56220
rect -33060 -57880 -32940 -57860
rect -33060 -57960 -33040 -57880
rect -32960 -57960 -32940 -57880
rect -33060 -58100 -32940 -57960
rect -33060 -58180 -33040 -58100
rect -32960 -58180 -32940 -58100
rect -33060 -58200 -32940 -58180
rect -32440 -57880 -32320 -57860
rect -32440 -57960 -32420 -57880
rect -32340 -57960 -32320 -57880
rect -32440 -58100 -32320 -57960
rect -32440 -58180 -32420 -58100
rect -32340 -58180 -32320 -58100
rect -32440 -58200 -32320 -58180
rect -31820 -57880 -31700 -57860
rect -31820 -57960 -31800 -57880
rect -31720 -57960 -31700 -57880
rect -31820 -58100 -31700 -57960
rect -31820 -58180 -31800 -58100
rect -31720 -58180 -31700 -58100
rect -31820 -58200 -31700 -58180
rect -20960 -57880 -20820 -57860
rect -20960 -57960 -20940 -57880
rect -20860 -57960 -20820 -57880
rect -20960 -58100 -20820 -57960
rect -20960 -58180 -20940 -58100
rect -20860 -58180 -20820 -58100
rect -20960 -58200 -20820 -58180
rect -20360 -57880 -20220 -57860
rect -20360 -57960 -20320 -57880
rect -20240 -57960 -20220 -57880
rect -20360 -58100 -20220 -57960
rect -20360 -58180 -20320 -58100
rect -20240 -58180 -20220 -58100
rect -20360 -58200 -20220 -58180
rect -19760 -57880 -19620 -57860
rect -19760 -57960 -19740 -57880
rect -19660 -57960 -19620 -57880
rect -19760 -58100 -19620 -57960
rect -19760 -58180 -19740 -58100
rect -19660 -58180 -19620 -58100
rect -19760 -58200 -19620 -58180
rect -32980 -59240 -31780 -58780
rect -20880 -59240 -19680 -58780
rect -33800 -59320 -29200 -59300
rect -33800 -59420 -33780 -59320
rect -33680 -59420 -33640 -59320
rect -33540 -59420 -33500 -59320
rect -33400 -59420 -33360 -59320
rect -33260 -59420 -33220 -59320
rect -33120 -59420 -33080 -59320
rect -32980 -59420 -32940 -59320
rect -32840 -59420 -32800 -59320
rect -32700 -59420 -32660 -59320
rect -32560 -59420 -32520 -59320
rect -32420 -59420 -32380 -59320
rect -32280 -59420 -32240 -59320
rect -32140 -59420 -32100 -59320
rect -32000 -59420 -31960 -59320
rect -31860 -59420 -31820 -59320
rect -31720 -59420 -31680 -59320
rect -31580 -59420 -31540 -59320
rect -31440 -59420 -31400 -59320
rect -31300 -59420 -31260 -59320
rect -31160 -59420 -31120 -59320
rect -31020 -59420 -29940 -59320
rect -29840 -59420 -29800 -59320
rect -29700 -59420 -29660 -59320
rect -29560 -59420 -29520 -59320
rect -29420 -59420 -29380 -59320
rect -29280 -59420 -29200 -59320
rect -33800 -59500 -29200 -59420
rect -33800 -59600 -33780 -59500
rect -33680 -59600 -33640 -59500
rect -33540 -59600 -33500 -59500
rect -33400 -59600 -33360 -59500
rect -33260 -59600 -33220 -59500
rect -33120 -59600 -33080 -59500
rect -32980 -59600 -32940 -59500
rect -32840 -59600 -32800 -59500
rect -32700 -59600 -32660 -59500
rect -32560 -59600 -32520 -59500
rect -32420 -59600 -32380 -59500
rect -32280 -59600 -32240 -59500
rect -32140 -59600 -32100 -59500
rect -32000 -59600 -31960 -59500
rect -31860 -59600 -31820 -59500
rect -31720 -59600 -31680 -59500
rect -31580 -59600 -31540 -59500
rect -31440 -59600 -31400 -59500
rect -31300 -59600 -31260 -59500
rect -31160 -59600 -31120 -59500
rect -31020 -59600 -29940 -59500
rect -29840 -59600 -29800 -59500
rect -29700 -59600 -29660 -59500
rect -29560 -59600 -29520 -59500
rect -29420 -59600 -29200 -59500
rect -33800 -59680 -29200 -59600
rect -33800 -59780 -33780 -59680
rect -33680 -59780 -33640 -59680
rect -33540 -59780 -33500 -59680
rect -33400 -59780 -33360 -59680
rect -33260 -59780 -33220 -59680
rect -33120 -59780 -33080 -59680
rect -32980 -59780 -32940 -59680
rect -32840 -59780 -32800 -59680
rect -32700 -59780 -32660 -59680
rect -32560 -59780 -32520 -59680
rect -32420 -59780 -32380 -59680
rect -32280 -59780 -32240 -59680
rect -32140 -59780 -32100 -59680
rect -32000 -59780 -31960 -59680
rect -31860 -59780 -31820 -59680
rect -31720 -59780 -31680 -59680
rect -31580 -59780 -31540 -59680
rect -31440 -59780 -31400 -59680
rect -31300 -59780 -31260 -59680
rect -31160 -59780 -31120 -59680
rect -31020 -59780 -29940 -59680
rect -29840 -59780 -29800 -59680
rect -29700 -59780 -29660 -59680
rect -29560 -59780 -29520 -59680
rect -29420 -59780 -29200 -59680
rect -33800 -59800 -29200 -59780
rect -23400 -59320 -18800 -59300
rect -23400 -59420 -23360 -59320
rect -23260 -59420 -23220 -59320
rect -23120 -59420 -23080 -59320
rect -22980 -59420 -22940 -59320
rect -22840 -59420 -22800 -59320
rect -22700 -59420 -21580 -59320
rect -21480 -59420 -21440 -59320
rect -21340 -59420 -21300 -59320
rect -21200 -59420 -21160 -59320
rect -21060 -59420 -21020 -59320
rect -20920 -59420 -20880 -59320
rect -20780 -59420 -20740 -59320
rect -20640 -59420 -20600 -59320
rect -20500 -59420 -20460 -59320
rect -20360 -59420 -20320 -59320
rect -20220 -59420 -20180 -59320
rect -20080 -59420 -20040 -59320
rect -19940 -59420 -19900 -59320
rect -19800 -59420 -19760 -59320
rect -19660 -59420 -19620 -59320
rect -19520 -59420 -19480 -59320
rect -19380 -59420 -19340 -59320
rect -19240 -59420 -19200 -59320
rect -19100 -59420 -19060 -59320
rect -18960 -59420 -18920 -59320
rect -18820 -59420 -18800 -59320
rect -23400 -59500 -18800 -59420
rect -23400 -59600 -23360 -59500
rect -23260 -59600 -23220 -59500
rect -23120 -59600 -23080 -59500
rect -22980 -59600 -22940 -59500
rect -22840 -59600 -22800 -59500
rect -22700 -59600 -21580 -59500
rect -21480 -59600 -21440 -59500
rect -21340 -59600 -21300 -59500
rect -21200 -59600 -21160 -59500
rect -21060 -59600 -21020 -59500
rect -20920 -59600 -20880 -59500
rect -20780 -59600 -20740 -59500
rect -20640 -59600 -20600 -59500
rect -20500 -59600 -20460 -59500
rect -20360 -59600 -20320 -59500
rect -20220 -59600 -20180 -59500
rect -20080 -59600 -20040 -59500
rect -19940 -59600 -19900 -59500
rect -19800 -59600 -19760 -59500
rect -19660 -59600 -19620 -59500
rect -19520 -59600 -19480 -59500
rect -19380 -59600 -19340 -59500
rect -19240 -59600 -19200 -59500
rect -19100 -59600 -19060 -59500
rect -18960 -59600 -18920 -59500
rect -18820 -59600 -18800 -59500
rect -23400 -59680 -18800 -59600
rect -23400 -59780 -23360 -59680
rect -23260 -59780 -23220 -59680
rect -23120 -59780 -23080 -59680
rect -22980 -59780 -22940 -59680
rect -22840 -59780 -22800 -59680
rect -22700 -59780 -21580 -59680
rect -21480 -59780 -21440 -59680
rect -21340 -59780 -21300 -59680
rect -21200 -59780 -21160 -59680
rect -21060 -59780 -21020 -59680
rect -20920 -59780 -20880 -59680
rect -20780 -59780 -20740 -59680
rect -20640 -59780 -20600 -59680
rect -20500 -59780 -20460 -59680
rect -20360 -59780 -20320 -59680
rect -20220 -59780 -20180 -59680
rect -20080 -59780 -20040 -59680
rect -19940 -59780 -19900 -59680
rect -19800 -59780 -19760 -59680
rect -19660 -59780 -19620 -59680
rect -19520 -59780 -19480 -59680
rect -19380 -59780 -19340 -59680
rect -19240 -59780 -19200 -59680
rect -19100 -59780 -19060 -59680
rect -18960 -59780 -18920 -59680
rect -18820 -59780 -18800 -59680
rect -23400 -59800 -18800 -59780
<< via1 >>
rect -33600 -51800 -33520 -51720
rect -33600 -52020 -33520 -51940
rect -33000 -51800 -32920 -51720
rect -33000 -52020 -32920 -51940
rect -32380 -51800 -32300 -51720
rect -32380 -52020 -32300 -51940
rect -31760 -51800 -31680 -51720
rect -31760 -52020 -31680 -51940
rect -31160 -51800 -31080 -51720
rect -31160 -52020 -31080 -51940
rect -21520 -51800 -21440 -51720
rect -21520 -52020 -21440 -51940
rect -20900 -51800 -20820 -51720
rect -20900 -52020 -20820 -51940
rect -20280 -51800 -20200 -51720
rect -20280 -52020 -20200 -51940
rect -19660 -51800 -19580 -51720
rect -19660 -52020 -19580 -51940
rect -19060 -51800 -18980 -51720
rect -19060 -52020 -18980 -51940
rect -30680 -52980 -30620 -52920
rect -30580 -52980 -30520 -52920
rect -30680 -53080 -30620 -53020
rect -30580 -53080 -30520 -53020
rect -22080 -52980 -22020 -52920
rect -21980 -52980 -21920 -52920
rect -22080 -53080 -22020 -53020
rect -21980 -53080 -21920 -53020
rect -32620 -53980 -32560 -53920
rect -32620 -54080 -32560 -54020
rect -32140 -53980 -32080 -53920
rect -32140 -54080 -32080 -54020
rect -20600 -53980 -20540 -53920
rect -20600 -54080 -20540 -54020
rect -20120 -53980 -20060 -53920
rect -20120 -54080 -20060 -54020
rect -33880 -54380 -33820 -54320
rect -33680 -54380 -33620 -54320
rect -33880 -54540 -33820 -54480
rect -33680 -54560 -33620 -54500
rect -33880 -54700 -33820 -54640
rect -33780 -54700 -33720 -54640
rect -33680 -54700 -33620 -54640
rect -32480 -54380 -32420 -54320
rect -32280 -54380 -32220 -54320
rect -32480 -54480 -32420 -54420
rect -32280 -54480 -32220 -54420
rect -32480 -54600 -32420 -54540
rect -32280 -54600 -32220 -54540
rect -32480 -54700 -32420 -54640
rect -32280 -54700 -32220 -54640
rect -20460 -54380 -20400 -54320
rect -20260 -54380 -20200 -54320
rect -20460 -54480 -20400 -54420
rect -20260 -54480 -20200 -54420
rect -20460 -54600 -20400 -54540
rect -20260 -54600 -20200 -54540
rect -20460 -54700 -20400 -54640
rect -20260 -54700 -20200 -54640
rect -18980 -54380 -18920 -54320
rect -18880 -54380 -18820 -54320
rect -18780 -54380 -18720 -54320
rect -18980 -54560 -18920 -54500
rect -18880 -54560 -18820 -54500
rect -18780 -54560 -18720 -54500
rect -18980 -54700 -18920 -54640
rect -18880 -54700 -18820 -54640
rect -18780 -54700 -18720 -54640
rect -23280 -55220 -23220 -55160
rect -23180 -55220 -23120 -55160
rect -23280 -55320 -23220 -55260
rect -23180 -55320 -23120 -55260
rect -29480 -55720 -29420 -55660
rect -29380 -55720 -29320 -55660
rect -29480 -55820 -29420 -55760
rect -29380 -55820 -29320 -55760
rect -33040 -57960 -32960 -57880
rect -33040 -58180 -32960 -58100
rect -32420 -57960 -32340 -57880
rect -32420 -58180 -32340 -58100
rect -31800 -57960 -31720 -57880
rect -31800 -58180 -31720 -58100
rect -20940 -57960 -20860 -57880
rect -20940 -58180 -20860 -58100
rect -20320 -57960 -20240 -57880
rect -20320 -58180 -20240 -58100
rect -19740 -57960 -19660 -57880
rect -19740 -58180 -19660 -58100
<< metal2 >>
rect -33960 -51720 -30760 -51700
rect -33960 -51800 -33600 -51720
rect -33520 -51800 -33000 -51720
rect -32920 -51800 -32380 -51720
rect -32300 -51800 -31760 -51720
rect -31680 -51800 -31160 -51720
rect -31080 -51800 -30760 -51720
rect -33960 -51940 -30760 -51800
rect -33960 -52020 -33600 -51940
rect -33520 -52020 -33000 -51940
rect -32920 -52020 -32380 -51940
rect -32300 -52020 -31760 -51940
rect -31680 -52020 -31160 -51940
rect -31080 -52020 -30760 -51940
rect -33960 -52040 -30760 -52020
rect -21860 -51720 -18660 -51700
rect -21860 -51800 -21520 -51720
rect -21440 -51800 -20900 -51720
rect -20820 -51800 -20280 -51720
rect -20200 -51800 -19660 -51720
rect -19580 -51800 -19060 -51720
rect -18980 -51800 -18660 -51720
rect -21860 -51940 -18660 -51800
rect -21860 -52020 -21520 -51940
rect -21440 -52020 -20900 -51940
rect -20820 -52020 -20280 -51940
rect -20200 -52020 -19660 -51940
rect -19580 -52020 -19060 -51940
rect -18980 -52020 -18660 -51940
rect -21860 -52040 -18660 -52020
rect -33900 -54320 -33600 -52040
rect -30700 -52920 -30500 -52900
rect -30700 -52980 -30680 -52920
rect -30620 -52980 -30580 -52920
rect -30520 -52980 -30500 -52920
rect -30700 -53020 -30500 -52980
rect -30700 -53080 -30680 -53020
rect -30620 -53080 -30580 -53020
rect -30520 -53080 -30500 -53020
rect -30700 -53100 -30500 -53080
rect -22100 -52920 -21900 -52900
rect -22100 -52980 -22080 -52920
rect -22020 -52980 -21980 -52920
rect -21920 -52980 -21900 -52920
rect -22100 -53020 -21900 -52980
rect -22100 -53080 -22080 -53020
rect -22020 -53080 -21980 -53020
rect -21920 -53080 -21900 -53020
rect -22100 -53100 -21900 -53080
rect -32660 -53920 -32520 -53900
rect -32660 -53980 -32620 -53920
rect -32560 -53980 -32520 -53920
rect -32660 -54020 -32520 -53980
rect -32660 -54080 -32620 -54020
rect -32560 -54080 -32520 -54020
rect -32660 -54100 -32520 -54080
rect -32180 -53920 -32040 -53900
rect -32180 -53980 -32140 -53920
rect -32080 -53980 -32040 -53920
rect -32180 -54020 -32040 -53980
rect -32180 -54080 -32140 -54020
rect -32080 -54080 -32040 -54020
rect -32180 -54100 -32040 -54080
rect -20620 -53920 -20520 -53900
rect -20620 -53980 -20600 -53920
rect -20540 -53980 -20520 -53920
rect -20620 -54020 -20520 -53980
rect -20620 -54080 -20600 -54020
rect -20540 -54080 -20520 -54020
rect -20620 -54100 -20520 -54080
rect -20140 -53920 -20040 -53900
rect -20140 -53980 -20120 -53920
rect -20060 -53980 -20040 -53920
rect -20140 -54020 -20040 -53980
rect -20140 -54080 -20120 -54020
rect -20060 -54080 -20040 -54020
rect -20140 -54100 -20040 -54080
rect -33900 -54380 -33880 -54320
rect -33820 -54380 -33780 -54320
rect -33720 -54380 -33680 -54320
rect -33620 -54380 -33600 -54320
rect -33900 -54480 -33600 -54380
rect -33900 -54560 -33880 -54480
rect -33820 -54500 -33600 -54480
rect -33820 -54560 -33780 -54500
rect -33720 -54560 -33680 -54500
rect -33620 -54560 -33600 -54500
rect -33900 -54640 -33600 -54560
rect -33900 -54700 -33880 -54640
rect -33820 -54700 -33780 -54640
rect -33720 -54700 -33680 -54640
rect -33620 -54700 -33600 -54640
rect -33900 -57860 -33600 -54700
rect -32500 -54320 -32200 -54300
rect -32500 -54380 -32480 -54320
rect -32420 -54380 -32380 -54320
rect -32320 -54380 -32280 -54320
rect -32220 -54380 -32200 -54320
rect -32500 -54420 -32200 -54380
rect -32500 -54480 -32480 -54420
rect -32420 -54480 -32380 -54420
rect -32320 -54480 -32280 -54420
rect -32220 -54480 -32200 -54420
rect -32500 -54540 -32200 -54480
rect -32500 -54600 -32480 -54540
rect -32420 -54600 -32380 -54540
rect -32320 -54600 -32280 -54540
rect -32220 -54600 -32200 -54540
rect -32500 -54640 -32200 -54600
rect -32500 -54700 -32480 -54640
rect -32420 -54700 -32380 -54640
rect -32320 -54700 -32280 -54640
rect -32220 -54700 -32200 -54640
rect -32500 -54720 -32200 -54700
rect -20480 -54320 -20180 -54300
rect -20480 -54380 -20460 -54320
rect -20400 -54380 -20360 -54320
rect -20300 -54380 -20260 -54320
rect -20200 -54380 -20180 -54320
rect -20480 -54420 -20180 -54380
rect -20480 -54480 -20460 -54420
rect -20400 -54480 -20360 -54420
rect -20300 -54480 -20260 -54420
rect -20200 -54480 -20180 -54420
rect -20480 -54540 -20180 -54480
rect -20480 -54600 -20460 -54540
rect -20400 -54600 -20360 -54540
rect -20300 -54600 -20260 -54540
rect -20200 -54600 -20180 -54540
rect -20480 -54640 -20180 -54600
rect -20480 -54700 -20460 -54640
rect -20400 -54700 -20360 -54640
rect -20300 -54700 -20260 -54640
rect -20200 -54700 -20180 -54640
rect -20480 -54720 -20180 -54700
rect -19000 -54320 -18700 -52040
rect -19000 -54380 -18980 -54320
rect -18920 -54380 -18880 -54320
rect -18820 -54380 -18780 -54320
rect -18720 -54380 -18700 -54320
rect -19000 -54480 -18700 -54380
rect -19000 -54560 -18980 -54480
rect -18920 -54500 -18780 -54480
rect -18920 -54560 -18880 -54500
rect -18820 -54560 -18780 -54500
rect -18720 -54560 -18700 -54480
rect -19000 -54640 -18700 -54560
rect -19000 -54700 -18980 -54640
rect -18920 -54700 -18880 -54640
rect -18820 -54700 -18780 -54640
rect -18720 -54700 -18700 -54640
rect -23300 -55160 -23100 -55140
rect -23300 -55220 -23280 -55160
rect -23220 -55220 -23180 -55160
rect -23120 -55220 -23100 -55160
rect -23300 -55260 -23100 -55220
rect -23300 -55320 -23280 -55260
rect -23220 -55320 -23180 -55260
rect -23120 -55320 -23100 -55260
rect -23300 -55340 -23100 -55320
rect -30140 -55380 -29900 -55360
rect -30140 -55460 -30120 -55380
rect -30040 -55460 -30000 -55380
rect -29920 -55460 -29900 -55380
rect -30140 -55540 -29900 -55460
rect -30140 -55620 -30120 -55540
rect -30040 -55620 -30000 -55540
rect -29920 -55620 -29900 -55540
rect -30140 -55640 -29900 -55620
rect -22740 -55380 -22500 -55360
rect -22740 -55460 -22720 -55380
rect -22640 -55460 -22600 -55380
rect -22520 -55460 -22500 -55380
rect -22740 -55540 -22500 -55460
rect -22740 -55620 -22720 -55540
rect -22640 -55620 -22600 -55540
rect -22520 -55620 -22500 -55540
rect -22740 -55640 -22500 -55620
rect -29500 -55660 -29300 -55640
rect -29500 -55720 -29480 -55660
rect -29420 -55720 -29380 -55660
rect -29320 -55720 -29300 -55660
rect -29500 -55760 -29300 -55720
rect -29500 -55820 -29480 -55760
rect -29420 -55820 -29380 -55760
rect -29320 -55820 -29300 -55760
rect -29500 -55840 -29300 -55820
rect -19000 -57860 -18700 -54700
rect -33940 -57880 -30740 -57860
rect -33940 -57960 -33040 -57880
rect -32960 -57960 -32420 -57880
rect -32340 -57960 -31800 -57880
rect -31720 -57960 -30740 -57880
rect -33940 -58100 -30740 -57960
rect -33940 -58180 -33040 -58100
rect -32960 -58180 -32420 -58100
rect -32340 -58180 -31800 -58100
rect -31720 -58180 -30740 -58100
rect -33940 -58200 -30740 -58180
rect -21820 -57880 -18620 -57860
rect -21820 -57960 -20940 -57880
rect -20860 -57960 -20320 -57880
rect -20240 -57960 -19740 -57880
rect -19660 -57960 -18620 -57880
rect -21820 -58100 -18620 -57960
rect -21820 -58180 -20940 -58100
rect -20860 -58180 -20320 -58100
rect -20240 -58180 -19740 -58100
rect -19660 -58180 -18620 -58100
rect -21820 -58200 -18620 -58180
rect -29620 -59000 -29320 -58580
rect -32980 -59240 -29320 -59000
rect -23320 -59000 -23020 -58580
rect -23320 -59240 -19660 -59000
<< via2 >>
rect -30680 -52980 -30620 -52920
rect -30580 -52980 -30520 -52920
rect -30680 -53080 -30620 -53020
rect -30580 -53080 -30520 -53020
rect -22080 -52980 -22020 -52920
rect -21980 -52980 -21920 -52920
rect -22080 -53080 -22020 -53020
rect -21980 -53080 -21920 -53020
rect -32620 -53980 -32560 -53920
rect -32620 -54080 -32560 -54020
rect -32140 -53980 -32080 -53920
rect -32140 -54080 -32080 -54020
rect -20600 -53980 -20540 -53920
rect -20600 -54080 -20540 -54020
rect -20120 -53980 -20060 -53920
rect -20120 -54080 -20060 -54020
rect -33880 -54380 -33820 -54320
rect -33780 -54380 -33720 -54320
rect -33680 -54380 -33620 -54320
rect -33880 -54540 -33820 -54500
rect -33880 -54560 -33820 -54540
rect -33780 -54560 -33720 -54500
rect -33680 -54560 -33620 -54500
rect -33880 -54700 -33820 -54640
rect -33780 -54700 -33720 -54640
rect -33680 -54700 -33620 -54640
rect -32380 -54380 -32320 -54320
rect -32380 -54480 -32320 -54420
rect -32380 -54600 -32320 -54540
rect -32380 -54700 -32320 -54640
rect -20360 -54380 -20300 -54320
rect -20360 -54480 -20300 -54420
rect -20360 -54600 -20300 -54540
rect -20360 -54700 -20300 -54640
rect -18980 -54380 -18920 -54320
rect -18880 -54380 -18820 -54320
rect -18780 -54380 -18720 -54320
rect -18980 -54500 -18920 -54480
rect -18780 -54500 -18720 -54480
rect -18980 -54540 -18920 -54500
rect -18880 -54560 -18820 -54500
rect -18780 -54540 -18720 -54500
rect -18980 -54700 -18920 -54640
rect -18880 -54700 -18820 -54640
rect -18780 -54700 -18720 -54640
rect -23280 -55220 -23220 -55160
rect -23180 -55220 -23120 -55160
rect -23280 -55320 -23220 -55260
rect -23180 -55320 -23120 -55260
rect -30120 -55460 -30040 -55380
rect -30000 -55460 -29920 -55380
rect -30120 -55620 -30040 -55540
rect -30000 -55620 -29920 -55540
rect -22720 -55460 -22640 -55380
rect -22600 -55460 -22520 -55380
rect -22720 -55620 -22640 -55540
rect -22600 -55620 -22520 -55540
rect -29480 -55720 -29420 -55660
rect -29380 -55720 -29320 -55660
rect -29480 -55820 -29420 -55760
rect -29380 -55820 -29320 -55760
<< metal3 >>
rect -30700 -52920 -30500 -52900
rect -30700 -53080 -30680 -52920
rect -30520 -53080 -30500 -52920
rect -30700 -53100 -30500 -53080
rect -22100 -52920 -21900 -52900
rect -22100 -53080 -22080 -52920
rect -21920 -53080 -21900 -52920
rect -22100 -53100 -21900 -53080
rect -34700 -53300 -34500 -53280
rect -34700 -53380 -34640 -53300
rect -34560 -53380 -34500 -53300
rect -34700 -53400 -34500 -53380
rect -34700 -53480 -34640 -53400
rect -34560 -53480 -34500 -53400
rect -34700 -53900 -34500 -53480
rect -18100 -53300 -17900 -53280
rect -18100 -53380 -18040 -53300
rect -17960 -53380 -17900 -53300
rect -18100 -53400 -17900 -53380
rect -18100 -53480 -18040 -53400
rect -17960 -53480 -17900 -53400
rect -18100 -53900 -17900 -53480
rect -34700 -53920 -31900 -53900
rect -34700 -53980 -32620 -53920
rect -32560 -53980 -32140 -53920
rect -32080 -53980 -31900 -53920
rect -34700 -54020 -31900 -53980
rect -34700 -54080 -32620 -54020
rect -32560 -54080 -32140 -54020
rect -32080 -54080 -31900 -54020
rect -34700 -54100 -31900 -54080
rect -20800 -53920 -17900 -53900
rect -20800 -53980 -20600 -53920
rect -20540 -53980 -20120 -53920
rect -20060 -53980 -17900 -53920
rect -20800 -54020 -17900 -53980
rect -20800 -54080 -20600 -54020
rect -20540 -54080 -20120 -54020
rect -20060 -54080 -17900 -54020
rect -20800 -54100 -17900 -54080
rect -33900 -54320 -33600 -54300
rect -33900 -54400 -33880 -54320
rect -33800 -54380 -33780 -54320
rect -33720 -54380 -33700 -54320
rect -33800 -54400 -33700 -54380
rect -33620 -54400 -33600 -54320
rect -33900 -54480 -33600 -54400
rect -33900 -54560 -33880 -54480
rect -33800 -54500 -33700 -54480
rect -33800 -54560 -33780 -54500
rect -33720 -54560 -33700 -54500
rect -33620 -54560 -33600 -54480
rect -33900 -54620 -33600 -54560
rect -33900 -54700 -33880 -54620
rect -33800 -54640 -33700 -54620
rect -33800 -54700 -33780 -54640
rect -33720 -54700 -33700 -54640
rect -33620 -54700 -33600 -54620
rect -33900 -54720 -33600 -54700
rect -32500 -54320 -32200 -54300
rect -32500 -54400 -32480 -54320
rect -32400 -54380 -32380 -54320
rect -32320 -54380 -32300 -54320
rect -32400 -54400 -32300 -54380
rect -32220 -54400 -32200 -54320
rect -32500 -54420 -32200 -54400
rect -32500 -54500 -32480 -54420
rect -32400 -54480 -32380 -54420
rect -32320 -54480 -32300 -54420
rect -32400 -54500 -32300 -54480
rect -32220 -54500 -32200 -54420
rect -32500 -54520 -32200 -54500
rect -32500 -54600 -32480 -54520
rect -32400 -54540 -32300 -54520
rect -32400 -54600 -32380 -54540
rect -32320 -54600 -32300 -54540
rect -32220 -54600 -32200 -54520
rect -32500 -54620 -32200 -54600
rect -32500 -54700 -32480 -54620
rect -32400 -54640 -32300 -54620
rect -32400 -54700 -32380 -54640
rect -32320 -54700 -32300 -54640
rect -32220 -54700 -32200 -54620
rect -32500 -54720 -32200 -54700
rect -20480 -54320 -20180 -54300
rect -20480 -54400 -20460 -54320
rect -20380 -54380 -20360 -54320
rect -20300 -54380 -20280 -54320
rect -20380 -54400 -20280 -54380
rect -20200 -54400 -20180 -54320
rect -20480 -54420 -20180 -54400
rect -20480 -54500 -20460 -54420
rect -20380 -54480 -20360 -54420
rect -20300 -54480 -20280 -54420
rect -20380 -54500 -20280 -54480
rect -20200 -54500 -20180 -54420
rect -20480 -54520 -20180 -54500
rect -20480 -54600 -20460 -54520
rect -20380 -54540 -20280 -54520
rect -20380 -54600 -20360 -54540
rect -20300 -54600 -20280 -54540
rect -20200 -54600 -20180 -54520
rect -20480 -54620 -20180 -54600
rect -20480 -54700 -20460 -54620
rect -20380 -54640 -20280 -54620
rect -20380 -54700 -20360 -54640
rect -20300 -54700 -20280 -54640
rect -20200 -54700 -20180 -54620
rect -20480 -54720 -20180 -54700
rect -19000 -54320 -18700 -54300
rect -19000 -54400 -18980 -54320
rect -18900 -54380 -18880 -54320
rect -18820 -54380 -18800 -54320
rect -18900 -54400 -18800 -54380
rect -18720 -54400 -18700 -54320
rect -19000 -54480 -18700 -54400
rect -19000 -54560 -18980 -54480
rect -18900 -54500 -18800 -54480
rect -18900 -54560 -18880 -54500
rect -18820 -54560 -18800 -54500
rect -18720 -54560 -18700 -54480
rect -19000 -54620 -18700 -54560
rect -19000 -54700 -18980 -54620
rect -18900 -54640 -18800 -54620
rect -18900 -54700 -18880 -54640
rect -18820 -54700 -18800 -54640
rect -18720 -54700 -18700 -54620
rect -19000 -54720 -18700 -54700
rect -23300 -55160 -23100 -55140
rect -23300 -55320 -23280 -55160
rect -23120 -55320 -23100 -55160
rect -23300 -55340 -23100 -55320
rect -30140 -55380 -29900 -55360
rect -30140 -55460 -30120 -55380
rect -30040 -55460 -30000 -55380
rect -29920 -55460 -29900 -55380
rect -30140 -55540 -29900 -55460
rect -30140 -55620 -30120 -55540
rect -30040 -55620 -30000 -55540
rect -29920 -55620 -29900 -55540
rect -30140 -55640 -29900 -55620
rect -22740 -55380 -22500 -55360
rect -22740 -55460 -22720 -55380
rect -22640 -55460 -22600 -55380
rect -22520 -55460 -22500 -55380
rect -22740 -55540 -22500 -55460
rect -22740 -55620 -22720 -55540
rect -22640 -55620 -22600 -55540
rect -22520 -55620 -22500 -55540
rect -22740 -55640 -22500 -55620
rect -29500 -55660 -29300 -55640
rect -29500 -55820 -29480 -55660
rect -29320 -55820 -29300 -55660
rect -29500 -55840 -29300 -55820
<< via3 >>
rect -30680 -52980 -30620 -52920
rect -30620 -52980 -30580 -52920
rect -30580 -52980 -30520 -52920
rect -30680 -53020 -30520 -52980
rect -30680 -53080 -30620 -53020
rect -30620 -53080 -30580 -53020
rect -30580 -53080 -30520 -53020
rect -22080 -52980 -22020 -52920
rect -22020 -52980 -21980 -52920
rect -21980 -52980 -21920 -52920
rect -22080 -53020 -21920 -52980
rect -22080 -53080 -22020 -53020
rect -22020 -53080 -21980 -53020
rect -21980 -53080 -21920 -53020
rect -34640 -53380 -34560 -53300
rect -34640 -53480 -34560 -53400
rect -18040 -53380 -17960 -53300
rect -18040 -53480 -17960 -53400
rect -33880 -54380 -33820 -54320
rect -33820 -54380 -33800 -54320
rect -33700 -54380 -33680 -54320
rect -33680 -54380 -33620 -54320
rect -33880 -54400 -33800 -54380
rect -33700 -54400 -33620 -54380
rect -33880 -54500 -33800 -54480
rect -33700 -54500 -33620 -54480
rect -33880 -54560 -33820 -54500
rect -33820 -54560 -33800 -54500
rect -33700 -54560 -33680 -54500
rect -33680 -54560 -33620 -54500
rect -33880 -54640 -33800 -54620
rect -33700 -54640 -33620 -54620
rect -33880 -54700 -33820 -54640
rect -33820 -54700 -33800 -54640
rect -33700 -54700 -33680 -54640
rect -33680 -54700 -33620 -54640
rect -32480 -54400 -32400 -54320
rect -32300 -54400 -32220 -54320
rect -32480 -54500 -32400 -54420
rect -32300 -54500 -32220 -54420
rect -32480 -54600 -32400 -54520
rect -32300 -54600 -32220 -54520
rect -32480 -54700 -32400 -54620
rect -32300 -54700 -32220 -54620
rect -20460 -54400 -20380 -54320
rect -20280 -54400 -20200 -54320
rect -20460 -54500 -20380 -54420
rect -20280 -54500 -20200 -54420
rect -20460 -54600 -20380 -54520
rect -20280 -54600 -20200 -54520
rect -20460 -54700 -20380 -54620
rect -20280 -54700 -20200 -54620
rect -18980 -54380 -18920 -54320
rect -18920 -54380 -18900 -54320
rect -18800 -54380 -18780 -54320
rect -18780 -54380 -18720 -54320
rect -18980 -54400 -18900 -54380
rect -18800 -54400 -18720 -54380
rect -18980 -54540 -18920 -54480
rect -18920 -54540 -18900 -54480
rect -18980 -54560 -18900 -54540
rect -18800 -54540 -18780 -54480
rect -18780 -54540 -18720 -54480
rect -18800 -54560 -18720 -54540
rect -18980 -54640 -18900 -54620
rect -18800 -54640 -18720 -54620
rect -18980 -54700 -18920 -54640
rect -18920 -54700 -18900 -54640
rect -18800 -54700 -18780 -54640
rect -18780 -54700 -18720 -54640
rect -23280 -55220 -23220 -55160
rect -23220 -55220 -23180 -55160
rect -23180 -55220 -23120 -55160
rect -23280 -55260 -23120 -55220
rect -23280 -55320 -23220 -55260
rect -23220 -55320 -23180 -55260
rect -23180 -55320 -23120 -55260
rect -30120 -55460 -30040 -55380
rect -30000 -55460 -29920 -55380
rect -30120 -55620 -30040 -55540
rect -30000 -55620 -29920 -55540
rect -22720 -55460 -22640 -55380
rect -22600 -55460 -22520 -55380
rect -22720 -55620 -22640 -55540
rect -22600 -55620 -22520 -55540
rect -29480 -55720 -29420 -55660
rect -29420 -55720 -29380 -55660
rect -29380 -55720 -29320 -55660
rect -29480 -55760 -29320 -55720
rect -29480 -55820 -29420 -55760
rect -29420 -55820 -29380 -55760
rect -29380 -55820 -29320 -55760
<< metal4 >>
rect -47800 -47300 -47400 -47100
rect -5000 -47300 -4600 -47100
rect -47800 -51300 -47600 -47300
rect -47800 -51500 -34500 -51300
rect -34700 -53300 -34500 -51500
rect -34700 -53380 -34640 -53300
rect -34560 -53380 -34500 -53300
rect -34700 -53400 -34500 -53380
rect -34700 -53480 -34640 -53400
rect -34560 -53480 -34500 -53400
rect -34700 -53500 -34500 -53480
rect -30700 -52920 -30500 -49900
rect -30700 -53080 -30680 -52920
rect -30520 -53080 -30500 -52920
rect -33900 -54320 -33600 -54300
rect -33900 -54700 -33880 -54320
rect -33800 -54380 -33700 -54320
rect -33800 -54700 -33700 -54640
rect -33620 -54700 -33600 -54320
rect -33900 -54720 -33600 -54700
rect -32500 -54320 -32200 -54300
rect -32500 -54700 -32480 -54320
rect -32400 -54380 -32300 -54320
rect -32400 -54700 -32300 -54640
rect -32220 -54700 -32200 -54320
rect -32500 -54720 -32200 -54700
rect -30700 -55400 -30500 -53080
rect -22100 -52920 -21900 -49900
rect -4800 -51300 -4600 -47300
rect -22100 -53080 -22080 -52920
rect -21920 -53080 -21900 -52920
rect -30140 -55380 -29900 -55360
rect -30140 -55400 -30120 -55380
rect -30700 -55460 -30120 -55400
rect -30040 -55460 -30000 -55380
rect -29920 -55400 -29900 -55380
rect -29920 -55460 -29600 -55400
rect -30700 -55540 -29600 -55460
rect -30700 -55600 -30120 -55540
rect -30140 -55620 -30120 -55600
rect -30040 -55620 -30000 -55540
rect -29920 -55600 -29600 -55540
rect -29920 -55620 -29900 -55600
rect -30140 -55640 -29900 -55620
rect -29500 -55660 -29300 -55100
rect -29500 -55820 -29480 -55660
rect -29320 -55820 -29300 -55660
rect -29500 -60600 -29300 -55820
rect -23300 -55160 -23100 -55100
rect -23300 -55320 -23280 -55160
rect -23120 -55320 -23100 -55160
rect -23300 -60600 -23100 -55320
rect -22740 -55380 -22500 -55360
rect -22740 -55400 -22720 -55380
rect -23000 -55460 -22720 -55400
rect -22640 -55460 -22600 -55380
rect -22520 -55400 -22500 -55380
rect -22100 -55400 -21900 -53080
rect -18100 -51500 -4600 -51300
rect -18100 -53300 -17900 -51500
rect -18100 -53380 -18040 -53300
rect -17960 -53380 -17900 -53300
rect -18100 -53400 -17900 -53380
rect -18100 -53480 -18040 -53400
rect -17960 -53480 -17900 -53400
rect -18100 -53500 -17900 -53480
rect -20480 -54320 -20180 -54300
rect -20480 -54700 -20460 -54320
rect -20380 -54380 -20280 -54320
rect -20380 -54700 -20280 -54640
rect -20200 -54700 -20180 -54320
rect -20480 -54720 -20180 -54700
rect -19000 -54320 -18700 -54300
rect -19000 -54700 -18980 -54320
rect -18900 -54380 -18800 -54320
rect -18900 -54700 -18800 -54640
rect -18720 -54700 -18700 -54320
rect -19000 -54720 -18700 -54700
rect -22520 -55460 -21900 -55400
rect -23000 -55540 -21900 -55460
rect -23000 -55600 -22720 -55540
rect -22740 -55620 -22720 -55600
rect -22640 -55620 -22600 -55540
rect -22520 -55600 -21900 -55540
rect -22520 -55620 -22500 -55600
rect -22740 -55640 -22500 -55620
<< via4 >>
rect -33880 -54400 -33800 -54380
rect -33800 -54400 -33700 -54380
rect -33700 -54400 -33620 -54380
rect -33880 -54480 -33620 -54400
rect -33880 -54560 -33800 -54480
rect -33800 -54560 -33700 -54480
rect -33700 -54560 -33620 -54480
rect -33880 -54620 -33620 -54560
rect -33880 -54640 -33800 -54620
rect -33800 -54640 -33700 -54620
rect -33700 -54640 -33620 -54620
rect -32480 -54400 -32400 -54380
rect -32400 -54400 -32300 -54380
rect -32300 -54400 -32220 -54380
rect -32480 -54420 -32220 -54400
rect -32480 -54500 -32400 -54420
rect -32400 -54500 -32300 -54420
rect -32300 -54500 -32220 -54420
rect -32480 -54520 -32220 -54500
rect -32480 -54600 -32400 -54520
rect -32400 -54600 -32300 -54520
rect -32300 -54600 -32220 -54520
rect -32480 -54620 -32220 -54600
rect -32480 -54640 -32400 -54620
rect -32400 -54640 -32300 -54620
rect -32300 -54640 -32220 -54620
rect -20460 -54400 -20380 -54380
rect -20380 -54400 -20280 -54380
rect -20280 -54400 -20200 -54380
rect -20460 -54420 -20200 -54400
rect -20460 -54500 -20380 -54420
rect -20380 -54500 -20280 -54420
rect -20280 -54500 -20200 -54420
rect -20460 -54520 -20200 -54500
rect -20460 -54600 -20380 -54520
rect -20380 -54600 -20280 -54520
rect -20280 -54600 -20200 -54520
rect -20460 -54620 -20200 -54600
rect -20460 -54640 -20380 -54620
rect -20380 -54640 -20280 -54620
rect -20280 -54640 -20200 -54620
rect -18980 -54400 -18900 -54380
rect -18900 -54400 -18800 -54380
rect -18800 -54400 -18720 -54380
rect -18980 -54480 -18720 -54400
rect -18980 -54560 -18900 -54480
rect -18900 -54560 -18800 -54480
rect -18800 -54560 -18720 -54480
rect -18980 -54620 -18720 -54560
rect -18980 -54640 -18900 -54620
rect -18900 -54640 -18800 -54620
rect -18800 -54640 -18720 -54620
<< metal5 >>
rect -34700 -54380 -17900 -54300
rect -34700 -54640 -33880 -54380
rect -33620 -54640 -32480 -54380
rect -32220 -54640 -20460 -54380
rect -20200 -54640 -18980 -54380
rect -18720 -54640 -17900 -54380
rect -34700 -54720 -17900 -54640
use 5t-ota_top  5t-ota_top_0 /foss/designs/icdec-biomedical-pmic/xschem/error-amplifier/schematics/sub-blocks
timestamp 1770013200
transform 1 0 -31518 0 1 -55548
box 1200 -5022 9200 5200
use sky130_fd_pr__cap_mim_m3_1_S7S847  sky130_fd_pr__cap_mim_m3_1_S7S847_0
timestamp 1770023980
transform 0 1 -26220 -1 0 -47314
box -2686 -21280 2686 21280
use sky130_fd_pr__nfet_g5v0d10v5_J76LUE  sky130_fd_pr__nfet_g5v0d10v5_J76LUE_0
timestamp 1770023980
transform 1 0 -32385 0 1 -58023
box -815 -977 815 977
use sky130_fd_pr__pfet_g5v0d10v5_AP3ZHE  sky130_fd_pr__pfet_g5v0d10v5_AP3ZHE_0
timestamp 1770023980
transform 1 0 -32353 0 1 -54318
box -467 -762 467 762
use sky130_fd_pr__pfet_g5v0d10v5_D6DL9T  sky130_fd_pr__pfet_g5v0d10v5_D6DL9T_0
timestamp 1770023980
transform 1 0 -32339 0 1 -51838
box -1461 -1262 1461 1262
use sky130_fd_pr__pfet_g5v0d10v5_D6DL9T  sky130_fd_pr__pfet_g5v0d10v5_D6DL9T_1
timestamp 1770023980
transform 1 0 -20239 0 1 -51838
box -1461 -1262 1461 1262
use sky130_fd_pr__nfet_g5v0d10v5_J76LUE  XM8
timestamp 1770023980
transform 1 0 -20285 0 1 -58023
box -815 -977 815 977
use sky130_fd_pr__pfet_g5v0d10v5_AP3ZHE  XM9
timestamp 1770023980
transform 1 0 -20333 0 1 -54338
box -467 -762 467 762
<< end >>
