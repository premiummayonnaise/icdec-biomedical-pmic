magic
tech sky130A
magscale 1 2
timestamp 1769436194
<< pwell >>
rect -10311 -2258 10311 2258
<< mvnmos >>
rect -10083 -2000 -9983 2000
rect -9925 -2000 -9825 2000
rect -9767 -2000 -9667 2000
rect -9609 -2000 -9509 2000
rect -9451 -2000 -9351 2000
rect -9293 -2000 -9193 2000
rect -9135 -2000 -9035 2000
rect -8977 -2000 -8877 2000
rect -8819 -2000 -8719 2000
rect -8661 -2000 -8561 2000
rect -8503 -2000 -8403 2000
rect -8345 -2000 -8245 2000
rect -8187 -2000 -8087 2000
rect -8029 -2000 -7929 2000
rect -7871 -2000 -7771 2000
rect -7713 -2000 -7613 2000
rect -7555 -2000 -7455 2000
rect -7397 -2000 -7297 2000
rect -7239 -2000 -7139 2000
rect -7081 -2000 -6981 2000
rect -6923 -2000 -6823 2000
rect -6765 -2000 -6665 2000
rect -6607 -2000 -6507 2000
rect -6449 -2000 -6349 2000
rect -6291 -2000 -6191 2000
rect -6133 -2000 -6033 2000
rect -5975 -2000 -5875 2000
rect -5817 -2000 -5717 2000
rect -5659 -2000 -5559 2000
rect -5501 -2000 -5401 2000
rect -5343 -2000 -5243 2000
rect -5185 -2000 -5085 2000
rect -5027 -2000 -4927 2000
rect -4869 -2000 -4769 2000
rect -4711 -2000 -4611 2000
rect -4553 -2000 -4453 2000
rect -4395 -2000 -4295 2000
rect -4237 -2000 -4137 2000
rect -4079 -2000 -3979 2000
rect -3921 -2000 -3821 2000
rect -3763 -2000 -3663 2000
rect -3605 -2000 -3505 2000
rect -3447 -2000 -3347 2000
rect -3289 -2000 -3189 2000
rect -3131 -2000 -3031 2000
rect -2973 -2000 -2873 2000
rect -2815 -2000 -2715 2000
rect -2657 -2000 -2557 2000
rect -2499 -2000 -2399 2000
rect -2341 -2000 -2241 2000
rect -2183 -2000 -2083 2000
rect -2025 -2000 -1925 2000
rect -1867 -2000 -1767 2000
rect -1709 -2000 -1609 2000
rect -1551 -2000 -1451 2000
rect -1393 -2000 -1293 2000
rect -1235 -2000 -1135 2000
rect -1077 -2000 -977 2000
rect -919 -2000 -819 2000
rect -761 -2000 -661 2000
rect -603 -2000 -503 2000
rect -445 -2000 -345 2000
rect -287 -2000 -187 2000
rect -129 -2000 -29 2000
rect 29 -2000 129 2000
rect 187 -2000 287 2000
rect 345 -2000 445 2000
rect 503 -2000 603 2000
rect 661 -2000 761 2000
rect 819 -2000 919 2000
rect 977 -2000 1077 2000
rect 1135 -2000 1235 2000
rect 1293 -2000 1393 2000
rect 1451 -2000 1551 2000
rect 1609 -2000 1709 2000
rect 1767 -2000 1867 2000
rect 1925 -2000 2025 2000
rect 2083 -2000 2183 2000
rect 2241 -2000 2341 2000
rect 2399 -2000 2499 2000
rect 2557 -2000 2657 2000
rect 2715 -2000 2815 2000
rect 2873 -2000 2973 2000
rect 3031 -2000 3131 2000
rect 3189 -2000 3289 2000
rect 3347 -2000 3447 2000
rect 3505 -2000 3605 2000
rect 3663 -2000 3763 2000
rect 3821 -2000 3921 2000
rect 3979 -2000 4079 2000
rect 4137 -2000 4237 2000
rect 4295 -2000 4395 2000
rect 4453 -2000 4553 2000
rect 4611 -2000 4711 2000
rect 4769 -2000 4869 2000
rect 4927 -2000 5027 2000
rect 5085 -2000 5185 2000
rect 5243 -2000 5343 2000
rect 5401 -2000 5501 2000
rect 5559 -2000 5659 2000
rect 5717 -2000 5817 2000
rect 5875 -2000 5975 2000
rect 6033 -2000 6133 2000
rect 6191 -2000 6291 2000
rect 6349 -2000 6449 2000
rect 6507 -2000 6607 2000
rect 6665 -2000 6765 2000
rect 6823 -2000 6923 2000
rect 6981 -2000 7081 2000
rect 7139 -2000 7239 2000
rect 7297 -2000 7397 2000
rect 7455 -2000 7555 2000
rect 7613 -2000 7713 2000
rect 7771 -2000 7871 2000
rect 7929 -2000 8029 2000
rect 8087 -2000 8187 2000
rect 8245 -2000 8345 2000
rect 8403 -2000 8503 2000
rect 8561 -2000 8661 2000
rect 8719 -2000 8819 2000
rect 8877 -2000 8977 2000
rect 9035 -2000 9135 2000
rect 9193 -2000 9293 2000
rect 9351 -2000 9451 2000
rect 9509 -2000 9609 2000
rect 9667 -2000 9767 2000
rect 9825 -2000 9925 2000
rect 9983 -2000 10083 2000
<< mvndiff >>
rect -10141 1988 -10083 2000
rect -10141 -1988 -10129 1988
rect -10095 -1988 -10083 1988
rect -10141 -2000 -10083 -1988
rect -9983 1988 -9925 2000
rect -9983 -1988 -9971 1988
rect -9937 -1988 -9925 1988
rect -9983 -2000 -9925 -1988
rect -9825 1988 -9767 2000
rect -9825 -1988 -9813 1988
rect -9779 -1988 -9767 1988
rect -9825 -2000 -9767 -1988
rect -9667 1988 -9609 2000
rect -9667 -1988 -9655 1988
rect -9621 -1988 -9609 1988
rect -9667 -2000 -9609 -1988
rect -9509 1988 -9451 2000
rect -9509 -1988 -9497 1988
rect -9463 -1988 -9451 1988
rect -9509 -2000 -9451 -1988
rect -9351 1988 -9293 2000
rect -9351 -1988 -9339 1988
rect -9305 -1988 -9293 1988
rect -9351 -2000 -9293 -1988
rect -9193 1988 -9135 2000
rect -9193 -1988 -9181 1988
rect -9147 -1988 -9135 1988
rect -9193 -2000 -9135 -1988
rect -9035 1988 -8977 2000
rect -9035 -1988 -9023 1988
rect -8989 -1988 -8977 1988
rect -9035 -2000 -8977 -1988
rect -8877 1988 -8819 2000
rect -8877 -1988 -8865 1988
rect -8831 -1988 -8819 1988
rect -8877 -2000 -8819 -1988
rect -8719 1988 -8661 2000
rect -8719 -1988 -8707 1988
rect -8673 -1988 -8661 1988
rect -8719 -2000 -8661 -1988
rect -8561 1988 -8503 2000
rect -8561 -1988 -8549 1988
rect -8515 -1988 -8503 1988
rect -8561 -2000 -8503 -1988
rect -8403 1988 -8345 2000
rect -8403 -1988 -8391 1988
rect -8357 -1988 -8345 1988
rect -8403 -2000 -8345 -1988
rect -8245 1988 -8187 2000
rect -8245 -1988 -8233 1988
rect -8199 -1988 -8187 1988
rect -8245 -2000 -8187 -1988
rect -8087 1988 -8029 2000
rect -8087 -1988 -8075 1988
rect -8041 -1988 -8029 1988
rect -8087 -2000 -8029 -1988
rect -7929 1988 -7871 2000
rect -7929 -1988 -7917 1988
rect -7883 -1988 -7871 1988
rect -7929 -2000 -7871 -1988
rect -7771 1988 -7713 2000
rect -7771 -1988 -7759 1988
rect -7725 -1988 -7713 1988
rect -7771 -2000 -7713 -1988
rect -7613 1988 -7555 2000
rect -7613 -1988 -7601 1988
rect -7567 -1988 -7555 1988
rect -7613 -2000 -7555 -1988
rect -7455 1988 -7397 2000
rect -7455 -1988 -7443 1988
rect -7409 -1988 -7397 1988
rect -7455 -2000 -7397 -1988
rect -7297 1988 -7239 2000
rect -7297 -1988 -7285 1988
rect -7251 -1988 -7239 1988
rect -7297 -2000 -7239 -1988
rect -7139 1988 -7081 2000
rect -7139 -1988 -7127 1988
rect -7093 -1988 -7081 1988
rect -7139 -2000 -7081 -1988
rect -6981 1988 -6923 2000
rect -6981 -1988 -6969 1988
rect -6935 -1988 -6923 1988
rect -6981 -2000 -6923 -1988
rect -6823 1988 -6765 2000
rect -6823 -1988 -6811 1988
rect -6777 -1988 -6765 1988
rect -6823 -2000 -6765 -1988
rect -6665 1988 -6607 2000
rect -6665 -1988 -6653 1988
rect -6619 -1988 -6607 1988
rect -6665 -2000 -6607 -1988
rect -6507 1988 -6449 2000
rect -6507 -1988 -6495 1988
rect -6461 -1988 -6449 1988
rect -6507 -2000 -6449 -1988
rect -6349 1988 -6291 2000
rect -6349 -1988 -6337 1988
rect -6303 -1988 -6291 1988
rect -6349 -2000 -6291 -1988
rect -6191 1988 -6133 2000
rect -6191 -1988 -6179 1988
rect -6145 -1988 -6133 1988
rect -6191 -2000 -6133 -1988
rect -6033 1988 -5975 2000
rect -6033 -1988 -6021 1988
rect -5987 -1988 -5975 1988
rect -6033 -2000 -5975 -1988
rect -5875 1988 -5817 2000
rect -5875 -1988 -5863 1988
rect -5829 -1988 -5817 1988
rect -5875 -2000 -5817 -1988
rect -5717 1988 -5659 2000
rect -5717 -1988 -5705 1988
rect -5671 -1988 -5659 1988
rect -5717 -2000 -5659 -1988
rect -5559 1988 -5501 2000
rect -5559 -1988 -5547 1988
rect -5513 -1988 -5501 1988
rect -5559 -2000 -5501 -1988
rect -5401 1988 -5343 2000
rect -5401 -1988 -5389 1988
rect -5355 -1988 -5343 1988
rect -5401 -2000 -5343 -1988
rect -5243 1988 -5185 2000
rect -5243 -1988 -5231 1988
rect -5197 -1988 -5185 1988
rect -5243 -2000 -5185 -1988
rect -5085 1988 -5027 2000
rect -5085 -1988 -5073 1988
rect -5039 -1988 -5027 1988
rect -5085 -2000 -5027 -1988
rect -4927 1988 -4869 2000
rect -4927 -1988 -4915 1988
rect -4881 -1988 -4869 1988
rect -4927 -2000 -4869 -1988
rect -4769 1988 -4711 2000
rect -4769 -1988 -4757 1988
rect -4723 -1988 -4711 1988
rect -4769 -2000 -4711 -1988
rect -4611 1988 -4553 2000
rect -4611 -1988 -4599 1988
rect -4565 -1988 -4553 1988
rect -4611 -2000 -4553 -1988
rect -4453 1988 -4395 2000
rect -4453 -1988 -4441 1988
rect -4407 -1988 -4395 1988
rect -4453 -2000 -4395 -1988
rect -4295 1988 -4237 2000
rect -4295 -1988 -4283 1988
rect -4249 -1988 -4237 1988
rect -4295 -2000 -4237 -1988
rect -4137 1988 -4079 2000
rect -4137 -1988 -4125 1988
rect -4091 -1988 -4079 1988
rect -4137 -2000 -4079 -1988
rect -3979 1988 -3921 2000
rect -3979 -1988 -3967 1988
rect -3933 -1988 -3921 1988
rect -3979 -2000 -3921 -1988
rect -3821 1988 -3763 2000
rect -3821 -1988 -3809 1988
rect -3775 -1988 -3763 1988
rect -3821 -2000 -3763 -1988
rect -3663 1988 -3605 2000
rect -3663 -1988 -3651 1988
rect -3617 -1988 -3605 1988
rect -3663 -2000 -3605 -1988
rect -3505 1988 -3447 2000
rect -3505 -1988 -3493 1988
rect -3459 -1988 -3447 1988
rect -3505 -2000 -3447 -1988
rect -3347 1988 -3289 2000
rect -3347 -1988 -3335 1988
rect -3301 -1988 -3289 1988
rect -3347 -2000 -3289 -1988
rect -3189 1988 -3131 2000
rect -3189 -1988 -3177 1988
rect -3143 -1988 -3131 1988
rect -3189 -2000 -3131 -1988
rect -3031 1988 -2973 2000
rect -3031 -1988 -3019 1988
rect -2985 -1988 -2973 1988
rect -3031 -2000 -2973 -1988
rect -2873 1988 -2815 2000
rect -2873 -1988 -2861 1988
rect -2827 -1988 -2815 1988
rect -2873 -2000 -2815 -1988
rect -2715 1988 -2657 2000
rect -2715 -1988 -2703 1988
rect -2669 -1988 -2657 1988
rect -2715 -2000 -2657 -1988
rect -2557 1988 -2499 2000
rect -2557 -1988 -2545 1988
rect -2511 -1988 -2499 1988
rect -2557 -2000 -2499 -1988
rect -2399 1988 -2341 2000
rect -2399 -1988 -2387 1988
rect -2353 -1988 -2341 1988
rect -2399 -2000 -2341 -1988
rect -2241 1988 -2183 2000
rect -2241 -1988 -2229 1988
rect -2195 -1988 -2183 1988
rect -2241 -2000 -2183 -1988
rect -2083 1988 -2025 2000
rect -2083 -1988 -2071 1988
rect -2037 -1988 -2025 1988
rect -2083 -2000 -2025 -1988
rect -1925 1988 -1867 2000
rect -1925 -1988 -1913 1988
rect -1879 -1988 -1867 1988
rect -1925 -2000 -1867 -1988
rect -1767 1988 -1709 2000
rect -1767 -1988 -1755 1988
rect -1721 -1988 -1709 1988
rect -1767 -2000 -1709 -1988
rect -1609 1988 -1551 2000
rect -1609 -1988 -1597 1988
rect -1563 -1988 -1551 1988
rect -1609 -2000 -1551 -1988
rect -1451 1988 -1393 2000
rect -1451 -1988 -1439 1988
rect -1405 -1988 -1393 1988
rect -1451 -2000 -1393 -1988
rect -1293 1988 -1235 2000
rect -1293 -1988 -1281 1988
rect -1247 -1988 -1235 1988
rect -1293 -2000 -1235 -1988
rect -1135 1988 -1077 2000
rect -1135 -1988 -1123 1988
rect -1089 -1988 -1077 1988
rect -1135 -2000 -1077 -1988
rect -977 1988 -919 2000
rect -977 -1988 -965 1988
rect -931 -1988 -919 1988
rect -977 -2000 -919 -1988
rect -819 1988 -761 2000
rect -819 -1988 -807 1988
rect -773 -1988 -761 1988
rect -819 -2000 -761 -1988
rect -661 1988 -603 2000
rect -661 -1988 -649 1988
rect -615 -1988 -603 1988
rect -661 -2000 -603 -1988
rect -503 1988 -445 2000
rect -503 -1988 -491 1988
rect -457 -1988 -445 1988
rect -503 -2000 -445 -1988
rect -345 1988 -287 2000
rect -345 -1988 -333 1988
rect -299 -1988 -287 1988
rect -345 -2000 -287 -1988
rect -187 1988 -129 2000
rect -187 -1988 -175 1988
rect -141 -1988 -129 1988
rect -187 -2000 -129 -1988
rect -29 1988 29 2000
rect -29 -1988 -17 1988
rect 17 -1988 29 1988
rect -29 -2000 29 -1988
rect 129 1988 187 2000
rect 129 -1988 141 1988
rect 175 -1988 187 1988
rect 129 -2000 187 -1988
rect 287 1988 345 2000
rect 287 -1988 299 1988
rect 333 -1988 345 1988
rect 287 -2000 345 -1988
rect 445 1988 503 2000
rect 445 -1988 457 1988
rect 491 -1988 503 1988
rect 445 -2000 503 -1988
rect 603 1988 661 2000
rect 603 -1988 615 1988
rect 649 -1988 661 1988
rect 603 -2000 661 -1988
rect 761 1988 819 2000
rect 761 -1988 773 1988
rect 807 -1988 819 1988
rect 761 -2000 819 -1988
rect 919 1988 977 2000
rect 919 -1988 931 1988
rect 965 -1988 977 1988
rect 919 -2000 977 -1988
rect 1077 1988 1135 2000
rect 1077 -1988 1089 1988
rect 1123 -1988 1135 1988
rect 1077 -2000 1135 -1988
rect 1235 1988 1293 2000
rect 1235 -1988 1247 1988
rect 1281 -1988 1293 1988
rect 1235 -2000 1293 -1988
rect 1393 1988 1451 2000
rect 1393 -1988 1405 1988
rect 1439 -1988 1451 1988
rect 1393 -2000 1451 -1988
rect 1551 1988 1609 2000
rect 1551 -1988 1563 1988
rect 1597 -1988 1609 1988
rect 1551 -2000 1609 -1988
rect 1709 1988 1767 2000
rect 1709 -1988 1721 1988
rect 1755 -1988 1767 1988
rect 1709 -2000 1767 -1988
rect 1867 1988 1925 2000
rect 1867 -1988 1879 1988
rect 1913 -1988 1925 1988
rect 1867 -2000 1925 -1988
rect 2025 1988 2083 2000
rect 2025 -1988 2037 1988
rect 2071 -1988 2083 1988
rect 2025 -2000 2083 -1988
rect 2183 1988 2241 2000
rect 2183 -1988 2195 1988
rect 2229 -1988 2241 1988
rect 2183 -2000 2241 -1988
rect 2341 1988 2399 2000
rect 2341 -1988 2353 1988
rect 2387 -1988 2399 1988
rect 2341 -2000 2399 -1988
rect 2499 1988 2557 2000
rect 2499 -1988 2511 1988
rect 2545 -1988 2557 1988
rect 2499 -2000 2557 -1988
rect 2657 1988 2715 2000
rect 2657 -1988 2669 1988
rect 2703 -1988 2715 1988
rect 2657 -2000 2715 -1988
rect 2815 1988 2873 2000
rect 2815 -1988 2827 1988
rect 2861 -1988 2873 1988
rect 2815 -2000 2873 -1988
rect 2973 1988 3031 2000
rect 2973 -1988 2985 1988
rect 3019 -1988 3031 1988
rect 2973 -2000 3031 -1988
rect 3131 1988 3189 2000
rect 3131 -1988 3143 1988
rect 3177 -1988 3189 1988
rect 3131 -2000 3189 -1988
rect 3289 1988 3347 2000
rect 3289 -1988 3301 1988
rect 3335 -1988 3347 1988
rect 3289 -2000 3347 -1988
rect 3447 1988 3505 2000
rect 3447 -1988 3459 1988
rect 3493 -1988 3505 1988
rect 3447 -2000 3505 -1988
rect 3605 1988 3663 2000
rect 3605 -1988 3617 1988
rect 3651 -1988 3663 1988
rect 3605 -2000 3663 -1988
rect 3763 1988 3821 2000
rect 3763 -1988 3775 1988
rect 3809 -1988 3821 1988
rect 3763 -2000 3821 -1988
rect 3921 1988 3979 2000
rect 3921 -1988 3933 1988
rect 3967 -1988 3979 1988
rect 3921 -2000 3979 -1988
rect 4079 1988 4137 2000
rect 4079 -1988 4091 1988
rect 4125 -1988 4137 1988
rect 4079 -2000 4137 -1988
rect 4237 1988 4295 2000
rect 4237 -1988 4249 1988
rect 4283 -1988 4295 1988
rect 4237 -2000 4295 -1988
rect 4395 1988 4453 2000
rect 4395 -1988 4407 1988
rect 4441 -1988 4453 1988
rect 4395 -2000 4453 -1988
rect 4553 1988 4611 2000
rect 4553 -1988 4565 1988
rect 4599 -1988 4611 1988
rect 4553 -2000 4611 -1988
rect 4711 1988 4769 2000
rect 4711 -1988 4723 1988
rect 4757 -1988 4769 1988
rect 4711 -2000 4769 -1988
rect 4869 1988 4927 2000
rect 4869 -1988 4881 1988
rect 4915 -1988 4927 1988
rect 4869 -2000 4927 -1988
rect 5027 1988 5085 2000
rect 5027 -1988 5039 1988
rect 5073 -1988 5085 1988
rect 5027 -2000 5085 -1988
rect 5185 1988 5243 2000
rect 5185 -1988 5197 1988
rect 5231 -1988 5243 1988
rect 5185 -2000 5243 -1988
rect 5343 1988 5401 2000
rect 5343 -1988 5355 1988
rect 5389 -1988 5401 1988
rect 5343 -2000 5401 -1988
rect 5501 1988 5559 2000
rect 5501 -1988 5513 1988
rect 5547 -1988 5559 1988
rect 5501 -2000 5559 -1988
rect 5659 1988 5717 2000
rect 5659 -1988 5671 1988
rect 5705 -1988 5717 1988
rect 5659 -2000 5717 -1988
rect 5817 1988 5875 2000
rect 5817 -1988 5829 1988
rect 5863 -1988 5875 1988
rect 5817 -2000 5875 -1988
rect 5975 1988 6033 2000
rect 5975 -1988 5987 1988
rect 6021 -1988 6033 1988
rect 5975 -2000 6033 -1988
rect 6133 1988 6191 2000
rect 6133 -1988 6145 1988
rect 6179 -1988 6191 1988
rect 6133 -2000 6191 -1988
rect 6291 1988 6349 2000
rect 6291 -1988 6303 1988
rect 6337 -1988 6349 1988
rect 6291 -2000 6349 -1988
rect 6449 1988 6507 2000
rect 6449 -1988 6461 1988
rect 6495 -1988 6507 1988
rect 6449 -2000 6507 -1988
rect 6607 1988 6665 2000
rect 6607 -1988 6619 1988
rect 6653 -1988 6665 1988
rect 6607 -2000 6665 -1988
rect 6765 1988 6823 2000
rect 6765 -1988 6777 1988
rect 6811 -1988 6823 1988
rect 6765 -2000 6823 -1988
rect 6923 1988 6981 2000
rect 6923 -1988 6935 1988
rect 6969 -1988 6981 1988
rect 6923 -2000 6981 -1988
rect 7081 1988 7139 2000
rect 7081 -1988 7093 1988
rect 7127 -1988 7139 1988
rect 7081 -2000 7139 -1988
rect 7239 1988 7297 2000
rect 7239 -1988 7251 1988
rect 7285 -1988 7297 1988
rect 7239 -2000 7297 -1988
rect 7397 1988 7455 2000
rect 7397 -1988 7409 1988
rect 7443 -1988 7455 1988
rect 7397 -2000 7455 -1988
rect 7555 1988 7613 2000
rect 7555 -1988 7567 1988
rect 7601 -1988 7613 1988
rect 7555 -2000 7613 -1988
rect 7713 1988 7771 2000
rect 7713 -1988 7725 1988
rect 7759 -1988 7771 1988
rect 7713 -2000 7771 -1988
rect 7871 1988 7929 2000
rect 7871 -1988 7883 1988
rect 7917 -1988 7929 1988
rect 7871 -2000 7929 -1988
rect 8029 1988 8087 2000
rect 8029 -1988 8041 1988
rect 8075 -1988 8087 1988
rect 8029 -2000 8087 -1988
rect 8187 1988 8245 2000
rect 8187 -1988 8199 1988
rect 8233 -1988 8245 1988
rect 8187 -2000 8245 -1988
rect 8345 1988 8403 2000
rect 8345 -1988 8357 1988
rect 8391 -1988 8403 1988
rect 8345 -2000 8403 -1988
rect 8503 1988 8561 2000
rect 8503 -1988 8515 1988
rect 8549 -1988 8561 1988
rect 8503 -2000 8561 -1988
rect 8661 1988 8719 2000
rect 8661 -1988 8673 1988
rect 8707 -1988 8719 1988
rect 8661 -2000 8719 -1988
rect 8819 1988 8877 2000
rect 8819 -1988 8831 1988
rect 8865 -1988 8877 1988
rect 8819 -2000 8877 -1988
rect 8977 1988 9035 2000
rect 8977 -1988 8989 1988
rect 9023 -1988 9035 1988
rect 8977 -2000 9035 -1988
rect 9135 1988 9193 2000
rect 9135 -1988 9147 1988
rect 9181 -1988 9193 1988
rect 9135 -2000 9193 -1988
rect 9293 1988 9351 2000
rect 9293 -1988 9305 1988
rect 9339 -1988 9351 1988
rect 9293 -2000 9351 -1988
rect 9451 1988 9509 2000
rect 9451 -1988 9463 1988
rect 9497 -1988 9509 1988
rect 9451 -2000 9509 -1988
rect 9609 1988 9667 2000
rect 9609 -1988 9621 1988
rect 9655 -1988 9667 1988
rect 9609 -2000 9667 -1988
rect 9767 1988 9825 2000
rect 9767 -1988 9779 1988
rect 9813 -1988 9825 1988
rect 9767 -2000 9825 -1988
rect 9925 1988 9983 2000
rect 9925 -1988 9937 1988
rect 9971 -1988 9983 1988
rect 9925 -2000 9983 -1988
rect 10083 1988 10141 2000
rect 10083 -1988 10095 1988
rect 10129 -1988 10141 1988
rect 10083 -2000 10141 -1988
<< mvndiffc >>
rect -10129 -1988 -10095 1988
rect -9971 -1988 -9937 1988
rect -9813 -1988 -9779 1988
rect -9655 -1988 -9621 1988
rect -9497 -1988 -9463 1988
rect -9339 -1988 -9305 1988
rect -9181 -1988 -9147 1988
rect -9023 -1988 -8989 1988
rect -8865 -1988 -8831 1988
rect -8707 -1988 -8673 1988
rect -8549 -1988 -8515 1988
rect -8391 -1988 -8357 1988
rect -8233 -1988 -8199 1988
rect -8075 -1988 -8041 1988
rect -7917 -1988 -7883 1988
rect -7759 -1988 -7725 1988
rect -7601 -1988 -7567 1988
rect -7443 -1988 -7409 1988
rect -7285 -1988 -7251 1988
rect -7127 -1988 -7093 1988
rect -6969 -1988 -6935 1988
rect -6811 -1988 -6777 1988
rect -6653 -1988 -6619 1988
rect -6495 -1988 -6461 1988
rect -6337 -1988 -6303 1988
rect -6179 -1988 -6145 1988
rect -6021 -1988 -5987 1988
rect -5863 -1988 -5829 1988
rect -5705 -1988 -5671 1988
rect -5547 -1988 -5513 1988
rect -5389 -1988 -5355 1988
rect -5231 -1988 -5197 1988
rect -5073 -1988 -5039 1988
rect -4915 -1988 -4881 1988
rect -4757 -1988 -4723 1988
rect -4599 -1988 -4565 1988
rect -4441 -1988 -4407 1988
rect -4283 -1988 -4249 1988
rect -4125 -1988 -4091 1988
rect -3967 -1988 -3933 1988
rect -3809 -1988 -3775 1988
rect -3651 -1988 -3617 1988
rect -3493 -1988 -3459 1988
rect -3335 -1988 -3301 1988
rect -3177 -1988 -3143 1988
rect -3019 -1988 -2985 1988
rect -2861 -1988 -2827 1988
rect -2703 -1988 -2669 1988
rect -2545 -1988 -2511 1988
rect -2387 -1988 -2353 1988
rect -2229 -1988 -2195 1988
rect -2071 -1988 -2037 1988
rect -1913 -1988 -1879 1988
rect -1755 -1988 -1721 1988
rect -1597 -1988 -1563 1988
rect -1439 -1988 -1405 1988
rect -1281 -1988 -1247 1988
rect -1123 -1988 -1089 1988
rect -965 -1988 -931 1988
rect -807 -1988 -773 1988
rect -649 -1988 -615 1988
rect -491 -1988 -457 1988
rect -333 -1988 -299 1988
rect -175 -1988 -141 1988
rect -17 -1988 17 1988
rect 141 -1988 175 1988
rect 299 -1988 333 1988
rect 457 -1988 491 1988
rect 615 -1988 649 1988
rect 773 -1988 807 1988
rect 931 -1988 965 1988
rect 1089 -1988 1123 1988
rect 1247 -1988 1281 1988
rect 1405 -1988 1439 1988
rect 1563 -1988 1597 1988
rect 1721 -1988 1755 1988
rect 1879 -1988 1913 1988
rect 2037 -1988 2071 1988
rect 2195 -1988 2229 1988
rect 2353 -1988 2387 1988
rect 2511 -1988 2545 1988
rect 2669 -1988 2703 1988
rect 2827 -1988 2861 1988
rect 2985 -1988 3019 1988
rect 3143 -1988 3177 1988
rect 3301 -1988 3335 1988
rect 3459 -1988 3493 1988
rect 3617 -1988 3651 1988
rect 3775 -1988 3809 1988
rect 3933 -1988 3967 1988
rect 4091 -1988 4125 1988
rect 4249 -1988 4283 1988
rect 4407 -1988 4441 1988
rect 4565 -1988 4599 1988
rect 4723 -1988 4757 1988
rect 4881 -1988 4915 1988
rect 5039 -1988 5073 1988
rect 5197 -1988 5231 1988
rect 5355 -1988 5389 1988
rect 5513 -1988 5547 1988
rect 5671 -1988 5705 1988
rect 5829 -1988 5863 1988
rect 5987 -1988 6021 1988
rect 6145 -1988 6179 1988
rect 6303 -1988 6337 1988
rect 6461 -1988 6495 1988
rect 6619 -1988 6653 1988
rect 6777 -1988 6811 1988
rect 6935 -1988 6969 1988
rect 7093 -1988 7127 1988
rect 7251 -1988 7285 1988
rect 7409 -1988 7443 1988
rect 7567 -1988 7601 1988
rect 7725 -1988 7759 1988
rect 7883 -1988 7917 1988
rect 8041 -1988 8075 1988
rect 8199 -1988 8233 1988
rect 8357 -1988 8391 1988
rect 8515 -1988 8549 1988
rect 8673 -1988 8707 1988
rect 8831 -1988 8865 1988
rect 8989 -1988 9023 1988
rect 9147 -1988 9181 1988
rect 9305 -1988 9339 1988
rect 9463 -1988 9497 1988
rect 9621 -1988 9655 1988
rect 9779 -1988 9813 1988
rect 9937 -1988 9971 1988
rect 10095 -1988 10129 1988
<< mvpsubdiff >>
rect -10275 2210 10275 2222
rect -10275 2176 -10167 2210
rect 10167 2176 10275 2210
rect -10275 2164 10275 2176
rect -10275 2114 -10217 2164
rect -10275 -2114 -10263 2114
rect -10229 -2114 -10217 2114
rect 10217 2114 10275 2164
rect -10275 -2164 -10217 -2114
rect 10217 -2114 10229 2114
rect 10263 -2114 10275 2114
rect 10217 -2164 10275 -2114
rect -10275 -2176 10275 -2164
rect -10275 -2210 -10167 -2176
rect 10167 -2210 10275 -2176
rect -10275 -2222 10275 -2210
<< mvpsubdiffcont >>
rect -10167 2176 10167 2210
rect -10263 -2114 -10229 2114
rect 10229 -2114 10263 2114
rect -10167 -2210 10167 -2176
<< poly >>
rect -10083 2072 -9983 2088
rect -10083 2038 -10067 2072
rect -9999 2038 -9983 2072
rect -10083 2000 -9983 2038
rect -9925 2072 -9825 2088
rect -9925 2038 -9909 2072
rect -9841 2038 -9825 2072
rect -9925 2000 -9825 2038
rect -9767 2072 -9667 2088
rect -9767 2038 -9751 2072
rect -9683 2038 -9667 2072
rect -9767 2000 -9667 2038
rect -9609 2072 -9509 2088
rect -9609 2038 -9593 2072
rect -9525 2038 -9509 2072
rect -9609 2000 -9509 2038
rect -9451 2072 -9351 2088
rect -9451 2038 -9435 2072
rect -9367 2038 -9351 2072
rect -9451 2000 -9351 2038
rect -9293 2072 -9193 2088
rect -9293 2038 -9277 2072
rect -9209 2038 -9193 2072
rect -9293 2000 -9193 2038
rect -9135 2072 -9035 2088
rect -9135 2038 -9119 2072
rect -9051 2038 -9035 2072
rect -9135 2000 -9035 2038
rect -8977 2072 -8877 2088
rect -8977 2038 -8961 2072
rect -8893 2038 -8877 2072
rect -8977 2000 -8877 2038
rect -8819 2072 -8719 2088
rect -8819 2038 -8803 2072
rect -8735 2038 -8719 2072
rect -8819 2000 -8719 2038
rect -8661 2072 -8561 2088
rect -8661 2038 -8645 2072
rect -8577 2038 -8561 2072
rect -8661 2000 -8561 2038
rect -8503 2072 -8403 2088
rect -8503 2038 -8487 2072
rect -8419 2038 -8403 2072
rect -8503 2000 -8403 2038
rect -8345 2072 -8245 2088
rect -8345 2038 -8329 2072
rect -8261 2038 -8245 2072
rect -8345 2000 -8245 2038
rect -8187 2072 -8087 2088
rect -8187 2038 -8171 2072
rect -8103 2038 -8087 2072
rect -8187 2000 -8087 2038
rect -8029 2072 -7929 2088
rect -8029 2038 -8013 2072
rect -7945 2038 -7929 2072
rect -8029 2000 -7929 2038
rect -7871 2072 -7771 2088
rect -7871 2038 -7855 2072
rect -7787 2038 -7771 2072
rect -7871 2000 -7771 2038
rect -7713 2072 -7613 2088
rect -7713 2038 -7697 2072
rect -7629 2038 -7613 2072
rect -7713 2000 -7613 2038
rect -7555 2072 -7455 2088
rect -7555 2038 -7539 2072
rect -7471 2038 -7455 2072
rect -7555 2000 -7455 2038
rect -7397 2072 -7297 2088
rect -7397 2038 -7381 2072
rect -7313 2038 -7297 2072
rect -7397 2000 -7297 2038
rect -7239 2072 -7139 2088
rect -7239 2038 -7223 2072
rect -7155 2038 -7139 2072
rect -7239 2000 -7139 2038
rect -7081 2072 -6981 2088
rect -7081 2038 -7065 2072
rect -6997 2038 -6981 2072
rect -7081 2000 -6981 2038
rect -6923 2072 -6823 2088
rect -6923 2038 -6907 2072
rect -6839 2038 -6823 2072
rect -6923 2000 -6823 2038
rect -6765 2072 -6665 2088
rect -6765 2038 -6749 2072
rect -6681 2038 -6665 2072
rect -6765 2000 -6665 2038
rect -6607 2072 -6507 2088
rect -6607 2038 -6591 2072
rect -6523 2038 -6507 2072
rect -6607 2000 -6507 2038
rect -6449 2072 -6349 2088
rect -6449 2038 -6433 2072
rect -6365 2038 -6349 2072
rect -6449 2000 -6349 2038
rect -6291 2072 -6191 2088
rect -6291 2038 -6275 2072
rect -6207 2038 -6191 2072
rect -6291 2000 -6191 2038
rect -6133 2072 -6033 2088
rect -6133 2038 -6117 2072
rect -6049 2038 -6033 2072
rect -6133 2000 -6033 2038
rect -5975 2072 -5875 2088
rect -5975 2038 -5959 2072
rect -5891 2038 -5875 2072
rect -5975 2000 -5875 2038
rect -5817 2072 -5717 2088
rect -5817 2038 -5801 2072
rect -5733 2038 -5717 2072
rect -5817 2000 -5717 2038
rect -5659 2072 -5559 2088
rect -5659 2038 -5643 2072
rect -5575 2038 -5559 2072
rect -5659 2000 -5559 2038
rect -5501 2072 -5401 2088
rect -5501 2038 -5485 2072
rect -5417 2038 -5401 2072
rect -5501 2000 -5401 2038
rect -5343 2072 -5243 2088
rect -5343 2038 -5327 2072
rect -5259 2038 -5243 2072
rect -5343 2000 -5243 2038
rect -5185 2072 -5085 2088
rect -5185 2038 -5169 2072
rect -5101 2038 -5085 2072
rect -5185 2000 -5085 2038
rect -5027 2072 -4927 2088
rect -5027 2038 -5011 2072
rect -4943 2038 -4927 2072
rect -5027 2000 -4927 2038
rect -4869 2072 -4769 2088
rect -4869 2038 -4853 2072
rect -4785 2038 -4769 2072
rect -4869 2000 -4769 2038
rect -4711 2072 -4611 2088
rect -4711 2038 -4695 2072
rect -4627 2038 -4611 2072
rect -4711 2000 -4611 2038
rect -4553 2072 -4453 2088
rect -4553 2038 -4537 2072
rect -4469 2038 -4453 2072
rect -4553 2000 -4453 2038
rect -4395 2072 -4295 2088
rect -4395 2038 -4379 2072
rect -4311 2038 -4295 2072
rect -4395 2000 -4295 2038
rect -4237 2072 -4137 2088
rect -4237 2038 -4221 2072
rect -4153 2038 -4137 2072
rect -4237 2000 -4137 2038
rect -4079 2072 -3979 2088
rect -4079 2038 -4063 2072
rect -3995 2038 -3979 2072
rect -4079 2000 -3979 2038
rect -3921 2072 -3821 2088
rect -3921 2038 -3905 2072
rect -3837 2038 -3821 2072
rect -3921 2000 -3821 2038
rect -3763 2072 -3663 2088
rect -3763 2038 -3747 2072
rect -3679 2038 -3663 2072
rect -3763 2000 -3663 2038
rect -3605 2072 -3505 2088
rect -3605 2038 -3589 2072
rect -3521 2038 -3505 2072
rect -3605 2000 -3505 2038
rect -3447 2072 -3347 2088
rect -3447 2038 -3431 2072
rect -3363 2038 -3347 2072
rect -3447 2000 -3347 2038
rect -3289 2072 -3189 2088
rect -3289 2038 -3273 2072
rect -3205 2038 -3189 2072
rect -3289 2000 -3189 2038
rect -3131 2072 -3031 2088
rect -3131 2038 -3115 2072
rect -3047 2038 -3031 2072
rect -3131 2000 -3031 2038
rect -2973 2072 -2873 2088
rect -2973 2038 -2957 2072
rect -2889 2038 -2873 2072
rect -2973 2000 -2873 2038
rect -2815 2072 -2715 2088
rect -2815 2038 -2799 2072
rect -2731 2038 -2715 2072
rect -2815 2000 -2715 2038
rect -2657 2072 -2557 2088
rect -2657 2038 -2641 2072
rect -2573 2038 -2557 2072
rect -2657 2000 -2557 2038
rect -2499 2072 -2399 2088
rect -2499 2038 -2483 2072
rect -2415 2038 -2399 2072
rect -2499 2000 -2399 2038
rect -2341 2072 -2241 2088
rect -2341 2038 -2325 2072
rect -2257 2038 -2241 2072
rect -2341 2000 -2241 2038
rect -2183 2072 -2083 2088
rect -2183 2038 -2167 2072
rect -2099 2038 -2083 2072
rect -2183 2000 -2083 2038
rect -2025 2072 -1925 2088
rect -2025 2038 -2009 2072
rect -1941 2038 -1925 2072
rect -2025 2000 -1925 2038
rect -1867 2072 -1767 2088
rect -1867 2038 -1851 2072
rect -1783 2038 -1767 2072
rect -1867 2000 -1767 2038
rect -1709 2072 -1609 2088
rect -1709 2038 -1693 2072
rect -1625 2038 -1609 2072
rect -1709 2000 -1609 2038
rect -1551 2072 -1451 2088
rect -1551 2038 -1535 2072
rect -1467 2038 -1451 2072
rect -1551 2000 -1451 2038
rect -1393 2072 -1293 2088
rect -1393 2038 -1377 2072
rect -1309 2038 -1293 2072
rect -1393 2000 -1293 2038
rect -1235 2072 -1135 2088
rect -1235 2038 -1219 2072
rect -1151 2038 -1135 2072
rect -1235 2000 -1135 2038
rect -1077 2072 -977 2088
rect -1077 2038 -1061 2072
rect -993 2038 -977 2072
rect -1077 2000 -977 2038
rect -919 2072 -819 2088
rect -919 2038 -903 2072
rect -835 2038 -819 2072
rect -919 2000 -819 2038
rect -761 2072 -661 2088
rect -761 2038 -745 2072
rect -677 2038 -661 2072
rect -761 2000 -661 2038
rect -603 2072 -503 2088
rect -603 2038 -587 2072
rect -519 2038 -503 2072
rect -603 2000 -503 2038
rect -445 2072 -345 2088
rect -445 2038 -429 2072
rect -361 2038 -345 2072
rect -445 2000 -345 2038
rect -287 2072 -187 2088
rect -287 2038 -271 2072
rect -203 2038 -187 2072
rect -287 2000 -187 2038
rect -129 2072 -29 2088
rect -129 2038 -113 2072
rect -45 2038 -29 2072
rect -129 2000 -29 2038
rect 29 2072 129 2088
rect 29 2038 45 2072
rect 113 2038 129 2072
rect 29 2000 129 2038
rect 187 2072 287 2088
rect 187 2038 203 2072
rect 271 2038 287 2072
rect 187 2000 287 2038
rect 345 2072 445 2088
rect 345 2038 361 2072
rect 429 2038 445 2072
rect 345 2000 445 2038
rect 503 2072 603 2088
rect 503 2038 519 2072
rect 587 2038 603 2072
rect 503 2000 603 2038
rect 661 2072 761 2088
rect 661 2038 677 2072
rect 745 2038 761 2072
rect 661 2000 761 2038
rect 819 2072 919 2088
rect 819 2038 835 2072
rect 903 2038 919 2072
rect 819 2000 919 2038
rect 977 2072 1077 2088
rect 977 2038 993 2072
rect 1061 2038 1077 2072
rect 977 2000 1077 2038
rect 1135 2072 1235 2088
rect 1135 2038 1151 2072
rect 1219 2038 1235 2072
rect 1135 2000 1235 2038
rect 1293 2072 1393 2088
rect 1293 2038 1309 2072
rect 1377 2038 1393 2072
rect 1293 2000 1393 2038
rect 1451 2072 1551 2088
rect 1451 2038 1467 2072
rect 1535 2038 1551 2072
rect 1451 2000 1551 2038
rect 1609 2072 1709 2088
rect 1609 2038 1625 2072
rect 1693 2038 1709 2072
rect 1609 2000 1709 2038
rect 1767 2072 1867 2088
rect 1767 2038 1783 2072
rect 1851 2038 1867 2072
rect 1767 2000 1867 2038
rect 1925 2072 2025 2088
rect 1925 2038 1941 2072
rect 2009 2038 2025 2072
rect 1925 2000 2025 2038
rect 2083 2072 2183 2088
rect 2083 2038 2099 2072
rect 2167 2038 2183 2072
rect 2083 2000 2183 2038
rect 2241 2072 2341 2088
rect 2241 2038 2257 2072
rect 2325 2038 2341 2072
rect 2241 2000 2341 2038
rect 2399 2072 2499 2088
rect 2399 2038 2415 2072
rect 2483 2038 2499 2072
rect 2399 2000 2499 2038
rect 2557 2072 2657 2088
rect 2557 2038 2573 2072
rect 2641 2038 2657 2072
rect 2557 2000 2657 2038
rect 2715 2072 2815 2088
rect 2715 2038 2731 2072
rect 2799 2038 2815 2072
rect 2715 2000 2815 2038
rect 2873 2072 2973 2088
rect 2873 2038 2889 2072
rect 2957 2038 2973 2072
rect 2873 2000 2973 2038
rect 3031 2072 3131 2088
rect 3031 2038 3047 2072
rect 3115 2038 3131 2072
rect 3031 2000 3131 2038
rect 3189 2072 3289 2088
rect 3189 2038 3205 2072
rect 3273 2038 3289 2072
rect 3189 2000 3289 2038
rect 3347 2072 3447 2088
rect 3347 2038 3363 2072
rect 3431 2038 3447 2072
rect 3347 2000 3447 2038
rect 3505 2072 3605 2088
rect 3505 2038 3521 2072
rect 3589 2038 3605 2072
rect 3505 2000 3605 2038
rect 3663 2072 3763 2088
rect 3663 2038 3679 2072
rect 3747 2038 3763 2072
rect 3663 2000 3763 2038
rect 3821 2072 3921 2088
rect 3821 2038 3837 2072
rect 3905 2038 3921 2072
rect 3821 2000 3921 2038
rect 3979 2072 4079 2088
rect 3979 2038 3995 2072
rect 4063 2038 4079 2072
rect 3979 2000 4079 2038
rect 4137 2072 4237 2088
rect 4137 2038 4153 2072
rect 4221 2038 4237 2072
rect 4137 2000 4237 2038
rect 4295 2072 4395 2088
rect 4295 2038 4311 2072
rect 4379 2038 4395 2072
rect 4295 2000 4395 2038
rect 4453 2072 4553 2088
rect 4453 2038 4469 2072
rect 4537 2038 4553 2072
rect 4453 2000 4553 2038
rect 4611 2072 4711 2088
rect 4611 2038 4627 2072
rect 4695 2038 4711 2072
rect 4611 2000 4711 2038
rect 4769 2072 4869 2088
rect 4769 2038 4785 2072
rect 4853 2038 4869 2072
rect 4769 2000 4869 2038
rect 4927 2072 5027 2088
rect 4927 2038 4943 2072
rect 5011 2038 5027 2072
rect 4927 2000 5027 2038
rect 5085 2072 5185 2088
rect 5085 2038 5101 2072
rect 5169 2038 5185 2072
rect 5085 2000 5185 2038
rect 5243 2072 5343 2088
rect 5243 2038 5259 2072
rect 5327 2038 5343 2072
rect 5243 2000 5343 2038
rect 5401 2072 5501 2088
rect 5401 2038 5417 2072
rect 5485 2038 5501 2072
rect 5401 2000 5501 2038
rect 5559 2072 5659 2088
rect 5559 2038 5575 2072
rect 5643 2038 5659 2072
rect 5559 2000 5659 2038
rect 5717 2072 5817 2088
rect 5717 2038 5733 2072
rect 5801 2038 5817 2072
rect 5717 2000 5817 2038
rect 5875 2072 5975 2088
rect 5875 2038 5891 2072
rect 5959 2038 5975 2072
rect 5875 2000 5975 2038
rect 6033 2072 6133 2088
rect 6033 2038 6049 2072
rect 6117 2038 6133 2072
rect 6033 2000 6133 2038
rect 6191 2072 6291 2088
rect 6191 2038 6207 2072
rect 6275 2038 6291 2072
rect 6191 2000 6291 2038
rect 6349 2072 6449 2088
rect 6349 2038 6365 2072
rect 6433 2038 6449 2072
rect 6349 2000 6449 2038
rect 6507 2072 6607 2088
rect 6507 2038 6523 2072
rect 6591 2038 6607 2072
rect 6507 2000 6607 2038
rect 6665 2072 6765 2088
rect 6665 2038 6681 2072
rect 6749 2038 6765 2072
rect 6665 2000 6765 2038
rect 6823 2072 6923 2088
rect 6823 2038 6839 2072
rect 6907 2038 6923 2072
rect 6823 2000 6923 2038
rect 6981 2072 7081 2088
rect 6981 2038 6997 2072
rect 7065 2038 7081 2072
rect 6981 2000 7081 2038
rect 7139 2072 7239 2088
rect 7139 2038 7155 2072
rect 7223 2038 7239 2072
rect 7139 2000 7239 2038
rect 7297 2072 7397 2088
rect 7297 2038 7313 2072
rect 7381 2038 7397 2072
rect 7297 2000 7397 2038
rect 7455 2072 7555 2088
rect 7455 2038 7471 2072
rect 7539 2038 7555 2072
rect 7455 2000 7555 2038
rect 7613 2072 7713 2088
rect 7613 2038 7629 2072
rect 7697 2038 7713 2072
rect 7613 2000 7713 2038
rect 7771 2072 7871 2088
rect 7771 2038 7787 2072
rect 7855 2038 7871 2072
rect 7771 2000 7871 2038
rect 7929 2072 8029 2088
rect 7929 2038 7945 2072
rect 8013 2038 8029 2072
rect 7929 2000 8029 2038
rect 8087 2072 8187 2088
rect 8087 2038 8103 2072
rect 8171 2038 8187 2072
rect 8087 2000 8187 2038
rect 8245 2072 8345 2088
rect 8245 2038 8261 2072
rect 8329 2038 8345 2072
rect 8245 2000 8345 2038
rect 8403 2072 8503 2088
rect 8403 2038 8419 2072
rect 8487 2038 8503 2072
rect 8403 2000 8503 2038
rect 8561 2072 8661 2088
rect 8561 2038 8577 2072
rect 8645 2038 8661 2072
rect 8561 2000 8661 2038
rect 8719 2072 8819 2088
rect 8719 2038 8735 2072
rect 8803 2038 8819 2072
rect 8719 2000 8819 2038
rect 8877 2072 8977 2088
rect 8877 2038 8893 2072
rect 8961 2038 8977 2072
rect 8877 2000 8977 2038
rect 9035 2072 9135 2088
rect 9035 2038 9051 2072
rect 9119 2038 9135 2072
rect 9035 2000 9135 2038
rect 9193 2072 9293 2088
rect 9193 2038 9209 2072
rect 9277 2038 9293 2072
rect 9193 2000 9293 2038
rect 9351 2072 9451 2088
rect 9351 2038 9367 2072
rect 9435 2038 9451 2072
rect 9351 2000 9451 2038
rect 9509 2072 9609 2088
rect 9509 2038 9525 2072
rect 9593 2038 9609 2072
rect 9509 2000 9609 2038
rect 9667 2072 9767 2088
rect 9667 2038 9683 2072
rect 9751 2038 9767 2072
rect 9667 2000 9767 2038
rect 9825 2072 9925 2088
rect 9825 2038 9841 2072
rect 9909 2038 9925 2072
rect 9825 2000 9925 2038
rect 9983 2072 10083 2088
rect 9983 2038 9999 2072
rect 10067 2038 10083 2072
rect 9983 2000 10083 2038
rect -10083 -2038 -9983 -2000
rect -10083 -2072 -10067 -2038
rect -9999 -2072 -9983 -2038
rect -10083 -2088 -9983 -2072
rect -9925 -2038 -9825 -2000
rect -9925 -2072 -9909 -2038
rect -9841 -2072 -9825 -2038
rect -9925 -2088 -9825 -2072
rect -9767 -2038 -9667 -2000
rect -9767 -2072 -9751 -2038
rect -9683 -2072 -9667 -2038
rect -9767 -2088 -9667 -2072
rect -9609 -2038 -9509 -2000
rect -9609 -2072 -9593 -2038
rect -9525 -2072 -9509 -2038
rect -9609 -2088 -9509 -2072
rect -9451 -2038 -9351 -2000
rect -9451 -2072 -9435 -2038
rect -9367 -2072 -9351 -2038
rect -9451 -2088 -9351 -2072
rect -9293 -2038 -9193 -2000
rect -9293 -2072 -9277 -2038
rect -9209 -2072 -9193 -2038
rect -9293 -2088 -9193 -2072
rect -9135 -2038 -9035 -2000
rect -9135 -2072 -9119 -2038
rect -9051 -2072 -9035 -2038
rect -9135 -2088 -9035 -2072
rect -8977 -2038 -8877 -2000
rect -8977 -2072 -8961 -2038
rect -8893 -2072 -8877 -2038
rect -8977 -2088 -8877 -2072
rect -8819 -2038 -8719 -2000
rect -8819 -2072 -8803 -2038
rect -8735 -2072 -8719 -2038
rect -8819 -2088 -8719 -2072
rect -8661 -2038 -8561 -2000
rect -8661 -2072 -8645 -2038
rect -8577 -2072 -8561 -2038
rect -8661 -2088 -8561 -2072
rect -8503 -2038 -8403 -2000
rect -8503 -2072 -8487 -2038
rect -8419 -2072 -8403 -2038
rect -8503 -2088 -8403 -2072
rect -8345 -2038 -8245 -2000
rect -8345 -2072 -8329 -2038
rect -8261 -2072 -8245 -2038
rect -8345 -2088 -8245 -2072
rect -8187 -2038 -8087 -2000
rect -8187 -2072 -8171 -2038
rect -8103 -2072 -8087 -2038
rect -8187 -2088 -8087 -2072
rect -8029 -2038 -7929 -2000
rect -8029 -2072 -8013 -2038
rect -7945 -2072 -7929 -2038
rect -8029 -2088 -7929 -2072
rect -7871 -2038 -7771 -2000
rect -7871 -2072 -7855 -2038
rect -7787 -2072 -7771 -2038
rect -7871 -2088 -7771 -2072
rect -7713 -2038 -7613 -2000
rect -7713 -2072 -7697 -2038
rect -7629 -2072 -7613 -2038
rect -7713 -2088 -7613 -2072
rect -7555 -2038 -7455 -2000
rect -7555 -2072 -7539 -2038
rect -7471 -2072 -7455 -2038
rect -7555 -2088 -7455 -2072
rect -7397 -2038 -7297 -2000
rect -7397 -2072 -7381 -2038
rect -7313 -2072 -7297 -2038
rect -7397 -2088 -7297 -2072
rect -7239 -2038 -7139 -2000
rect -7239 -2072 -7223 -2038
rect -7155 -2072 -7139 -2038
rect -7239 -2088 -7139 -2072
rect -7081 -2038 -6981 -2000
rect -7081 -2072 -7065 -2038
rect -6997 -2072 -6981 -2038
rect -7081 -2088 -6981 -2072
rect -6923 -2038 -6823 -2000
rect -6923 -2072 -6907 -2038
rect -6839 -2072 -6823 -2038
rect -6923 -2088 -6823 -2072
rect -6765 -2038 -6665 -2000
rect -6765 -2072 -6749 -2038
rect -6681 -2072 -6665 -2038
rect -6765 -2088 -6665 -2072
rect -6607 -2038 -6507 -2000
rect -6607 -2072 -6591 -2038
rect -6523 -2072 -6507 -2038
rect -6607 -2088 -6507 -2072
rect -6449 -2038 -6349 -2000
rect -6449 -2072 -6433 -2038
rect -6365 -2072 -6349 -2038
rect -6449 -2088 -6349 -2072
rect -6291 -2038 -6191 -2000
rect -6291 -2072 -6275 -2038
rect -6207 -2072 -6191 -2038
rect -6291 -2088 -6191 -2072
rect -6133 -2038 -6033 -2000
rect -6133 -2072 -6117 -2038
rect -6049 -2072 -6033 -2038
rect -6133 -2088 -6033 -2072
rect -5975 -2038 -5875 -2000
rect -5975 -2072 -5959 -2038
rect -5891 -2072 -5875 -2038
rect -5975 -2088 -5875 -2072
rect -5817 -2038 -5717 -2000
rect -5817 -2072 -5801 -2038
rect -5733 -2072 -5717 -2038
rect -5817 -2088 -5717 -2072
rect -5659 -2038 -5559 -2000
rect -5659 -2072 -5643 -2038
rect -5575 -2072 -5559 -2038
rect -5659 -2088 -5559 -2072
rect -5501 -2038 -5401 -2000
rect -5501 -2072 -5485 -2038
rect -5417 -2072 -5401 -2038
rect -5501 -2088 -5401 -2072
rect -5343 -2038 -5243 -2000
rect -5343 -2072 -5327 -2038
rect -5259 -2072 -5243 -2038
rect -5343 -2088 -5243 -2072
rect -5185 -2038 -5085 -2000
rect -5185 -2072 -5169 -2038
rect -5101 -2072 -5085 -2038
rect -5185 -2088 -5085 -2072
rect -5027 -2038 -4927 -2000
rect -5027 -2072 -5011 -2038
rect -4943 -2072 -4927 -2038
rect -5027 -2088 -4927 -2072
rect -4869 -2038 -4769 -2000
rect -4869 -2072 -4853 -2038
rect -4785 -2072 -4769 -2038
rect -4869 -2088 -4769 -2072
rect -4711 -2038 -4611 -2000
rect -4711 -2072 -4695 -2038
rect -4627 -2072 -4611 -2038
rect -4711 -2088 -4611 -2072
rect -4553 -2038 -4453 -2000
rect -4553 -2072 -4537 -2038
rect -4469 -2072 -4453 -2038
rect -4553 -2088 -4453 -2072
rect -4395 -2038 -4295 -2000
rect -4395 -2072 -4379 -2038
rect -4311 -2072 -4295 -2038
rect -4395 -2088 -4295 -2072
rect -4237 -2038 -4137 -2000
rect -4237 -2072 -4221 -2038
rect -4153 -2072 -4137 -2038
rect -4237 -2088 -4137 -2072
rect -4079 -2038 -3979 -2000
rect -4079 -2072 -4063 -2038
rect -3995 -2072 -3979 -2038
rect -4079 -2088 -3979 -2072
rect -3921 -2038 -3821 -2000
rect -3921 -2072 -3905 -2038
rect -3837 -2072 -3821 -2038
rect -3921 -2088 -3821 -2072
rect -3763 -2038 -3663 -2000
rect -3763 -2072 -3747 -2038
rect -3679 -2072 -3663 -2038
rect -3763 -2088 -3663 -2072
rect -3605 -2038 -3505 -2000
rect -3605 -2072 -3589 -2038
rect -3521 -2072 -3505 -2038
rect -3605 -2088 -3505 -2072
rect -3447 -2038 -3347 -2000
rect -3447 -2072 -3431 -2038
rect -3363 -2072 -3347 -2038
rect -3447 -2088 -3347 -2072
rect -3289 -2038 -3189 -2000
rect -3289 -2072 -3273 -2038
rect -3205 -2072 -3189 -2038
rect -3289 -2088 -3189 -2072
rect -3131 -2038 -3031 -2000
rect -3131 -2072 -3115 -2038
rect -3047 -2072 -3031 -2038
rect -3131 -2088 -3031 -2072
rect -2973 -2038 -2873 -2000
rect -2973 -2072 -2957 -2038
rect -2889 -2072 -2873 -2038
rect -2973 -2088 -2873 -2072
rect -2815 -2038 -2715 -2000
rect -2815 -2072 -2799 -2038
rect -2731 -2072 -2715 -2038
rect -2815 -2088 -2715 -2072
rect -2657 -2038 -2557 -2000
rect -2657 -2072 -2641 -2038
rect -2573 -2072 -2557 -2038
rect -2657 -2088 -2557 -2072
rect -2499 -2038 -2399 -2000
rect -2499 -2072 -2483 -2038
rect -2415 -2072 -2399 -2038
rect -2499 -2088 -2399 -2072
rect -2341 -2038 -2241 -2000
rect -2341 -2072 -2325 -2038
rect -2257 -2072 -2241 -2038
rect -2341 -2088 -2241 -2072
rect -2183 -2038 -2083 -2000
rect -2183 -2072 -2167 -2038
rect -2099 -2072 -2083 -2038
rect -2183 -2088 -2083 -2072
rect -2025 -2038 -1925 -2000
rect -2025 -2072 -2009 -2038
rect -1941 -2072 -1925 -2038
rect -2025 -2088 -1925 -2072
rect -1867 -2038 -1767 -2000
rect -1867 -2072 -1851 -2038
rect -1783 -2072 -1767 -2038
rect -1867 -2088 -1767 -2072
rect -1709 -2038 -1609 -2000
rect -1709 -2072 -1693 -2038
rect -1625 -2072 -1609 -2038
rect -1709 -2088 -1609 -2072
rect -1551 -2038 -1451 -2000
rect -1551 -2072 -1535 -2038
rect -1467 -2072 -1451 -2038
rect -1551 -2088 -1451 -2072
rect -1393 -2038 -1293 -2000
rect -1393 -2072 -1377 -2038
rect -1309 -2072 -1293 -2038
rect -1393 -2088 -1293 -2072
rect -1235 -2038 -1135 -2000
rect -1235 -2072 -1219 -2038
rect -1151 -2072 -1135 -2038
rect -1235 -2088 -1135 -2072
rect -1077 -2038 -977 -2000
rect -1077 -2072 -1061 -2038
rect -993 -2072 -977 -2038
rect -1077 -2088 -977 -2072
rect -919 -2038 -819 -2000
rect -919 -2072 -903 -2038
rect -835 -2072 -819 -2038
rect -919 -2088 -819 -2072
rect -761 -2038 -661 -2000
rect -761 -2072 -745 -2038
rect -677 -2072 -661 -2038
rect -761 -2088 -661 -2072
rect -603 -2038 -503 -2000
rect -603 -2072 -587 -2038
rect -519 -2072 -503 -2038
rect -603 -2088 -503 -2072
rect -445 -2038 -345 -2000
rect -445 -2072 -429 -2038
rect -361 -2072 -345 -2038
rect -445 -2088 -345 -2072
rect -287 -2038 -187 -2000
rect -287 -2072 -271 -2038
rect -203 -2072 -187 -2038
rect -287 -2088 -187 -2072
rect -129 -2038 -29 -2000
rect -129 -2072 -113 -2038
rect -45 -2072 -29 -2038
rect -129 -2088 -29 -2072
rect 29 -2038 129 -2000
rect 29 -2072 45 -2038
rect 113 -2072 129 -2038
rect 29 -2088 129 -2072
rect 187 -2038 287 -2000
rect 187 -2072 203 -2038
rect 271 -2072 287 -2038
rect 187 -2088 287 -2072
rect 345 -2038 445 -2000
rect 345 -2072 361 -2038
rect 429 -2072 445 -2038
rect 345 -2088 445 -2072
rect 503 -2038 603 -2000
rect 503 -2072 519 -2038
rect 587 -2072 603 -2038
rect 503 -2088 603 -2072
rect 661 -2038 761 -2000
rect 661 -2072 677 -2038
rect 745 -2072 761 -2038
rect 661 -2088 761 -2072
rect 819 -2038 919 -2000
rect 819 -2072 835 -2038
rect 903 -2072 919 -2038
rect 819 -2088 919 -2072
rect 977 -2038 1077 -2000
rect 977 -2072 993 -2038
rect 1061 -2072 1077 -2038
rect 977 -2088 1077 -2072
rect 1135 -2038 1235 -2000
rect 1135 -2072 1151 -2038
rect 1219 -2072 1235 -2038
rect 1135 -2088 1235 -2072
rect 1293 -2038 1393 -2000
rect 1293 -2072 1309 -2038
rect 1377 -2072 1393 -2038
rect 1293 -2088 1393 -2072
rect 1451 -2038 1551 -2000
rect 1451 -2072 1467 -2038
rect 1535 -2072 1551 -2038
rect 1451 -2088 1551 -2072
rect 1609 -2038 1709 -2000
rect 1609 -2072 1625 -2038
rect 1693 -2072 1709 -2038
rect 1609 -2088 1709 -2072
rect 1767 -2038 1867 -2000
rect 1767 -2072 1783 -2038
rect 1851 -2072 1867 -2038
rect 1767 -2088 1867 -2072
rect 1925 -2038 2025 -2000
rect 1925 -2072 1941 -2038
rect 2009 -2072 2025 -2038
rect 1925 -2088 2025 -2072
rect 2083 -2038 2183 -2000
rect 2083 -2072 2099 -2038
rect 2167 -2072 2183 -2038
rect 2083 -2088 2183 -2072
rect 2241 -2038 2341 -2000
rect 2241 -2072 2257 -2038
rect 2325 -2072 2341 -2038
rect 2241 -2088 2341 -2072
rect 2399 -2038 2499 -2000
rect 2399 -2072 2415 -2038
rect 2483 -2072 2499 -2038
rect 2399 -2088 2499 -2072
rect 2557 -2038 2657 -2000
rect 2557 -2072 2573 -2038
rect 2641 -2072 2657 -2038
rect 2557 -2088 2657 -2072
rect 2715 -2038 2815 -2000
rect 2715 -2072 2731 -2038
rect 2799 -2072 2815 -2038
rect 2715 -2088 2815 -2072
rect 2873 -2038 2973 -2000
rect 2873 -2072 2889 -2038
rect 2957 -2072 2973 -2038
rect 2873 -2088 2973 -2072
rect 3031 -2038 3131 -2000
rect 3031 -2072 3047 -2038
rect 3115 -2072 3131 -2038
rect 3031 -2088 3131 -2072
rect 3189 -2038 3289 -2000
rect 3189 -2072 3205 -2038
rect 3273 -2072 3289 -2038
rect 3189 -2088 3289 -2072
rect 3347 -2038 3447 -2000
rect 3347 -2072 3363 -2038
rect 3431 -2072 3447 -2038
rect 3347 -2088 3447 -2072
rect 3505 -2038 3605 -2000
rect 3505 -2072 3521 -2038
rect 3589 -2072 3605 -2038
rect 3505 -2088 3605 -2072
rect 3663 -2038 3763 -2000
rect 3663 -2072 3679 -2038
rect 3747 -2072 3763 -2038
rect 3663 -2088 3763 -2072
rect 3821 -2038 3921 -2000
rect 3821 -2072 3837 -2038
rect 3905 -2072 3921 -2038
rect 3821 -2088 3921 -2072
rect 3979 -2038 4079 -2000
rect 3979 -2072 3995 -2038
rect 4063 -2072 4079 -2038
rect 3979 -2088 4079 -2072
rect 4137 -2038 4237 -2000
rect 4137 -2072 4153 -2038
rect 4221 -2072 4237 -2038
rect 4137 -2088 4237 -2072
rect 4295 -2038 4395 -2000
rect 4295 -2072 4311 -2038
rect 4379 -2072 4395 -2038
rect 4295 -2088 4395 -2072
rect 4453 -2038 4553 -2000
rect 4453 -2072 4469 -2038
rect 4537 -2072 4553 -2038
rect 4453 -2088 4553 -2072
rect 4611 -2038 4711 -2000
rect 4611 -2072 4627 -2038
rect 4695 -2072 4711 -2038
rect 4611 -2088 4711 -2072
rect 4769 -2038 4869 -2000
rect 4769 -2072 4785 -2038
rect 4853 -2072 4869 -2038
rect 4769 -2088 4869 -2072
rect 4927 -2038 5027 -2000
rect 4927 -2072 4943 -2038
rect 5011 -2072 5027 -2038
rect 4927 -2088 5027 -2072
rect 5085 -2038 5185 -2000
rect 5085 -2072 5101 -2038
rect 5169 -2072 5185 -2038
rect 5085 -2088 5185 -2072
rect 5243 -2038 5343 -2000
rect 5243 -2072 5259 -2038
rect 5327 -2072 5343 -2038
rect 5243 -2088 5343 -2072
rect 5401 -2038 5501 -2000
rect 5401 -2072 5417 -2038
rect 5485 -2072 5501 -2038
rect 5401 -2088 5501 -2072
rect 5559 -2038 5659 -2000
rect 5559 -2072 5575 -2038
rect 5643 -2072 5659 -2038
rect 5559 -2088 5659 -2072
rect 5717 -2038 5817 -2000
rect 5717 -2072 5733 -2038
rect 5801 -2072 5817 -2038
rect 5717 -2088 5817 -2072
rect 5875 -2038 5975 -2000
rect 5875 -2072 5891 -2038
rect 5959 -2072 5975 -2038
rect 5875 -2088 5975 -2072
rect 6033 -2038 6133 -2000
rect 6033 -2072 6049 -2038
rect 6117 -2072 6133 -2038
rect 6033 -2088 6133 -2072
rect 6191 -2038 6291 -2000
rect 6191 -2072 6207 -2038
rect 6275 -2072 6291 -2038
rect 6191 -2088 6291 -2072
rect 6349 -2038 6449 -2000
rect 6349 -2072 6365 -2038
rect 6433 -2072 6449 -2038
rect 6349 -2088 6449 -2072
rect 6507 -2038 6607 -2000
rect 6507 -2072 6523 -2038
rect 6591 -2072 6607 -2038
rect 6507 -2088 6607 -2072
rect 6665 -2038 6765 -2000
rect 6665 -2072 6681 -2038
rect 6749 -2072 6765 -2038
rect 6665 -2088 6765 -2072
rect 6823 -2038 6923 -2000
rect 6823 -2072 6839 -2038
rect 6907 -2072 6923 -2038
rect 6823 -2088 6923 -2072
rect 6981 -2038 7081 -2000
rect 6981 -2072 6997 -2038
rect 7065 -2072 7081 -2038
rect 6981 -2088 7081 -2072
rect 7139 -2038 7239 -2000
rect 7139 -2072 7155 -2038
rect 7223 -2072 7239 -2038
rect 7139 -2088 7239 -2072
rect 7297 -2038 7397 -2000
rect 7297 -2072 7313 -2038
rect 7381 -2072 7397 -2038
rect 7297 -2088 7397 -2072
rect 7455 -2038 7555 -2000
rect 7455 -2072 7471 -2038
rect 7539 -2072 7555 -2038
rect 7455 -2088 7555 -2072
rect 7613 -2038 7713 -2000
rect 7613 -2072 7629 -2038
rect 7697 -2072 7713 -2038
rect 7613 -2088 7713 -2072
rect 7771 -2038 7871 -2000
rect 7771 -2072 7787 -2038
rect 7855 -2072 7871 -2038
rect 7771 -2088 7871 -2072
rect 7929 -2038 8029 -2000
rect 7929 -2072 7945 -2038
rect 8013 -2072 8029 -2038
rect 7929 -2088 8029 -2072
rect 8087 -2038 8187 -2000
rect 8087 -2072 8103 -2038
rect 8171 -2072 8187 -2038
rect 8087 -2088 8187 -2072
rect 8245 -2038 8345 -2000
rect 8245 -2072 8261 -2038
rect 8329 -2072 8345 -2038
rect 8245 -2088 8345 -2072
rect 8403 -2038 8503 -2000
rect 8403 -2072 8419 -2038
rect 8487 -2072 8503 -2038
rect 8403 -2088 8503 -2072
rect 8561 -2038 8661 -2000
rect 8561 -2072 8577 -2038
rect 8645 -2072 8661 -2038
rect 8561 -2088 8661 -2072
rect 8719 -2038 8819 -2000
rect 8719 -2072 8735 -2038
rect 8803 -2072 8819 -2038
rect 8719 -2088 8819 -2072
rect 8877 -2038 8977 -2000
rect 8877 -2072 8893 -2038
rect 8961 -2072 8977 -2038
rect 8877 -2088 8977 -2072
rect 9035 -2038 9135 -2000
rect 9035 -2072 9051 -2038
rect 9119 -2072 9135 -2038
rect 9035 -2088 9135 -2072
rect 9193 -2038 9293 -2000
rect 9193 -2072 9209 -2038
rect 9277 -2072 9293 -2038
rect 9193 -2088 9293 -2072
rect 9351 -2038 9451 -2000
rect 9351 -2072 9367 -2038
rect 9435 -2072 9451 -2038
rect 9351 -2088 9451 -2072
rect 9509 -2038 9609 -2000
rect 9509 -2072 9525 -2038
rect 9593 -2072 9609 -2038
rect 9509 -2088 9609 -2072
rect 9667 -2038 9767 -2000
rect 9667 -2072 9683 -2038
rect 9751 -2072 9767 -2038
rect 9667 -2088 9767 -2072
rect 9825 -2038 9925 -2000
rect 9825 -2072 9841 -2038
rect 9909 -2072 9925 -2038
rect 9825 -2088 9925 -2072
rect 9983 -2038 10083 -2000
rect 9983 -2072 9999 -2038
rect 10067 -2072 10083 -2038
rect 9983 -2088 10083 -2072
<< polycont >>
rect -10067 2038 -9999 2072
rect -9909 2038 -9841 2072
rect -9751 2038 -9683 2072
rect -9593 2038 -9525 2072
rect -9435 2038 -9367 2072
rect -9277 2038 -9209 2072
rect -9119 2038 -9051 2072
rect -8961 2038 -8893 2072
rect -8803 2038 -8735 2072
rect -8645 2038 -8577 2072
rect -8487 2038 -8419 2072
rect -8329 2038 -8261 2072
rect -8171 2038 -8103 2072
rect -8013 2038 -7945 2072
rect -7855 2038 -7787 2072
rect -7697 2038 -7629 2072
rect -7539 2038 -7471 2072
rect -7381 2038 -7313 2072
rect -7223 2038 -7155 2072
rect -7065 2038 -6997 2072
rect -6907 2038 -6839 2072
rect -6749 2038 -6681 2072
rect -6591 2038 -6523 2072
rect -6433 2038 -6365 2072
rect -6275 2038 -6207 2072
rect -6117 2038 -6049 2072
rect -5959 2038 -5891 2072
rect -5801 2038 -5733 2072
rect -5643 2038 -5575 2072
rect -5485 2038 -5417 2072
rect -5327 2038 -5259 2072
rect -5169 2038 -5101 2072
rect -5011 2038 -4943 2072
rect -4853 2038 -4785 2072
rect -4695 2038 -4627 2072
rect -4537 2038 -4469 2072
rect -4379 2038 -4311 2072
rect -4221 2038 -4153 2072
rect -4063 2038 -3995 2072
rect -3905 2038 -3837 2072
rect -3747 2038 -3679 2072
rect -3589 2038 -3521 2072
rect -3431 2038 -3363 2072
rect -3273 2038 -3205 2072
rect -3115 2038 -3047 2072
rect -2957 2038 -2889 2072
rect -2799 2038 -2731 2072
rect -2641 2038 -2573 2072
rect -2483 2038 -2415 2072
rect -2325 2038 -2257 2072
rect -2167 2038 -2099 2072
rect -2009 2038 -1941 2072
rect -1851 2038 -1783 2072
rect -1693 2038 -1625 2072
rect -1535 2038 -1467 2072
rect -1377 2038 -1309 2072
rect -1219 2038 -1151 2072
rect -1061 2038 -993 2072
rect -903 2038 -835 2072
rect -745 2038 -677 2072
rect -587 2038 -519 2072
rect -429 2038 -361 2072
rect -271 2038 -203 2072
rect -113 2038 -45 2072
rect 45 2038 113 2072
rect 203 2038 271 2072
rect 361 2038 429 2072
rect 519 2038 587 2072
rect 677 2038 745 2072
rect 835 2038 903 2072
rect 993 2038 1061 2072
rect 1151 2038 1219 2072
rect 1309 2038 1377 2072
rect 1467 2038 1535 2072
rect 1625 2038 1693 2072
rect 1783 2038 1851 2072
rect 1941 2038 2009 2072
rect 2099 2038 2167 2072
rect 2257 2038 2325 2072
rect 2415 2038 2483 2072
rect 2573 2038 2641 2072
rect 2731 2038 2799 2072
rect 2889 2038 2957 2072
rect 3047 2038 3115 2072
rect 3205 2038 3273 2072
rect 3363 2038 3431 2072
rect 3521 2038 3589 2072
rect 3679 2038 3747 2072
rect 3837 2038 3905 2072
rect 3995 2038 4063 2072
rect 4153 2038 4221 2072
rect 4311 2038 4379 2072
rect 4469 2038 4537 2072
rect 4627 2038 4695 2072
rect 4785 2038 4853 2072
rect 4943 2038 5011 2072
rect 5101 2038 5169 2072
rect 5259 2038 5327 2072
rect 5417 2038 5485 2072
rect 5575 2038 5643 2072
rect 5733 2038 5801 2072
rect 5891 2038 5959 2072
rect 6049 2038 6117 2072
rect 6207 2038 6275 2072
rect 6365 2038 6433 2072
rect 6523 2038 6591 2072
rect 6681 2038 6749 2072
rect 6839 2038 6907 2072
rect 6997 2038 7065 2072
rect 7155 2038 7223 2072
rect 7313 2038 7381 2072
rect 7471 2038 7539 2072
rect 7629 2038 7697 2072
rect 7787 2038 7855 2072
rect 7945 2038 8013 2072
rect 8103 2038 8171 2072
rect 8261 2038 8329 2072
rect 8419 2038 8487 2072
rect 8577 2038 8645 2072
rect 8735 2038 8803 2072
rect 8893 2038 8961 2072
rect 9051 2038 9119 2072
rect 9209 2038 9277 2072
rect 9367 2038 9435 2072
rect 9525 2038 9593 2072
rect 9683 2038 9751 2072
rect 9841 2038 9909 2072
rect 9999 2038 10067 2072
rect -10067 -2072 -9999 -2038
rect -9909 -2072 -9841 -2038
rect -9751 -2072 -9683 -2038
rect -9593 -2072 -9525 -2038
rect -9435 -2072 -9367 -2038
rect -9277 -2072 -9209 -2038
rect -9119 -2072 -9051 -2038
rect -8961 -2072 -8893 -2038
rect -8803 -2072 -8735 -2038
rect -8645 -2072 -8577 -2038
rect -8487 -2072 -8419 -2038
rect -8329 -2072 -8261 -2038
rect -8171 -2072 -8103 -2038
rect -8013 -2072 -7945 -2038
rect -7855 -2072 -7787 -2038
rect -7697 -2072 -7629 -2038
rect -7539 -2072 -7471 -2038
rect -7381 -2072 -7313 -2038
rect -7223 -2072 -7155 -2038
rect -7065 -2072 -6997 -2038
rect -6907 -2072 -6839 -2038
rect -6749 -2072 -6681 -2038
rect -6591 -2072 -6523 -2038
rect -6433 -2072 -6365 -2038
rect -6275 -2072 -6207 -2038
rect -6117 -2072 -6049 -2038
rect -5959 -2072 -5891 -2038
rect -5801 -2072 -5733 -2038
rect -5643 -2072 -5575 -2038
rect -5485 -2072 -5417 -2038
rect -5327 -2072 -5259 -2038
rect -5169 -2072 -5101 -2038
rect -5011 -2072 -4943 -2038
rect -4853 -2072 -4785 -2038
rect -4695 -2072 -4627 -2038
rect -4537 -2072 -4469 -2038
rect -4379 -2072 -4311 -2038
rect -4221 -2072 -4153 -2038
rect -4063 -2072 -3995 -2038
rect -3905 -2072 -3837 -2038
rect -3747 -2072 -3679 -2038
rect -3589 -2072 -3521 -2038
rect -3431 -2072 -3363 -2038
rect -3273 -2072 -3205 -2038
rect -3115 -2072 -3047 -2038
rect -2957 -2072 -2889 -2038
rect -2799 -2072 -2731 -2038
rect -2641 -2072 -2573 -2038
rect -2483 -2072 -2415 -2038
rect -2325 -2072 -2257 -2038
rect -2167 -2072 -2099 -2038
rect -2009 -2072 -1941 -2038
rect -1851 -2072 -1783 -2038
rect -1693 -2072 -1625 -2038
rect -1535 -2072 -1467 -2038
rect -1377 -2072 -1309 -2038
rect -1219 -2072 -1151 -2038
rect -1061 -2072 -993 -2038
rect -903 -2072 -835 -2038
rect -745 -2072 -677 -2038
rect -587 -2072 -519 -2038
rect -429 -2072 -361 -2038
rect -271 -2072 -203 -2038
rect -113 -2072 -45 -2038
rect 45 -2072 113 -2038
rect 203 -2072 271 -2038
rect 361 -2072 429 -2038
rect 519 -2072 587 -2038
rect 677 -2072 745 -2038
rect 835 -2072 903 -2038
rect 993 -2072 1061 -2038
rect 1151 -2072 1219 -2038
rect 1309 -2072 1377 -2038
rect 1467 -2072 1535 -2038
rect 1625 -2072 1693 -2038
rect 1783 -2072 1851 -2038
rect 1941 -2072 2009 -2038
rect 2099 -2072 2167 -2038
rect 2257 -2072 2325 -2038
rect 2415 -2072 2483 -2038
rect 2573 -2072 2641 -2038
rect 2731 -2072 2799 -2038
rect 2889 -2072 2957 -2038
rect 3047 -2072 3115 -2038
rect 3205 -2072 3273 -2038
rect 3363 -2072 3431 -2038
rect 3521 -2072 3589 -2038
rect 3679 -2072 3747 -2038
rect 3837 -2072 3905 -2038
rect 3995 -2072 4063 -2038
rect 4153 -2072 4221 -2038
rect 4311 -2072 4379 -2038
rect 4469 -2072 4537 -2038
rect 4627 -2072 4695 -2038
rect 4785 -2072 4853 -2038
rect 4943 -2072 5011 -2038
rect 5101 -2072 5169 -2038
rect 5259 -2072 5327 -2038
rect 5417 -2072 5485 -2038
rect 5575 -2072 5643 -2038
rect 5733 -2072 5801 -2038
rect 5891 -2072 5959 -2038
rect 6049 -2072 6117 -2038
rect 6207 -2072 6275 -2038
rect 6365 -2072 6433 -2038
rect 6523 -2072 6591 -2038
rect 6681 -2072 6749 -2038
rect 6839 -2072 6907 -2038
rect 6997 -2072 7065 -2038
rect 7155 -2072 7223 -2038
rect 7313 -2072 7381 -2038
rect 7471 -2072 7539 -2038
rect 7629 -2072 7697 -2038
rect 7787 -2072 7855 -2038
rect 7945 -2072 8013 -2038
rect 8103 -2072 8171 -2038
rect 8261 -2072 8329 -2038
rect 8419 -2072 8487 -2038
rect 8577 -2072 8645 -2038
rect 8735 -2072 8803 -2038
rect 8893 -2072 8961 -2038
rect 9051 -2072 9119 -2038
rect 9209 -2072 9277 -2038
rect 9367 -2072 9435 -2038
rect 9525 -2072 9593 -2038
rect 9683 -2072 9751 -2038
rect 9841 -2072 9909 -2038
rect 9999 -2072 10067 -2038
<< locali >>
rect -10263 2176 -10167 2210
rect 10167 2176 10263 2210
rect -10263 2114 -10229 2176
rect 10229 2114 10263 2176
rect -10083 2038 -10067 2072
rect -9999 2038 -9983 2072
rect -9925 2038 -9909 2072
rect -9841 2038 -9825 2072
rect -9767 2038 -9751 2072
rect -9683 2038 -9667 2072
rect -9609 2038 -9593 2072
rect -9525 2038 -9509 2072
rect -9451 2038 -9435 2072
rect -9367 2038 -9351 2072
rect -9293 2038 -9277 2072
rect -9209 2038 -9193 2072
rect -9135 2038 -9119 2072
rect -9051 2038 -9035 2072
rect -8977 2038 -8961 2072
rect -8893 2038 -8877 2072
rect -8819 2038 -8803 2072
rect -8735 2038 -8719 2072
rect -8661 2038 -8645 2072
rect -8577 2038 -8561 2072
rect -8503 2038 -8487 2072
rect -8419 2038 -8403 2072
rect -8345 2038 -8329 2072
rect -8261 2038 -8245 2072
rect -8187 2038 -8171 2072
rect -8103 2038 -8087 2072
rect -8029 2038 -8013 2072
rect -7945 2038 -7929 2072
rect -7871 2038 -7855 2072
rect -7787 2038 -7771 2072
rect -7713 2038 -7697 2072
rect -7629 2038 -7613 2072
rect -7555 2038 -7539 2072
rect -7471 2038 -7455 2072
rect -7397 2038 -7381 2072
rect -7313 2038 -7297 2072
rect -7239 2038 -7223 2072
rect -7155 2038 -7139 2072
rect -7081 2038 -7065 2072
rect -6997 2038 -6981 2072
rect -6923 2038 -6907 2072
rect -6839 2038 -6823 2072
rect -6765 2038 -6749 2072
rect -6681 2038 -6665 2072
rect -6607 2038 -6591 2072
rect -6523 2038 -6507 2072
rect -6449 2038 -6433 2072
rect -6365 2038 -6349 2072
rect -6291 2038 -6275 2072
rect -6207 2038 -6191 2072
rect -6133 2038 -6117 2072
rect -6049 2038 -6033 2072
rect -5975 2038 -5959 2072
rect -5891 2038 -5875 2072
rect -5817 2038 -5801 2072
rect -5733 2038 -5717 2072
rect -5659 2038 -5643 2072
rect -5575 2038 -5559 2072
rect -5501 2038 -5485 2072
rect -5417 2038 -5401 2072
rect -5343 2038 -5327 2072
rect -5259 2038 -5243 2072
rect -5185 2038 -5169 2072
rect -5101 2038 -5085 2072
rect -5027 2038 -5011 2072
rect -4943 2038 -4927 2072
rect -4869 2038 -4853 2072
rect -4785 2038 -4769 2072
rect -4711 2038 -4695 2072
rect -4627 2038 -4611 2072
rect -4553 2038 -4537 2072
rect -4469 2038 -4453 2072
rect -4395 2038 -4379 2072
rect -4311 2038 -4295 2072
rect -4237 2038 -4221 2072
rect -4153 2038 -4137 2072
rect -4079 2038 -4063 2072
rect -3995 2038 -3979 2072
rect -3921 2038 -3905 2072
rect -3837 2038 -3821 2072
rect -3763 2038 -3747 2072
rect -3679 2038 -3663 2072
rect -3605 2038 -3589 2072
rect -3521 2038 -3505 2072
rect -3447 2038 -3431 2072
rect -3363 2038 -3347 2072
rect -3289 2038 -3273 2072
rect -3205 2038 -3189 2072
rect -3131 2038 -3115 2072
rect -3047 2038 -3031 2072
rect -2973 2038 -2957 2072
rect -2889 2038 -2873 2072
rect -2815 2038 -2799 2072
rect -2731 2038 -2715 2072
rect -2657 2038 -2641 2072
rect -2573 2038 -2557 2072
rect -2499 2038 -2483 2072
rect -2415 2038 -2399 2072
rect -2341 2038 -2325 2072
rect -2257 2038 -2241 2072
rect -2183 2038 -2167 2072
rect -2099 2038 -2083 2072
rect -2025 2038 -2009 2072
rect -1941 2038 -1925 2072
rect -1867 2038 -1851 2072
rect -1783 2038 -1767 2072
rect -1709 2038 -1693 2072
rect -1625 2038 -1609 2072
rect -1551 2038 -1535 2072
rect -1467 2038 -1451 2072
rect -1393 2038 -1377 2072
rect -1309 2038 -1293 2072
rect -1235 2038 -1219 2072
rect -1151 2038 -1135 2072
rect -1077 2038 -1061 2072
rect -993 2038 -977 2072
rect -919 2038 -903 2072
rect -835 2038 -819 2072
rect -761 2038 -745 2072
rect -677 2038 -661 2072
rect -603 2038 -587 2072
rect -519 2038 -503 2072
rect -445 2038 -429 2072
rect -361 2038 -345 2072
rect -287 2038 -271 2072
rect -203 2038 -187 2072
rect -129 2038 -113 2072
rect -45 2038 -29 2072
rect 29 2038 45 2072
rect 113 2038 129 2072
rect 187 2038 203 2072
rect 271 2038 287 2072
rect 345 2038 361 2072
rect 429 2038 445 2072
rect 503 2038 519 2072
rect 587 2038 603 2072
rect 661 2038 677 2072
rect 745 2038 761 2072
rect 819 2038 835 2072
rect 903 2038 919 2072
rect 977 2038 993 2072
rect 1061 2038 1077 2072
rect 1135 2038 1151 2072
rect 1219 2038 1235 2072
rect 1293 2038 1309 2072
rect 1377 2038 1393 2072
rect 1451 2038 1467 2072
rect 1535 2038 1551 2072
rect 1609 2038 1625 2072
rect 1693 2038 1709 2072
rect 1767 2038 1783 2072
rect 1851 2038 1867 2072
rect 1925 2038 1941 2072
rect 2009 2038 2025 2072
rect 2083 2038 2099 2072
rect 2167 2038 2183 2072
rect 2241 2038 2257 2072
rect 2325 2038 2341 2072
rect 2399 2038 2415 2072
rect 2483 2038 2499 2072
rect 2557 2038 2573 2072
rect 2641 2038 2657 2072
rect 2715 2038 2731 2072
rect 2799 2038 2815 2072
rect 2873 2038 2889 2072
rect 2957 2038 2973 2072
rect 3031 2038 3047 2072
rect 3115 2038 3131 2072
rect 3189 2038 3205 2072
rect 3273 2038 3289 2072
rect 3347 2038 3363 2072
rect 3431 2038 3447 2072
rect 3505 2038 3521 2072
rect 3589 2038 3605 2072
rect 3663 2038 3679 2072
rect 3747 2038 3763 2072
rect 3821 2038 3837 2072
rect 3905 2038 3921 2072
rect 3979 2038 3995 2072
rect 4063 2038 4079 2072
rect 4137 2038 4153 2072
rect 4221 2038 4237 2072
rect 4295 2038 4311 2072
rect 4379 2038 4395 2072
rect 4453 2038 4469 2072
rect 4537 2038 4553 2072
rect 4611 2038 4627 2072
rect 4695 2038 4711 2072
rect 4769 2038 4785 2072
rect 4853 2038 4869 2072
rect 4927 2038 4943 2072
rect 5011 2038 5027 2072
rect 5085 2038 5101 2072
rect 5169 2038 5185 2072
rect 5243 2038 5259 2072
rect 5327 2038 5343 2072
rect 5401 2038 5417 2072
rect 5485 2038 5501 2072
rect 5559 2038 5575 2072
rect 5643 2038 5659 2072
rect 5717 2038 5733 2072
rect 5801 2038 5817 2072
rect 5875 2038 5891 2072
rect 5959 2038 5975 2072
rect 6033 2038 6049 2072
rect 6117 2038 6133 2072
rect 6191 2038 6207 2072
rect 6275 2038 6291 2072
rect 6349 2038 6365 2072
rect 6433 2038 6449 2072
rect 6507 2038 6523 2072
rect 6591 2038 6607 2072
rect 6665 2038 6681 2072
rect 6749 2038 6765 2072
rect 6823 2038 6839 2072
rect 6907 2038 6923 2072
rect 6981 2038 6997 2072
rect 7065 2038 7081 2072
rect 7139 2038 7155 2072
rect 7223 2038 7239 2072
rect 7297 2038 7313 2072
rect 7381 2038 7397 2072
rect 7455 2038 7471 2072
rect 7539 2038 7555 2072
rect 7613 2038 7629 2072
rect 7697 2038 7713 2072
rect 7771 2038 7787 2072
rect 7855 2038 7871 2072
rect 7929 2038 7945 2072
rect 8013 2038 8029 2072
rect 8087 2038 8103 2072
rect 8171 2038 8187 2072
rect 8245 2038 8261 2072
rect 8329 2038 8345 2072
rect 8403 2038 8419 2072
rect 8487 2038 8503 2072
rect 8561 2038 8577 2072
rect 8645 2038 8661 2072
rect 8719 2038 8735 2072
rect 8803 2038 8819 2072
rect 8877 2038 8893 2072
rect 8961 2038 8977 2072
rect 9035 2038 9051 2072
rect 9119 2038 9135 2072
rect 9193 2038 9209 2072
rect 9277 2038 9293 2072
rect 9351 2038 9367 2072
rect 9435 2038 9451 2072
rect 9509 2038 9525 2072
rect 9593 2038 9609 2072
rect 9667 2038 9683 2072
rect 9751 2038 9767 2072
rect 9825 2038 9841 2072
rect 9909 2038 9925 2072
rect 9983 2038 9999 2072
rect 10067 2038 10083 2072
rect -10129 1988 -10095 2004
rect -10129 -2004 -10095 -1988
rect -9971 1988 -9937 2004
rect -9971 -2004 -9937 -1988
rect -9813 1988 -9779 2004
rect -9813 -2004 -9779 -1988
rect -9655 1988 -9621 2004
rect -9655 -2004 -9621 -1988
rect -9497 1988 -9463 2004
rect -9497 -2004 -9463 -1988
rect -9339 1988 -9305 2004
rect -9339 -2004 -9305 -1988
rect -9181 1988 -9147 2004
rect -9181 -2004 -9147 -1988
rect -9023 1988 -8989 2004
rect -9023 -2004 -8989 -1988
rect -8865 1988 -8831 2004
rect -8865 -2004 -8831 -1988
rect -8707 1988 -8673 2004
rect -8707 -2004 -8673 -1988
rect -8549 1988 -8515 2004
rect -8549 -2004 -8515 -1988
rect -8391 1988 -8357 2004
rect -8391 -2004 -8357 -1988
rect -8233 1988 -8199 2004
rect -8233 -2004 -8199 -1988
rect -8075 1988 -8041 2004
rect -8075 -2004 -8041 -1988
rect -7917 1988 -7883 2004
rect -7917 -2004 -7883 -1988
rect -7759 1988 -7725 2004
rect -7759 -2004 -7725 -1988
rect -7601 1988 -7567 2004
rect -7601 -2004 -7567 -1988
rect -7443 1988 -7409 2004
rect -7443 -2004 -7409 -1988
rect -7285 1988 -7251 2004
rect -7285 -2004 -7251 -1988
rect -7127 1988 -7093 2004
rect -7127 -2004 -7093 -1988
rect -6969 1988 -6935 2004
rect -6969 -2004 -6935 -1988
rect -6811 1988 -6777 2004
rect -6811 -2004 -6777 -1988
rect -6653 1988 -6619 2004
rect -6653 -2004 -6619 -1988
rect -6495 1988 -6461 2004
rect -6495 -2004 -6461 -1988
rect -6337 1988 -6303 2004
rect -6337 -2004 -6303 -1988
rect -6179 1988 -6145 2004
rect -6179 -2004 -6145 -1988
rect -6021 1988 -5987 2004
rect -6021 -2004 -5987 -1988
rect -5863 1988 -5829 2004
rect -5863 -2004 -5829 -1988
rect -5705 1988 -5671 2004
rect -5705 -2004 -5671 -1988
rect -5547 1988 -5513 2004
rect -5547 -2004 -5513 -1988
rect -5389 1988 -5355 2004
rect -5389 -2004 -5355 -1988
rect -5231 1988 -5197 2004
rect -5231 -2004 -5197 -1988
rect -5073 1988 -5039 2004
rect -5073 -2004 -5039 -1988
rect -4915 1988 -4881 2004
rect -4915 -2004 -4881 -1988
rect -4757 1988 -4723 2004
rect -4757 -2004 -4723 -1988
rect -4599 1988 -4565 2004
rect -4599 -2004 -4565 -1988
rect -4441 1988 -4407 2004
rect -4441 -2004 -4407 -1988
rect -4283 1988 -4249 2004
rect -4283 -2004 -4249 -1988
rect -4125 1988 -4091 2004
rect -4125 -2004 -4091 -1988
rect -3967 1988 -3933 2004
rect -3967 -2004 -3933 -1988
rect -3809 1988 -3775 2004
rect -3809 -2004 -3775 -1988
rect -3651 1988 -3617 2004
rect -3651 -2004 -3617 -1988
rect -3493 1988 -3459 2004
rect -3493 -2004 -3459 -1988
rect -3335 1988 -3301 2004
rect -3335 -2004 -3301 -1988
rect -3177 1988 -3143 2004
rect -3177 -2004 -3143 -1988
rect -3019 1988 -2985 2004
rect -3019 -2004 -2985 -1988
rect -2861 1988 -2827 2004
rect -2861 -2004 -2827 -1988
rect -2703 1988 -2669 2004
rect -2703 -2004 -2669 -1988
rect -2545 1988 -2511 2004
rect -2545 -2004 -2511 -1988
rect -2387 1988 -2353 2004
rect -2387 -2004 -2353 -1988
rect -2229 1988 -2195 2004
rect -2229 -2004 -2195 -1988
rect -2071 1988 -2037 2004
rect -2071 -2004 -2037 -1988
rect -1913 1988 -1879 2004
rect -1913 -2004 -1879 -1988
rect -1755 1988 -1721 2004
rect -1755 -2004 -1721 -1988
rect -1597 1988 -1563 2004
rect -1597 -2004 -1563 -1988
rect -1439 1988 -1405 2004
rect -1439 -2004 -1405 -1988
rect -1281 1988 -1247 2004
rect -1281 -2004 -1247 -1988
rect -1123 1988 -1089 2004
rect -1123 -2004 -1089 -1988
rect -965 1988 -931 2004
rect -965 -2004 -931 -1988
rect -807 1988 -773 2004
rect -807 -2004 -773 -1988
rect -649 1988 -615 2004
rect -649 -2004 -615 -1988
rect -491 1988 -457 2004
rect -491 -2004 -457 -1988
rect -333 1988 -299 2004
rect -333 -2004 -299 -1988
rect -175 1988 -141 2004
rect -175 -2004 -141 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 141 1988 175 2004
rect 141 -2004 175 -1988
rect 299 1988 333 2004
rect 299 -2004 333 -1988
rect 457 1988 491 2004
rect 457 -2004 491 -1988
rect 615 1988 649 2004
rect 615 -2004 649 -1988
rect 773 1988 807 2004
rect 773 -2004 807 -1988
rect 931 1988 965 2004
rect 931 -2004 965 -1988
rect 1089 1988 1123 2004
rect 1089 -2004 1123 -1988
rect 1247 1988 1281 2004
rect 1247 -2004 1281 -1988
rect 1405 1988 1439 2004
rect 1405 -2004 1439 -1988
rect 1563 1988 1597 2004
rect 1563 -2004 1597 -1988
rect 1721 1988 1755 2004
rect 1721 -2004 1755 -1988
rect 1879 1988 1913 2004
rect 1879 -2004 1913 -1988
rect 2037 1988 2071 2004
rect 2037 -2004 2071 -1988
rect 2195 1988 2229 2004
rect 2195 -2004 2229 -1988
rect 2353 1988 2387 2004
rect 2353 -2004 2387 -1988
rect 2511 1988 2545 2004
rect 2511 -2004 2545 -1988
rect 2669 1988 2703 2004
rect 2669 -2004 2703 -1988
rect 2827 1988 2861 2004
rect 2827 -2004 2861 -1988
rect 2985 1988 3019 2004
rect 2985 -2004 3019 -1988
rect 3143 1988 3177 2004
rect 3143 -2004 3177 -1988
rect 3301 1988 3335 2004
rect 3301 -2004 3335 -1988
rect 3459 1988 3493 2004
rect 3459 -2004 3493 -1988
rect 3617 1988 3651 2004
rect 3617 -2004 3651 -1988
rect 3775 1988 3809 2004
rect 3775 -2004 3809 -1988
rect 3933 1988 3967 2004
rect 3933 -2004 3967 -1988
rect 4091 1988 4125 2004
rect 4091 -2004 4125 -1988
rect 4249 1988 4283 2004
rect 4249 -2004 4283 -1988
rect 4407 1988 4441 2004
rect 4407 -2004 4441 -1988
rect 4565 1988 4599 2004
rect 4565 -2004 4599 -1988
rect 4723 1988 4757 2004
rect 4723 -2004 4757 -1988
rect 4881 1988 4915 2004
rect 4881 -2004 4915 -1988
rect 5039 1988 5073 2004
rect 5039 -2004 5073 -1988
rect 5197 1988 5231 2004
rect 5197 -2004 5231 -1988
rect 5355 1988 5389 2004
rect 5355 -2004 5389 -1988
rect 5513 1988 5547 2004
rect 5513 -2004 5547 -1988
rect 5671 1988 5705 2004
rect 5671 -2004 5705 -1988
rect 5829 1988 5863 2004
rect 5829 -2004 5863 -1988
rect 5987 1988 6021 2004
rect 5987 -2004 6021 -1988
rect 6145 1988 6179 2004
rect 6145 -2004 6179 -1988
rect 6303 1988 6337 2004
rect 6303 -2004 6337 -1988
rect 6461 1988 6495 2004
rect 6461 -2004 6495 -1988
rect 6619 1988 6653 2004
rect 6619 -2004 6653 -1988
rect 6777 1988 6811 2004
rect 6777 -2004 6811 -1988
rect 6935 1988 6969 2004
rect 6935 -2004 6969 -1988
rect 7093 1988 7127 2004
rect 7093 -2004 7127 -1988
rect 7251 1988 7285 2004
rect 7251 -2004 7285 -1988
rect 7409 1988 7443 2004
rect 7409 -2004 7443 -1988
rect 7567 1988 7601 2004
rect 7567 -2004 7601 -1988
rect 7725 1988 7759 2004
rect 7725 -2004 7759 -1988
rect 7883 1988 7917 2004
rect 7883 -2004 7917 -1988
rect 8041 1988 8075 2004
rect 8041 -2004 8075 -1988
rect 8199 1988 8233 2004
rect 8199 -2004 8233 -1988
rect 8357 1988 8391 2004
rect 8357 -2004 8391 -1988
rect 8515 1988 8549 2004
rect 8515 -2004 8549 -1988
rect 8673 1988 8707 2004
rect 8673 -2004 8707 -1988
rect 8831 1988 8865 2004
rect 8831 -2004 8865 -1988
rect 8989 1988 9023 2004
rect 8989 -2004 9023 -1988
rect 9147 1988 9181 2004
rect 9147 -2004 9181 -1988
rect 9305 1988 9339 2004
rect 9305 -2004 9339 -1988
rect 9463 1988 9497 2004
rect 9463 -2004 9497 -1988
rect 9621 1988 9655 2004
rect 9621 -2004 9655 -1988
rect 9779 1988 9813 2004
rect 9779 -2004 9813 -1988
rect 9937 1988 9971 2004
rect 9937 -2004 9971 -1988
rect 10095 1988 10129 2004
rect 10095 -2004 10129 -1988
rect -10083 -2072 -10067 -2038
rect -9999 -2072 -9983 -2038
rect -9925 -2072 -9909 -2038
rect -9841 -2072 -9825 -2038
rect -9767 -2072 -9751 -2038
rect -9683 -2072 -9667 -2038
rect -9609 -2072 -9593 -2038
rect -9525 -2072 -9509 -2038
rect -9451 -2072 -9435 -2038
rect -9367 -2072 -9351 -2038
rect -9293 -2072 -9277 -2038
rect -9209 -2072 -9193 -2038
rect -9135 -2072 -9119 -2038
rect -9051 -2072 -9035 -2038
rect -8977 -2072 -8961 -2038
rect -8893 -2072 -8877 -2038
rect -8819 -2072 -8803 -2038
rect -8735 -2072 -8719 -2038
rect -8661 -2072 -8645 -2038
rect -8577 -2072 -8561 -2038
rect -8503 -2072 -8487 -2038
rect -8419 -2072 -8403 -2038
rect -8345 -2072 -8329 -2038
rect -8261 -2072 -8245 -2038
rect -8187 -2072 -8171 -2038
rect -8103 -2072 -8087 -2038
rect -8029 -2072 -8013 -2038
rect -7945 -2072 -7929 -2038
rect -7871 -2072 -7855 -2038
rect -7787 -2072 -7771 -2038
rect -7713 -2072 -7697 -2038
rect -7629 -2072 -7613 -2038
rect -7555 -2072 -7539 -2038
rect -7471 -2072 -7455 -2038
rect -7397 -2072 -7381 -2038
rect -7313 -2072 -7297 -2038
rect -7239 -2072 -7223 -2038
rect -7155 -2072 -7139 -2038
rect -7081 -2072 -7065 -2038
rect -6997 -2072 -6981 -2038
rect -6923 -2072 -6907 -2038
rect -6839 -2072 -6823 -2038
rect -6765 -2072 -6749 -2038
rect -6681 -2072 -6665 -2038
rect -6607 -2072 -6591 -2038
rect -6523 -2072 -6507 -2038
rect -6449 -2072 -6433 -2038
rect -6365 -2072 -6349 -2038
rect -6291 -2072 -6275 -2038
rect -6207 -2072 -6191 -2038
rect -6133 -2072 -6117 -2038
rect -6049 -2072 -6033 -2038
rect -5975 -2072 -5959 -2038
rect -5891 -2072 -5875 -2038
rect -5817 -2072 -5801 -2038
rect -5733 -2072 -5717 -2038
rect -5659 -2072 -5643 -2038
rect -5575 -2072 -5559 -2038
rect -5501 -2072 -5485 -2038
rect -5417 -2072 -5401 -2038
rect -5343 -2072 -5327 -2038
rect -5259 -2072 -5243 -2038
rect -5185 -2072 -5169 -2038
rect -5101 -2072 -5085 -2038
rect -5027 -2072 -5011 -2038
rect -4943 -2072 -4927 -2038
rect -4869 -2072 -4853 -2038
rect -4785 -2072 -4769 -2038
rect -4711 -2072 -4695 -2038
rect -4627 -2072 -4611 -2038
rect -4553 -2072 -4537 -2038
rect -4469 -2072 -4453 -2038
rect -4395 -2072 -4379 -2038
rect -4311 -2072 -4295 -2038
rect -4237 -2072 -4221 -2038
rect -4153 -2072 -4137 -2038
rect -4079 -2072 -4063 -2038
rect -3995 -2072 -3979 -2038
rect -3921 -2072 -3905 -2038
rect -3837 -2072 -3821 -2038
rect -3763 -2072 -3747 -2038
rect -3679 -2072 -3663 -2038
rect -3605 -2072 -3589 -2038
rect -3521 -2072 -3505 -2038
rect -3447 -2072 -3431 -2038
rect -3363 -2072 -3347 -2038
rect -3289 -2072 -3273 -2038
rect -3205 -2072 -3189 -2038
rect -3131 -2072 -3115 -2038
rect -3047 -2072 -3031 -2038
rect -2973 -2072 -2957 -2038
rect -2889 -2072 -2873 -2038
rect -2815 -2072 -2799 -2038
rect -2731 -2072 -2715 -2038
rect -2657 -2072 -2641 -2038
rect -2573 -2072 -2557 -2038
rect -2499 -2072 -2483 -2038
rect -2415 -2072 -2399 -2038
rect -2341 -2072 -2325 -2038
rect -2257 -2072 -2241 -2038
rect -2183 -2072 -2167 -2038
rect -2099 -2072 -2083 -2038
rect -2025 -2072 -2009 -2038
rect -1941 -2072 -1925 -2038
rect -1867 -2072 -1851 -2038
rect -1783 -2072 -1767 -2038
rect -1709 -2072 -1693 -2038
rect -1625 -2072 -1609 -2038
rect -1551 -2072 -1535 -2038
rect -1467 -2072 -1451 -2038
rect -1393 -2072 -1377 -2038
rect -1309 -2072 -1293 -2038
rect -1235 -2072 -1219 -2038
rect -1151 -2072 -1135 -2038
rect -1077 -2072 -1061 -2038
rect -993 -2072 -977 -2038
rect -919 -2072 -903 -2038
rect -835 -2072 -819 -2038
rect -761 -2072 -745 -2038
rect -677 -2072 -661 -2038
rect -603 -2072 -587 -2038
rect -519 -2072 -503 -2038
rect -445 -2072 -429 -2038
rect -361 -2072 -345 -2038
rect -287 -2072 -271 -2038
rect -203 -2072 -187 -2038
rect -129 -2072 -113 -2038
rect -45 -2072 -29 -2038
rect 29 -2072 45 -2038
rect 113 -2072 129 -2038
rect 187 -2072 203 -2038
rect 271 -2072 287 -2038
rect 345 -2072 361 -2038
rect 429 -2072 445 -2038
rect 503 -2072 519 -2038
rect 587 -2072 603 -2038
rect 661 -2072 677 -2038
rect 745 -2072 761 -2038
rect 819 -2072 835 -2038
rect 903 -2072 919 -2038
rect 977 -2072 993 -2038
rect 1061 -2072 1077 -2038
rect 1135 -2072 1151 -2038
rect 1219 -2072 1235 -2038
rect 1293 -2072 1309 -2038
rect 1377 -2072 1393 -2038
rect 1451 -2072 1467 -2038
rect 1535 -2072 1551 -2038
rect 1609 -2072 1625 -2038
rect 1693 -2072 1709 -2038
rect 1767 -2072 1783 -2038
rect 1851 -2072 1867 -2038
rect 1925 -2072 1941 -2038
rect 2009 -2072 2025 -2038
rect 2083 -2072 2099 -2038
rect 2167 -2072 2183 -2038
rect 2241 -2072 2257 -2038
rect 2325 -2072 2341 -2038
rect 2399 -2072 2415 -2038
rect 2483 -2072 2499 -2038
rect 2557 -2072 2573 -2038
rect 2641 -2072 2657 -2038
rect 2715 -2072 2731 -2038
rect 2799 -2072 2815 -2038
rect 2873 -2072 2889 -2038
rect 2957 -2072 2973 -2038
rect 3031 -2072 3047 -2038
rect 3115 -2072 3131 -2038
rect 3189 -2072 3205 -2038
rect 3273 -2072 3289 -2038
rect 3347 -2072 3363 -2038
rect 3431 -2072 3447 -2038
rect 3505 -2072 3521 -2038
rect 3589 -2072 3605 -2038
rect 3663 -2072 3679 -2038
rect 3747 -2072 3763 -2038
rect 3821 -2072 3837 -2038
rect 3905 -2072 3921 -2038
rect 3979 -2072 3995 -2038
rect 4063 -2072 4079 -2038
rect 4137 -2072 4153 -2038
rect 4221 -2072 4237 -2038
rect 4295 -2072 4311 -2038
rect 4379 -2072 4395 -2038
rect 4453 -2072 4469 -2038
rect 4537 -2072 4553 -2038
rect 4611 -2072 4627 -2038
rect 4695 -2072 4711 -2038
rect 4769 -2072 4785 -2038
rect 4853 -2072 4869 -2038
rect 4927 -2072 4943 -2038
rect 5011 -2072 5027 -2038
rect 5085 -2072 5101 -2038
rect 5169 -2072 5185 -2038
rect 5243 -2072 5259 -2038
rect 5327 -2072 5343 -2038
rect 5401 -2072 5417 -2038
rect 5485 -2072 5501 -2038
rect 5559 -2072 5575 -2038
rect 5643 -2072 5659 -2038
rect 5717 -2072 5733 -2038
rect 5801 -2072 5817 -2038
rect 5875 -2072 5891 -2038
rect 5959 -2072 5975 -2038
rect 6033 -2072 6049 -2038
rect 6117 -2072 6133 -2038
rect 6191 -2072 6207 -2038
rect 6275 -2072 6291 -2038
rect 6349 -2072 6365 -2038
rect 6433 -2072 6449 -2038
rect 6507 -2072 6523 -2038
rect 6591 -2072 6607 -2038
rect 6665 -2072 6681 -2038
rect 6749 -2072 6765 -2038
rect 6823 -2072 6839 -2038
rect 6907 -2072 6923 -2038
rect 6981 -2072 6997 -2038
rect 7065 -2072 7081 -2038
rect 7139 -2072 7155 -2038
rect 7223 -2072 7239 -2038
rect 7297 -2072 7313 -2038
rect 7381 -2072 7397 -2038
rect 7455 -2072 7471 -2038
rect 7539 -2072 7555 -2038
rect 7613 -2072 7629 -2038
rect 7697 -2072 7713 -2038
rect 7771 -2072 7787 -2038
rect 7855 -2072 7871 -2038
rect 7929 -2072 7945 -2038
rect 8013 -2072 8029 -2038
rect 8087 -2072 8103 -2038
rect 8171 -2072 8187 -2038
rect 8245 -2072 8261 -2038
rect 8329 -2072 8345 -2038
rect 8403 -2072 8419 -2038
rect 8487 -2072 8503 -2038
rect 8561 -2072 8577 -2038
rect 8645 -2072 8661 -2038
rect 8719 -2072 8735 -2038
rect 8803 -2072 8819 -2038
rect 8877 -2072 8893 -2038
rect 8961 -2072 8977 -2038
rect 9035 -2072 9051 -2038
rect 9119 -2072 9135 -2038
rect 9193 -2072 9209 -2038
rect 9277 -2072 9293 -2038
rect 9351 -2072 9367 -2038
rect 9435 -2072 9451 -2038
rect 9509 -2072 9525 -2038
rect 9593 -2072 9609 -2038
rect 9667 -2072 9683 -2038
rect 9751 -2072 9767 -2038
rect 9825 -2072 9841 -2038
rect 9909 -2072 9925 -2038
rect 9983 -2072 9999 -2038
rect 10067 -2072 10083 -2038
rect -10263 -2176 -10229 -2114
rect 10229 -2176 10263 -2114
rect -10263 -2210 -10167 -2176
rect 10167 -2210 10263 -2176
<< viali >>
rect -10067 2038 -9999 2072
rect -9909 2038 -9841 2072
rect -9751 2038 -9683 2072
rect -9593 2038 -9525 2072
rect -9435 2038 -9367 2072
rect -9277 2038 -9209 2072
rect -9119 2038 -9051 2072
rect -8961 2038 -8893 2072
rect -8803 2038 -8735 2072
rect -8645 2038 -8577 2072
rect -8487 2038 -8419 2072
rect -8329 2038 -8261 2072
rect -8171 2038 -8103 2072
rect -8013 2038 -7945 2072
rect -7855 2038 -7787 2072
rect -7697 2038 -7629 2072
rect -7539 2038 -7471 2072
rect -7381 2038 -7313 2072
rect -7223 2038 -7155 2072
rect -7065 2038 -6997 2072
rect -6907 2038 -6839 2072
rect -6749 2038 -6681 2072
rect -6591 2038 -6523 2072
rect -6433 2038 -6365 2072
rect -6275 2038 -6207 2072
rect -6117 2038 -6049 2072
rect -5959 2038 -5891 2072
rect -5801 2038 -5733 2072
rect -5643 2038 -5575 2072
rect -5485 2038 -5417 2072
rect -5327 2038 -5259 2072
rect -5169 2038 -5101 2072
rect -5011 2038 -4943 2072
rect -4853 2038 -4785 2072
rect -4695 2038 -4627 2072
rect -4537 2038 -4469 2072
rect -4379 2038 -4311 2072
rect -4221 2038 -4153 2072
rect -4063 2038 -3995 2072
rect -3905 2038 -3837 2072
rect -3747 2038 -3679 2072
rect -3589 2038 -3521 2072
rect -3431 2038 -3363 2072
rect -3273 2038 -3205 2072
rect -3115 2038 -3047 2072
rect -2957 2038 -2889 2072
rect -2799 2038 -2731 2072
rect -2641 2038 -2573 2072
rect -2483 2038 -2415 2072
rect -2325 2038 -2257 2072
rect -2167 2038 -2099 2072
rect -2009 2038 -1941 2072
rect -1851 2038 -1783 2072
rect -1693 2038 -1625 2072
rect -1535 2038 -1467 2072
rect -1377 2038 -1309 2072
rect -1219 2038 -1151 2072
rect -1061 2038 -993 2072
rect -903 2038 -835 2072
rect -745 2038 -677 2072
rect -587 2038 -519 2072
rect -429 2038 -361 2072
rect -271 2038 -203 2072
rect -113 2038 -45 2072
rect 45 2038 113 2072
rect 203 2038 271 2072
rect 361 2038 429 2072
rect 519 2038 587 2072
rect 677 2038 745 2072
rect 835 2038 903 2072
rect 993 2038 1061 2072
rect 1151 2038 1219 2072
rect 1309 2038 1377 2072
rect 1467 2038 1535 2072
rect 1625 2038 1693 2072
rect 1783 2038 1851 2072
rect 1941 2038 2009 2072
rect 2099 2038 2167 2072
rect 2257 2038 2325 2072
rect 2415 2038 2483 2072
rect 2573 2038 2641 2072
rect 2731 2038 2799 2072
rect 2889 2038 2957 2072
rect 3047 2038 3115 2072
rect 3205 2038 3273 2072
rect 3363 2038 3431 2072
rect 3521 2038 3589 2072
rect 3679 2038 3747 2072
rect 3837 2038 3905 2072
rect 3995 2038 4063 2072
rect 4153 2038 4221 2072
rect 4311 2038 4379 2072
rect 4469 2038 4537 2072
rect 4627 2038 4695 2072
rect 4785 2038 4853 2072
rect 4943 2038 5011 2072
rect 5101 2038 5169 2072
rect 5259 2038 5327 2072
rect 5417 2038 5485 2072
rect 5575 2038 5643 2072
rect 5733 2038 5801 2072
rect 5891 2038 5959 2072
rect 6049 2038 6117 2072
rect 6207 2038 6275 2072
rect 6365 2038 6433 2072
rect 6523 2038 6591 2072
rect 6681 2038 6749 2072
rect 6839 2038 6907 2072
rect 6997 2038 7065 2072
rect 7155 2038 7223 2072
rect 7313 2038 7381 2072
rect 7471 2038 7539 2072
rect 7629 2038 7697 2072
rect 7787 2038 7855 2072
rect 7945 2038 8013 2072
rect 8103 2038 8171 2072
rect 8261 2038 8329 2072
rect 8419 2038 8487 2072
rect 8577 2038 8645 2072
rect 8735 2038 8803 2072
rect 8893 2038 8961 2072
rect 9051 2038 9119 2072
rect 9209 2038 9277 2072
rect 9367 2038 9435 2072
rect 9525 2038 9593 2072
rect 9683 2038 9751 2072
rect 9841 2038 9909 2072
rect 9999 2038 10067 2072
rect -10129 -1988 -10095 1988
rect -9971 -1988 -9937 1988
rect -9813 -1988 -9779 1988
rect -9655 -1988 -9621 1988
rect -9497 -1988 -9463 1988
rect -9339 -1988 -9305 1988
rect -9181 -1988 -9147 1988
rect -9023 -1988 -8989 1988
rect -8865 -1988 -8831 1988
rect -8707 -1988 -8673 1988
rect -8549 -1988 -8515 1988
rect -8391 -1988 -8357 1988
rect -8233 -1988 -8199 1988
rect -8075 -1988 -8041 1988
rect -7917 -1988 -7883 1988
rect -7759 -1988 -7725 1988
rect -7601 -1988 -7567 1988
rect -7443 -1988 -7409 1988
rect -7285 -1988 -7251 1988
rect -7127 -1988 -7093 1988
rect -6969 -1988 -6935 1988
rect -6811 -1988 -6777 1988
rect -6653 -1988 -6619 1988
rect -6495 -1988 -6461 1988
rect -6337 -1988 -6303 1988
rect -6179 -1988 -6145 1988
rect -6021 -1988 -5987 1988
rect -5863 -1988 -5829 1988
rect -5705 -1988 -5671 1988
rect -5547 -1988 -5513 1988
rect -5389 -1988 -5355 1988
rect -5231 -1988 -5197 1988
rect -5073 -1988 -5039 1988
rect -4915 -1988 -4881 1988
rect -4757 -1988 -4723 1988
rect -4599 -1988 -4565 1988
rect -4441 -1988 -4407 1988
rect -4283 -1988 -4249 1988
rect -4125 -1988 -4091 1988
rect -3967 -1988 -3933 1988
rect -3809 -1988 -3775 1988
rect -3651 -1988 -3617 1988
rect -3493 -1988 -3459 1988
rect -3335 -1988 -3301 1988
rect -3177 -1988 -3143 1988
rect -3019 -1988 -2985 1988
rect -2861 -1988 -2827 1988
rect -2703 -1988 -2669 1988
rect -2545 -1988 -2511 1988
rect -2387 -1988 -2353 1988
rect -2229 -1988 -2195 1988
rect -2071 -1988 -2037 1988
rect -1913 -1988 -1879 1988
rect -1755 -1988 -1721 1988
rect -1597 -1988 -1563 1988
rect -1439 -1988 -1405 1988
rect -1281 -1988 -1247 1988
rect -1123 -1988 -1089 1988
rect -965 -1988 -931 1988
rect -807 -1988 -773 1988
rect -649 -1988 -615 1988
rect -491 -1988 -457 1988
rect -333 -1988 -299 1988
rect -175 -1988 -141 1988
rect -17 -1988 17 1988
rect 141 -1988 175 1988
rect 299 -1988 333 1988
rect 457 -1988 491 1988
rect 615 -1988 649 1988
rect 773 -1988 807 1988
rect 931 -1988 965 1988
rect 1089 -1988 1123 1988
rect 1247 -1988 1281 1988
rect 1405 -1988 1439 1988
rect 1563 -1988 1597 1988
rect 1721 -1988 1755 1988
rect 1879 -1988 1913 1988
rect 2037 -1988 2071 1988
rect 2195 -1988 2229 1988
rect 2353 -1988 2387 1988
rect 2511 -1988 2545 1988
rect 2669 -1988 2703 1988
rect 2827 -1988 2861 1988
rect 2985 -1988 3019 1988
rect 3143 -1988 3177 1988
rect 3301 -1988 3335 1988
rect 3459 -1988 3493 1988
rect 3617 -1988 3651 1988
rect 3775 -1988 3809 1988
rect 3933 -1988 3967 1988
rect 4091 -1988 4125 1988
rect 4249 -1988 4283 1988
rect 4407 -1988 4441 1988
rect 4565 -1988 4599 1988
rect 4723 -1988 4757 1988
rect 4881 -1988 4915 1988
rect 5039 -1988 5073 1988
rect 5197 -1988 5231 1988
rect 5355 -1988 5389 1988
rect 5513 -1988 5547 1988
rect 5671 -1988 5705 1988
rect 5829 -1988 5863 1988
rect 5987 -1988 6021 1988
rect 6145 -1988 6179 1988
rect 6303 -1988 6337 1988
rect 6461 -1988 6495 1988
rect 6619 -1988 6653 1988
rect 6777 -1988 6811 1988
rect 6935 -1988 6969 1988
rect 7093 -1988 7127 1988
rect 7251 -1988 7285 1988
rect 7409 -1988 7443 1988
rect 7567 -1988 7601 1988
rect 7725 -1988 7759 1988
rect 7883 -1988 7917 1988
rect 8041 -1988 8075 1988
rect 8199 -1988 8233 1988
rect 8357 -1988 8391 1988
rect 8515 -1988 8549 1988
rect 8673 -1988 8707 1988
rect 8831 -1988 8865 1988
rect 8989 -1988 9023 1988
rect 9147 -1988 9181 1988
rect 9305 -1988 9339 1988
rect 9463 -1988 9497 1988
rect 9621 -1988 9655 1988
rect 9779 -1988 9813 1988
rect 9937 -1988 9971 1988
rect 10095 -1988 10129 1988
rect -10067 -2072 -9999 -2038
rect -9909 -2072 -9841 -2038
rect -9751 -2072 -9683 -2038
rect -9593 -2072 -9525 -2038
rect -9435 -2072 -9367 -2038
rect -9277 -2072 -9209 -2038
rect -9119 -2072 -9051 -2038
rect -8961 -2072 -8893 -2038
rect -8803 -2072 -8735 -2038
rect -8645 -2072 -8577 -2038
rect -8487 -2072 -8419 -2038
rect -8329 -2072 -8261 -2038
rect -8171 -2072 -8103 -2038
rect -8013 -2072 -7945 -2038
rect -7855 -2072 -7787 -2038
rect -7697 -2072 -7629 -2038
rect -7539 -2072 -7471 -2038
rect -7381 -2072 -7313 -2038
rect -7223 -2072 -7155 -2038
rect -7065 -2072 -6997 -2038
rect -6907 -2072 -6839 -2038
rect -6749 -2072 -6681 -2038
rect -6591 -2072 -6523 -2038
rect -6433 -2072 -6365 -2038
rect -6275 -2072 -6207 -2038
rect -6117 -2072 -6049 -2038
rect -5959 -2072 -5891 -2038
rect -5801 -2072 -5733 -2038
rect -5643 -2072 -5575 -2038
rect -5485 -2072 -5417 -2038
rect -5327 -2072 -5259 -2038
rect -5169 -2072 -5101 -2038
rect -5011 -2072 -4943 -2038
rect -4853 -2072 -4785 -2038
rect -4695 -2072 -4627 -2038
rect -4537 -2072 -4469 -2038
rect -4379 -2072 -4311 -2038
rect -4221 -2072 -4153 -2038
rect -4063 -2072 -3995 -2038
rect -3905 -2072 -3837 -2038
rect -3747 -2072 -3679 -2038
rect -3589 -2072 -3521 -2038
rect -3431 -2072 -3363 -2038
rect -3273 -2072 -3205 -2038
rect -3115 -2072 -3047 -2038
rect -2957 -2072 -2889 -2038
rect -2799 -2072 -2731 -2038
rect -2641 -2072 -2573 -2038
rect -2483 -2072 -2415 -2038
rect -2325 -2072 -2257 -2038
rect -2167 -2072 -2099 -2038
rect -2009 -2072 -1941 -2038
rect -1851 -2072 -1783 -2038
rect -1693 -2072 -1625 -2038
rect -1535 -2072 -1467 -2038
rect -1377 -2072 -1309 -2038
rect -1219 -2072 -1151 -2038
rect -1061 -2072 -993 -2038
rect -903 -2072 -835 -2038
rect -745 -2072 -677 -2038
rect -587 -2072 -519 -2038
rect -429 -2072 -361 -2038
rect -271 -2072 -203 -2038
rect -113 -2072 -45 -2038
rect 45 -2072 113 -2038
rect 203 -2072 271 -2038
rect 361 -2072 429 -2038
rect 519 -2072 587 -2038
rect 677 -2072 745 -2038
rect 835 -2072 903 -2038
rect 993 -2072 1061 -2038
rect 1151 -2072 1219 -2038
rect 1309 -2072 1377 -2038
rect 1467 -2072 1535 -2038
rect 1625 -2072 1693 -2038
rect 1783 -2072 1851 -2038
rect 1941 -2072 2009 -2038
rect 2099 -2072 2167 -2038
rect 2257 -2072 2325 -2038
rect 2415 -2072 2483 -2038
rect 2573 -2072 2641 -2038
rect 2731 -2072 2799 -2038
rect 2889 -2072 2957 -2038
rect 3047 -2072 3115 -2038
rect 3205 -2072 3273 -2038
rect 3363 -2072 3431 -2038
rect 3521 -2072 3589 -2038
rect 3679 -2072 3747 -2038
rect 3837 -2072 3905 -2038
rect 3995 -2072 4063 -2038
rect 4153 -2072 4221 -2038
rect 4311 -2072 4379 -2038
rect 4469 -2072 4537 -2038
rect 4627 -2072 4695 -2038
rect 4785 -2072 4853 -2038
rect 4943 -2072 5011 -2038
rect 5101 -2072 5169 -2038
rect 5259 -2072 5327 -2038
rect 5417 -2072 5485 -2038
rect 5575 -2072 5643 -2038
rect 5733 -2072 5801 -2038
rect 5891 -2072 5959 -2038
rect 6049 -2072 6117 -2038
rect 6207 -2072 6275 -2038
rect 6365 -2072 6433 -2038
rect 6523 -2072 6591 -2038
rect 6681 -2072 6749 -2038
rect 6839 -2072 6907 -2038
rect 6997 -2072 7065 -2038
rect 7155 -2072 7223 -2038
rect 7313 -2072 7381 -2038
rect 7471 -2072 7539 -2038
rect 7629 -2072 7697 -2038
rect 7787 -2072 7855 -2038
rect 7945 -2072 8013 -2038
rect 8103 -2072 8171 -2038
rect 8261 -2072 8329 -2038
rect 8419 -2072 8487 -2038
rect 8577 -2072 8645 -2038
rect 8735 -2072 8803 -2038
rect 8893 -2072 8961 -2038
rect 9051 -2072 9119 -2038
rect 9209 -2072 9277 -2038
rect 9367 -2072 9435 -2038
rect 9525 -2072 9593 -2038
rect 9683 -2072 9751 -2038
rect 9841 -2072 9909 -2038
rect 9999 -2072 10067 -2038
<< metal1 >>
rect -10079 2072 -9987 2078
rect -10079 2038 -10067 2072
rect -9999 2038 -9987 2072
rect -10079 2032 -9987 2038
rect -9921 2072 -9829 2078
rect -9921 2038 -9909 2072
rect -9841 2038 -9829 2072
rect -9921 2032 -9829 2038
rect -9763 2072 -9671 2078
rect -9763 2038 -9751 2072
rect -9683 2038 -9671 2072
rect -9763 2032 -9671 2038
rect -9605 2072 -9513 2078
rect -9605 2038 -9593 2072
rect -9525 2038 -9513 2072
rect -9605 2032 -9513 2038
rect -9447 2072 -9355 2078
rect -9447 2038 -9435 2072
rect -9367 2038 -9355 2072
rect -9447 2032 -9355 2038
rect -9289 2072 -9197 2078
rect -9289 2038 -9277 2072
rect -9209 2038 -9197 2072
rect -9289 2032 -9197 2038
rect -9131 2072 -9039 2078
rect -9131 2038 -9119 2072
rect -9051 2038 -9039 2072
rect -9131 2032 -9039 2038
rect -8973 2072 -8881 2078
rect -8973 2038 -8961 2072
rect -8893 2038 -8881 2072
rect -8973 2032 -8881 2038
rect -8815 2072 -8723 2078
rect -8815 2038 -8803 2072
rect -8735 2038 -8723 2072
rect -8815 2032 -8723 2038
rect -8657 2072 -8565 2078
rect -8657 2038 -8645 2072
rect -8577 2038 -8565 2072
rect -8657 2032 -8565 2038
rect -8499 2072 -8407 2078
rect -8499 2038 -8487 2072
rect -8419 2038 -8407 2072
rect -8499 2032 -8407 2038
rect -8341 2072 -8249 2078
rect -8341 2038 -8329 2072
rect -8261 2038 -8249 2072
rect -8341 2032 -8249 2038
rect -8183 2072 -8091 2078
rect -8183 2038 -8171 2072
rect -8103 2038 -8091 2072
rect -8183 2032 -8091 2038
rect -8025 2072 -7933 2078
rect -8025 2038 -8013 2072
rect -7945 2038 -7933 2072
rect -8025 2032 -7933 2038
rect -7867 2072 -7775 2078
rect -7867 2038 -7855 2072
rect -7787 2038 -7775 2072
rect -7867 2032 -7775 2038
rect -7709 2072 -7617 2078
rect -7709 2038 -7697 2072
rect -7629 2038 -7617 2072
rect -7709 2032 -7617 2038
rect -7551 2072 -7459 2078
rect -7551 2038 -7539 2072
rect -7471 2038 -7459 2072
rect -7551 2032 -7459 2038
rect -7393 2072 -7301 2078
rect -7393 2038 -7381 2072
rect -7313 2038 -7301 2072
rect -7393 2032 -7301 2038
rect -7235 2072 -7143 2078
rect -7235 2038 -7223 2072
rect -7155 2038 -7143 2072
rect -7235 2032 -7143 2038
rect -7077 2072 -6985 2078
rect -7077 2038 -7065 2072
rect -6997 2038 -6985 2072
rect -7077 2032 -6985 2038
rect -6919 2072 -6827 2078
rect -6919 2038 -6907 2072
rect -6839 2038 -6827 2072
rect -6919 2032 -6827 2038
rect -6761 2072 -6669 2078
rect -6761 2038 -6749 2072
rect -6681 2038 -6669 2072
rect -6761 2032 -6669 2038
rect -6603 2072 -6511 2078
rect -6603 2038 -6591 2072
rect -6523 2038 -6511 2072
rect -6603 2032 -6511 2038
rect -6445 2072 -6353 2078
rect -6445 2038 -6433 2072
rect -6365 2038 -6353 2072
rect -6445 2032 -6353 2038
rect -6287 2072 -6195 2078
rect -6287 2038 -6275 2072
rect -6207 2038 -6195 2072
rect -6287 2032 -6195 2038
rect -6129 2072 -6037 2078
rect -6129 2038 -6117 2072
rect -6049 2038 -6037 2072
rect -6129 2032 -6037 2038
rect -5971 2072 -5879 2078
rect -5971 2038 -5959 2072
rect -5891 2038 -5879 2072
rect -5971 2032 -5879 2038
rect -5813 2072 -5721 2078
rect -5813 2038 -5801 2072
rect -5733 2038 -5721 2072
rect -5813 2032 -5721 2038
rect -5655 2072 -5563 2078
rect -5655 2038 -5643 2072
rect -5575 2038 -5563 2072
rect -5655 2032 -5563 2038
rect -5497 2072 -5405 2078
rect -5497 2038 -5485 2072
rect -5417 2038 -5405 2072
rect -5497 2032 -5405 2038
rect -5339 2072 -5247 2078
rect -5339 2038 -5327 2072
rect -5259 2038 -5247 2072
rect -5339 2032 -5247 2038
rect -5181 2072 -5089 2078
rect -5181 2038 -5169 2072
rect -5101 2038 -5089 2072
rect -5181 2032 -5089 2038
rect -5023 2072 -4931 2078
rect -5023 2038 -5011 2072
rect -4943 2038 -4931 2072
rect -5023 2032 -4931 2038
rect -4865 2072 -4773 2078
rect -4865 2038 -4853 2072
rect -4785 2038 -4773 2072
rect -4865 2032 -4773 2038
rect -4707 2072 -4615 2078
rect -4707 2038 -4695 2072
rect -4627 2038 -4615 2072
rect -4707 2032 -4615 2038
rect -4549 2072 -4457 2078
rect -4549 2038 -4537 2072
rect -4469 2038 -4457 2072
rect -4549 2032 -4457 2038
rect -4391 2072 -4299 2078
rect -4391 2038 -4379 2072
rect -4311 2038 -4299 2072
rect -4391 2032 -4299 2038
rect -4233 2072 -4141 2078
rect -4233 2038 -4221 2072
rect -4153 2038 -4141 2072
rect -4233 2032 -4141 2038
rect -4075 2072 -3983 2078
rect -4075 2038 -4063 2072
rect -3995 2038 -3983 2072
rect -4075 2032 -3983 2038
rect -3917 2072 -3825 2078
rect -3917 2038 -3905 2072
rect -3837 2038 -3825 2072
rect -3917 2032 -3825 2038
rect -3759 2072 -3667 2078
rect -3759 2038 -3747 2072
rect -3679 2038 -3667 2072
rect -3759 2032 -3667 2038
rect -3601 2072 -3509 2078
rect -3601 2038 -3589 2072
rect -3521 2038 -3509 2072
rect -3601 2032 -3509 2038
rect -3443 2072 -3351 2078
rect -3443 2038 -3431 2072
rect -3363 2038 -3351 2072
rect -3443 2032 -3351 2038
rect -3285 2072 -3193 2078
rect -3285 2038 -3273 2072
rect -3205 2038 -3193 2072
rect -3285 2032 -3193 2038
rect -3127 2072 -3035 2078
rect -3127 2038 -3115 2072
rect -3047 2038 -3035 2072
rect -3127 2032 -3035 2038
rect -2969 2072 -2877 2078
rect -2969 2038 -2957 2072
rect -2889 2038 -2877 2072
rect -2969 2032 -2877 2038
rect -2811 2072 -2719 2078
rect -2811 2038 -2799 2072
rect -2731 2038 -2719 2072
rect -2811 2032 -2719 2038
rect -2653 2072 -2561 2078
rect -2653 2038 -2641 2072
rect -2573 2038 -2561 2072
rect -2653 2032 -2561 2038
rect -2495 2072 -2403 2078
rect -2495 2038 -2483 2072
rect -2415 2038 -2403 2072
rect -2495 2032 -2403 2038
rect -2337 2072 -2245 2078
rect -2337 2038 -2325 2072
rect -2257 2038 -2245 2072
rect -2337 2032 -2245 2038
rect -2179 2072 -2087 2078
rect -2179 2038 -2167 2072
rect -2099 2038 -2087 2072
rect -2179 2032 -2087 2038
rect -2021 2072 -1929 2078
rect -2021 2038 -2009 2072
rect -1941 2038 -1929 2072
rect -2021 2032 -1929 2038
rect -1863 2072 -1771 2078
rect -1863 2038 -1851 2072
rect -1783 2038 -1771 2072
rect -1863 2032 -1771 2038
rect -1705 2072 -1613 2078
rect -1705 2038 -1693 2072
rect -1625 2038 -1613 2072
rect -1705 2032 -1613 2038
rect -1547 2072 -1455 2078
rect -1547 2038 -1535 2072
rect -1467 2038 -1455 2072
rect -1547 2032 -1455 2038
rect -1389 2072 -1297 2078
rect -1389 2038 -1377 2072
rect -1309 2038 -1297 2072
rect -1389 2032 -1297 2038
rect -1231 2072 -1139 2078
rect -1231 2038 -1219 2072
rect -1151 2038 -1139 2072
rect -1231 2032 -1139 2038
rect -1073 2072 -981 2078
rect -1073 2038 -1061 2072
rect -993 2038 -981 2072
rect -1073 2032 -981 2038
rect -915 2072 -823 2078
rect -915 2038 -903 2072
rect -835 2038 -823 2072
rect -915 2032 -823 2038
rect -757 2072 -665 2078
rect -757 2038 -745 2072
rect -677 2038 -665 2072
rect -757 2032 -665 2038
rect -599 2072 -507 2078
rect -599 2038 -587 2072
rect -519 2038 -507 2072
rect -599 2032 -507 2038
rect -441 2072 -349 2078
rect -441 2038 -429 2072
rect -361 2038 -349 2072
rect -441 2032 -349 2038
rect -283 2072 -191 2078
rect -283 2038 -271 2072
rect -203 2038 -191 2072
rect -283 2032 -191 2038
rect -125 2072 -33 2078
rect -125 2038 -113 2072
rect -45 2038 -33 2072
rect -125 2032 -33 2038
rect 33 2072 125 2078
rect 33 2038 45 2072
rect 113 2038 125 2072
rect 33 2032 125 2038
rect 191 2072 283 2078
rect 191 2038 203 2072
rect 271 2038 283 2072
rect 191 2032 283 2038
rect 349 2072 441 2078
rect 349 2038 361 2072
rect 429 2038 441 2072
rect 349 2032 441 2038
rect 507 2072 599 2078
rect 507 2038 519 2072
rect 587 2038 599 2072
rect 507 2032 599 2038
rect 665 2072 757 2078
rect 665 2038 677 2072
rect 745 2038 757 2072
rect 665 2032 757 2038
rect 823 2072 915 2078
rect 823 2038 835 2072
rect 903 2038 915 2072
rect 823 2032 915 2038
rect 981 2072 1073 2078
rect 981 2038 993 2072
rect 1061 2038 1073 2072
rect 981 2032 1073 2038
rect 1139 2072 1231 2078
rect 1139 2038 1151 2072
rect 1219 2038 1231 2072
rect 1139 2032 1231 2038
rect 1297 2072 1389 2078
rect 1297 2038 1309 2072
rect 1377 2038 1389 2072
rect 1297 2032 1389 2038
rect 1455 2072 1547 2078
rect 1455 2038 1467 2072
rect 1535 2038 1547 2072
rect 1455 2032 1547 2038
rect 1613 2072 1705 2078
rect 1613 2038 1625 2072
rect 1693 2038 1705 2072
rect 1613 2032 1705 2038
rect 1771 2072 1863 2078
rect 1771 2038 1783 2072
rect 1851 2038 1863 2072
rect 1771 2032 1863 2038
rect 1929 2072 2021 2078
rect 1929 2038 1941 2072
rect 2009 2038 2021 2072
rect 1929 2032 2021 2038
rect 2087 2072 2179 2078
rect 2087 2038 2099 2072
rect 2167 2038 2179 2072
rect 2087 2032 2179 2038
rect 2245 2072 2337 2078
rect 2245 2038 2257 2072
rect 2325 2038 2337 2072
rect 2245 2032 2337 2038
rect 2403 2072 2495 2078
rect 2403 2038 2415 2072
rect 2483 2038 2495 2072
rect 2403 2032 2495 2038
rect 2561 2072 2653 2078
rect 2561 2038 2573 2072
rect 2641 2038 2653 2072
rect 2561 2032 2653 2038
rect 2719 2072 2811 2078
rect 2719 2038 2731 2072
rect 2799 2038 2811 2072
rect 2719 2032 2811 2038
rect 2877 2072 2969 2078
rect 2877 2038 2889 2072
rect 2957 2038 2969 2072
rect 2877 2032 2969 2038
rect 3035 2072 3127 2078
rect 3035 2038 3047 2072
rect 3115 2038 3127 2072
rect 3035 2032 3127 2038
rect 3193 2072 3285 2078
rect 3193 2038 3205 2072
rect 3273 2038 3285 2072
rect 3193 2032 3285 2038
rect 3351 2072 3443 2078
rect 3351 2038 3363 2072
rect 3431 2038 3443 2072
rect 3351 2032 3443 2038
rect 3509 2072 3601 2078
rect 3509 2038 3521 2072
rect 3589 2038 3601 2072
rect 3509 2032 3601 2038
rect 3667 2072 3759 2078
rect 3667 2038 3679 2072
rect 3747 2038 3759 2072
rect 3667 2032 3759 2038
rect 3825 2072 3917 2078
rect 3825 2038 3837 2072
rect 3905 2038 3917 2072
rect 3825 2032 3917 2038
rect 3983 2072 4075 2078
rect 3983 2038 3995 2072
rect 4063 2038 4075 2072
rect 3983 2032 4075 2038
rect 4141 2072 4233 2078
rect 4141 2038 4153 2072
rect 4221 2038 4233 2072
rect 4141 2032 4233 2038
rect 4299 2072 4391 2078
rect 4299 2038 4311 2072
rect 4379 2038 4391 2072
rect 4299 2032 4391 2038
rect 4457 2072 4549 2078
rect 4457 2038 4469 2072
rect 4537 2038 4549 2072
rect 4457 2032 4549 2038
rect 4615 2072 4707 2078
rect 4615 2038 4627 2072
rect 4695 2038 4707 2072
rect 4615 2032 4707 2038
rect 4773 2072 4865 2078
rect 4773 2038 4785 2072
rect 4853 2038 4865 2072
rect 4773 2032 4865 2038
rect 4931 2072 5023 2078
rect 4931 2038 4943 2072
rect 5011 2038 5023 2072
rect 4931 2032 5023 2038
rect 5089 2072 5181 2078
rect 5089 2038 5101 2072
rect 5169 2038 5181 2072
rect 5089 2032 5181 2038
rect 5247 2072 5339 2078
rect 5247 2038 5259 2072
rect 5327 2038 5339 2072
rect 5247 2032 5339 2038
rect 5405 2072 5497 2078
rect 5405 2038 5417 2072
rect 5485 2038 5497 2072
rect 5405 2032 5497 2038
rect 5563 2072 5655 2078
rect 5563 2038 5575 2072
rect 5643 2038 5655 2072
rect 5563 2032 5655 2038
rect 5721 2072 5813 2078
rect 5721 2038 5733 2072
rect 5801 2038 5813 2072
rect 5721 2032 5813 2038
rect 5879 2072 5971 2078
rect 5879 2038 5891 2072
rect 5959 2038 5971 2072
rect 5879 2032 5971 2038
rect 6037 2072 6129 2078
rect 6037 2038 6049 2072
rect 6117 2038 6129 2072
rect 6037 2032 6129 2038
rect 6195 2072 6287 2078
rect 6195 2038 6207 2072
rect 6275 2038 6287 2072
rect 6195 2032 6287 2038
rect 6353 2072 6445 2078
rect 6353 2038 6365 2072
rect 6433 2038 6445 2072
rect 6353 2032 6445 2038
rect 6511 2072 6603 2078
rect 6511 2038 6523 2072
rect 6591 2038 6603 2072
rect 6511 2032 6603 2038
rect 6669 2072 6761 2078
rect 6669 2038 6681 2072
rect 6749 2038 6761 2072
rect 6669 2032 6761 2038
rect 6827 2072 6919 2078
rect 6827 2038 6839 2072
rect 6907 2038 6919 2072
rect 6827 2032 6919 2038
rect 6985 2072 7077 2078
rect 6985 2038 6997 2072
rect 7065 2038 7077 2072
rect 6985 2032 7077 2038
rect 7143 2072 7235 2078
rect 7143 2038 7155 2072
rect 7223 2038 7235 2072
rect 7143 2032 7235 2038
rect 7301 2072 7393 2078
rect 7301 2038 7313 2072
rect 7381 2038 7393 2072
rect 7301 2032 7393 2038
rect 7459 2072 7551 2078
rect 7459 2038 7471 2072
rect 7539 2038 7551 2072
rect 7459 2032 7551 2038
rect 7617 2072 7709 2078
rect 7617 2038 7629 2072
rect 7697 2038 7709 2072
rect 7617 2032 7709 2038
rect 7775 2072 7867 2078
rect 7775 2038 7787 2072
rect 7855 2038 7867 2072
rect 7775 2032 7867 2038
rect 7933 2072 8025 2078
rect 7933 2038 7945 2072
rect 8013 2038 8025 2072
rect 7933 2032 8025 2038
rect 8091 2072 8183 2078
rect 8091 2038 8103 2072
rect 8171 2038 8183 2072
rect 8091 2032 8183 2038
rect 8249 2072 8341 2078
rect 8249 2038 8261 2072
rect 8329 2038 8341 2072
rect 8249 2032 8341 2038
rect 8407 2072 8499 2078
rect 8407 2038 8419 2072
rect 8487 2038 8499 2072
rect 8407 2032 8499 2038
rect 8565 2072 8657 2078
rect 8565 2038 8577 2072
rect 8645 2038 8657 2072
rect 8565 2032 8657 2038
rect 8723 2072 8815 2078
rect 8723 2038 8735 2072
rect 8803 2038 8815 2072
rect 8723 2032 8815 2038
rect 8881 2072 8973 2078
rect 8881 2038 8893 2072
rect 8961 2038 8973 2072
rect 8881 2032 8973 2038
rect 9039 2072 9131 2078
rect 9039 2038 9051 2072
rect 9119 2038 9131 2072
rect 9039 2032 9131 2038
rect 9197 2072 9289 2078
rect 9197 2038 9209 2072
rect 9277 2038 9289 2072
rect 9197 2032 9289 2038
rect 9355 2072 9447 2078
rect 9355 2038 9367 2072
rect 9435 2038 9447 2072
rect 9355 2032 9447 2038
rect 9513 2072 9605 2078
rect 9513 2038 9525 2072
rect 9593 2038 9605 2072
rect 9513 2032 9605 2038
rect 9671 2072 9763 2078
rect 9671 2038 9683 2072
rect 9751 2038 9763 2072
rect 9671 2032 9763 2038
rect 9829 2072 9921 2078
rect 9829 2038 9841 2072
rect 9909 2038 9921 2072
rect 9829 2032 9921 2038
rect 9987 2072 10079 2078
rect 9987 2038 9999 2072
rect 10067 2038 10079 2072
rect 9987 2032 10079 2038
rect -10135 1988 -10089 2000
rect -10135 -1988 -10129 1988
rect -10095 -1988 -10089 1988
rect -10135 -2000 -10089 -1988
rect -9977 1988 -9931 2000
rect -9977 -1988 -9971 1988
rect -9937 -1988 -9931 1988
rect -9977 -2000 -9931 -1988
rect -9819 1988 -9773 2000
rect -9819 -1988 -9813 1988
rect -9779 -1988 -9773 1988
rect -9819 -2000 -9773 -1988
rect -9661 1988 -9615 2000
rect -9661 -1988 -9655 1988
rect -9621 -1988 -9615 1988
rect -9661 -2000 -9615 -1988
rect -9503 1988 -9457 2000
rect -9503 -1988 -9497 1988
rect -9463 -1988 -9457 1988
rect -9503 -2000 -9457 -1988
rect -9345 1988 -9299 2000
rect -9345 -1988 -9339 1988
rect -9305 -1988 -9299 1988
rect -9345 -2000 -9299 -1988
rect -9187 1988 -9141 2000
rect -9187 -1988 -9181 1988
rect -9147 -1988 -9141 1988
rect -9187 -2000 -9141 -1988
rect -9029 1988 -8983 2000
rect -9029 -1988 -9023 1988
rect -8989 -1988 -8983 1988
rect -9029 -2000 -8983 -1988
rect -8871 1988 -8825 2000
rect -8871 -1988 -8865 1988
rect -8831 -1988 -8825 1988
rect -8871 -2000 -8825 -1988
rect -8713 1988 -8667 2000
rect -8713 -1988 -8707 1988
rect -8673 -1988 -8667 1988
rect -8713 -2000 -8667 -1988
rect -8555 1988 -8509 2000
rect -8555 -1988 -8549 1988
rect -8515 -1988 -8509 1988
rect -8555 -2000 -8509 -1988
rect -8397 1988 -8351 2000
rect -8397 -1988 -8391 1988
rect -8357 -1988 -8351 1988
rect -8397 -2000 -8351 -1988
rect -8239 1988 -8193 2000
rect -8239 -1988 -8233 1988
rect -8199 -1988 -8193 1988
rect -8239 -2000 -8193 -1988
rect -8081 1988 -8035 2000
rect -8081 -1988 -8075 1988
rect -8041 -1988 -8035 1988
rect -8081 -2000 -8035 -1988
rect -7923 1988 -7877 2000
rect -7923 -1988 -7917 1988
rect -7883 -1988 -7877 1988
rect -7923 -2000 -7877 -1988
rect -7765 1988 -7719 2000
rect -7765 -1988 -7759 1988
rect -7725 -1988 -7719 1988
rect -7765 -2000 -7719 -1988
rect -7607 1988 -7561 2000
rect -7607 -1988 -7601 1988
rect -7567 -1988 -7561 1988
rect -7607 -2000 -7561 -1988
rect -7449 1988 -7403 2000
rect -7449 -1988 -7443 1988
rect -7409 -1988 -7403 1988
rect -7449 -2000 -7403 -1988
rect -7291 1988 -7245 2000
rect -7291 -1988 -7285 1988
rect -7251 -1988 -7245 1988
rect -7291 -2000 -7245 -1988
rect -7133 1988 -7087 2000
rect -7133 -1988 -7127 1988
rect -7093 -1988 -7087 1988
rect -7133 -2000 -7087 -1988
rect -6975 1988 -6929 2000
rect -6975 -1988 -6969 1988
rect -6935 -1988 -6929 1988
rect -6975 -2000 -6929 -1988
rect -6817 1988 -6771 2000
rect -6817 -1988 -6811 1988
rect -6777 -1988 -6771 1988
rect -6817 -2000 -6771 -1988
rect -6659 1988 -6613 2000
rect -6659 -1988 -6653 1988
rect -6619 -1988 -6613 1988
rect -6659 -2000 -6613 -1988
rect -6501 1988 -6455 2000
rect -6501 -1988 -6495 1988
rect -6461 -1988 -6455 1988
rect -6501 -2000 -6455 -1988
rect -6343 1988 -6297 2000
rect -6343 -1988 -6337 1988
rect -6303 -1988 -6297 1988
rect -6343 -2000 -6297 -1988
rect -6185 1988 -6139 2000
rect -6185 -1988 -6179 1988
rect -6145 -1988 -6139 1988
rect -6185 -2000 -6139 -1988
rect -6027 1988 -5981 2000
rect -6027 -1988 -6021 1988
rect -5987 -1988 -5981 1988
rect -6027 -2000 -5981 -1988
rect -5869 1988 -5823 2000
rect -5869 -1988 -5863 1988
rect -5829 -1988 -5823 1988
rect -5869 -2000 -5823 -1988
rect -5711 1988 -5665 2000
rect -5711 -1988 -5705 1988
rect -5671 -1988 -5665 1988
rect -5711 -2000 -5665 -1988
rect -5553 1988 -5507 2000
rect -5553 -1988 -5547 1988
rect -5513 -1988 -5507 1988
rect -5553 -2000 -5507 -1988
rect -5395 1988 -5349 2000
rect -5395 -1988 -5389 1988
rect -5355 -1988 -5349 1988
rect -5395 -2000 -5349 -1988
rect -5237 1988 -5191 2000
rect -5237 -1988 -5231 1988
rect -5197 -1988 -5191 1988
rect -5237 -2000 -5191 -1988
rect -5079 1988 -5033 2000
rect -5079 -1988 -5073 1988
rect -5039 -1988 -5033 1988
rect -5079 -2000 -5033 -1988
rect -4921 1988 -4875 2000
rect -4921 -1988 -4915 1988
rect -4881 -1988 -4875 1988
rect -4921 -2000 -4875 -1988
rect -4763 1988 -4717 2000
rect -4763 -1988 -4757 1988
rect -4723 -1988 -4717 1988
rect -4763 -2000 -4717 -1988
rect -4605 1988 -4559 2000
rect -4605 -1988 -4599 1988
rect -4565 -1988 -4559 1988
rect -4605 -2000 -4559 -1988
rect -4447 1988 -4401 2000
rect -4447 -1988 -4441 1988
rect -4407 -1988 -4401 1988
rect -4447 -2000 -4401 -1988
rect -4289 1988 -4243 2000
rect -4289 -1988 -4283 1988
rect -4249 -1988 -4243 1988
rect -4289 -2000 -4243 -1988
rect -4131 1988 -4085 2000
rect -4131 -1988 -4125 1988
rect -4091 -1988 -4085 1988
rect -4131 -2000 -4085 -1988
rect -3973 1988 -3927 2000
rect -3973 -1988 -3967 1988
rect -3933 -1988 -3927 1988
rect -3973 -2000 -3927 -1988
rect -3815 1988 -3769 2000
rect -3815 -1988 -3809 1988
rect -3775 -1988 -3769 1988
rect -3815 -2000 -3769 -1988
rect -3657 1988 -3611 2000
rect -3657 -1988 -3651 1988
rect -3617 -1988 -3611 1988
rect -3657 -2000 -3611 -1988
rect -3499 1988 -3453 2000
rect -3499 -1988 -3493 1988
rect -3459 -1988 -3453 1988
rect -3499 -2000 -3453 -1988
rect -3341 1988 -3295 2000
rect -3341 -1988 -3335 1988
rect -3301 -1988 -3295 1988
rect -3341 -2000 -3295 -1988
rect -3183 1988 -3137 2000
rect -3183 -1988 -3177 1988
rect -3143 -1988 -3137 1988
rect -3183 -2000 -3137 -1988
rect -3025 1988 -2979 2000
rect -3025 -1988 -3019 1988
rect -2985 -1988 -2979 1988
rect -3025 -2000 -2979 -1988
rect -2867 1988 -2821 2000
rect -2867 -1988 -2861 1988
rect -2827 -1988 -2821 1988
rect -2867 -2000 -2821 -1988
rect -2709 1988 -2663 2000
rect -2709 -1988 -2703 1988
rect -2669 -1988 -2663 1988
rect -2709 -2000 -2663 -1988
rect -2551 1988 -2505 2000
rect -2551 -1988 -2545 1988
rect -2511 -1988 -2505 1988
rect -2551 -2000 -2505 -1988
rect -2393 1988 -2347 2000
rect -2393 -1988 -2387 1988
rect -2353 -1988 -2347 1988
rect -2393 -2000 -2347 -1988
rect -2235 1988 -2189 2000
rect -2235 -1988 -2229 1988
rect -2195 -1988 -2189 1988
rect -2235 -2000 -2189 -1988
rect -2077 1988 -2031 2000
rect -2077 -1988 -2071 1988
rect -2037 -1988 -2031 1988
rect -2077 -2000 -2031 -1988
rect -1919 1988 -1873 2000
rect -1919 -1988 -1913 1988
rect -1879 -1988 -1873 1988
rect -1919 -2000 -1873 -1988
rect -1761 1988 -1715 2000
rect -1761 -1988 -1755 1988
rect -1721 -1988 -1715 1988
rect -1761 -2000 -1715 -1988
rect -1603 1988 -1557 2000
rect -1603 -1988 -1597 1988
rect -1563 -1988 -1557 1988
rect -1603 -2000 -1557 -1988
rect -1445 1988 -1399 2000
rect -1445 -1988 -1439 1988
rect -1405 -1988 -1399 1988
rect -1445 -2000 -1399 -1988
rect -1287 1988 -1241 2000
rect -1287 -1988 -1281 1988
rect -1247 -1988 -1241 1988
rect -1287 -2000 -1241 -1988
rect -1129 1988 -1083 2000
rect -1129 -1988 -1123 1988
rect -1089 -1988 -1083 1988
rect -1129 -2000 -1083 -1988
rect -971 1988 -925 2000
rect -971 -1988 -965 1988
rect -931 -1988 -925 1988
rect -971 -2000 -925 -1988
rect -813 1988 -767 2000
rect -813 -1988 -807 1988
rect -773 -1988 -767 1988
rect -813 -2000 -767 -1988
rect -655 1988 -609 2000
rect -655 -1988 -649 1988
rect -615 -1988 -609 1988
rect -655 -2000 -609 -1988
rect -497 1988 -451 2000
rect -497 -1988 -491 1988
rect -457 -1988 -451 1988
rect -497 -2000 -451 -1988
rect -339 1988 -293 2000
rect -339 -1988 -333 1988
rect -299 -1988 -293 1988
rect -339 -2000 -293 -1988
rect -181 1988 -135 2000
rect -181 -1988 -175 1988
rect -141 -1988 -135 1988
rect -181 -2000 -135 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 135 1988 181 2000
rect 135 -1988 141 1988
rect 175 -1988 181 1988
rect 135 -2000 181 -1988
rect 293 1988 339 2000
rect 293 -1988 299 1988
rect 333 -1988 339 1988
rect 293 -2000 339 -1988
rect 451 1988 497 2000
rect 451 -1988 457 1988
rect 491 -1988 497 1988
rect 451 -2000 497 -1988
rect 609 1988 655 2000
rect 609 -1988 615 1988
rect 649 -1988 655 1988
rect 609 -2000 655 -1988
rect 767 1988 813 2000
rect 767 -1988 773 1988
rect 807 -1988 813 1988
rect 767 -2000 813 -1988
rect 925 1988 971 2000
rect 925 -1988 931 1988
rect 965 -1988 971 1988
rect 925 -2000 971 -1988
rect 1083 1988 1129 2000
rect 1083 -1988 1089 1988
rect 1123 -1988 1129 1988
rect 1083 -2000 1129 -1988
rect 1241 1988 1287 2000
rect 1241 -1988 1247 1988
rect 1281 -1988 1287 1988
rect 1241 -2000 1287 -1988
rect 1399 1988 1445 2000
rect 1399 -1988 1405 1988
rect 1439 -1988 1445 1988
rect 1399 -2000 1445 -1988
rect 1557 1988 1603 2000
rect 1557 -1988 1563 1988
rect 1597 -1988 1603 1988
rect 1557 -2000 1603 -1988
rect 1715 1988 1761 2000
rect 1715 -1988 1721 1988
rect 1755 -1988 1761 1988
rect 1715 -2000 1761 -1988
rect 1873 1988 1919 2000
rect 1873 -1988 1879 1988
rect 1913 -1988 1919 1988
rect 1873 -2000 1919 -1988
rect 2031 1988 2077 2000
rect 2031 -1988 2037 1988
rect 2071 -1988 2077 1988
rect 2031 -2000 2077 -1988
rect 2189 1988 2235 2000
rect 2189 -1988 2195 1988
rect 2229 -1988 2235 1988
rect 2189 -2000 2235 -1988
rect 2347 1988 2393 2000
rect 2347 -1988 2353 1988
rect 2387 -1988 2393 1988
rect 2347 -2000 2393 -1988
rect 2505 1988 2551 2000
rect 2505 -1988 2511 1988
rect 2545 -1988 2551 1988
rect 2505 -2000 2551 -1988
rect 2663 1988 2709 2000
rect 2663 -1988 2669 1988
rect 2703 -1988 2709 1988
rect 2663 -2000 2709 -1988
rect 2821 1988 2867 2000
rect 2821 -1988 2827 1988
rect 2861 -1988 2867 1988
rect 2821 -2000 2867 -1988
rect 2979 1988 3025 2000
rect 2979 -1988 2985 1988
rect 3019 -1988 3025 1988
rect 2979 -2000 3025 -1988
rect 3137 1988 3183 2000
rect 3137 -1988 3143 1988
rect 3177 -1988 3183 1988
rect 3137 -2000 3183 -1988
rect 3295 1988 3341 2000
rect 3295 -1988 3301 1988
rect 3335 -1988 3341 1988
rect 3295 -2000 3341 -1988
rect 3453 1988 3499 2000
rect 3453 -1988 3459 1988
rect 3493 -1988 3499 1988
rect 3453 -2000 3499 -1988
rect 3611 1988 3657 2000
rect 3611 -1988 3617 1988
rect 3651 -1988 3657 1988
rect 3611 -2000 3657 -1988
rect 3769 1988 3815 2000
rect 3769 -1988 3775 1988
rect 3809 -1988 3815 1988
rect 3769 -2000 3815 -1988
rect 3927 1988 3973 2000
rect 3927 -1988 3933 1988
rect 3967 -1988 3973 1988
rect 3927 -2000 3973 -1988
rect 4085 1988 4131 2000
rect 4085 -1988 4091 1988
rect 4125 -1988 4131 1988
rect 4085 -2000 4131 -1988
rect 4243 1988 4289 2000
rect 4243 -1988 4249 1988
rect 4283 -1988 4289 1988
rect 4243 -2000 4289 -1988
rect 4401 1988 4447 2000
rect 4401 -1988 4407 1988
rect 4441 -1988 4447 1988
rect 4401 -2000 4447 -1988
rect 4559 1988 4605 2000
rect 4559 -1988 4565 1988
rect 4599 -1988 4605 1988
rect 4559 -2000 4605 -1988
rect 4717 1988 4763 2000
rect 4717 -1988 4723 1988
rect 4757 -1988 4763 1988
rect 4717 -2000 4763 -1988
rect 4875 1988 4921 2000
rect 4875 -1988 4881 1988
rect 4915 -1988 4921 1988
rect 4875 -2000 4921 -1988
rect 5033 1988 5079 2000
rect 5033 -1988 5039 1988
rect 5073 -1988 5079 1988
rect 5033 -2000 5079 -1988
rect 5191 1988 5237 2000
rect 5191 -1988 5197 1988
rect 5231 -1988 5237 1988
rect 5191 -2000 5237 -1988
rect 5349 1988 5395 2000
rect 5349 -1988 5355 1988
rect 5389 -1988 5395 1988
rect 5349 -2000 5395 -1988
rect 5507 1988 5553 2000
rect 5507 -1988 5513 1988
rect 5547 -1988 5553 1988
rect 5507 -2000 5553 -1988
rect 5665 1988 5711 2000
rect 5665 -1988 5671 1988
rect 5705 -1988 5711 1988
rect 5665 -2000 5711 -1988
rect 5823 1988 5869 2000
rect 5823 -1988 5829 1988
rect 5863 -1988 5869 1988
rect 5823 -2000 5869 -1988
rect 5981 1988 6027 2000
rect 5981 -1988 5987 1988
rect 6021 -1988 6027 1988
rect 5981 -2000 6027 -1988
rect 6139 1988 6185 2000
rect 6139 -1988 6145 1988
rect 6179 -1988 6185 1988
rect 6139 -2000 6185 -1988
rect 6297 1988 6343 2000
rect 6297 -1988 6303 1988
rect 6337 -1988 6343 1988
rect 6297 -2000 6343 -1988
rect 6455 1988 6501 2000
rect 6455 -1988 6461 1988
rect 6495 -1988 6501 1988
rect 6455 -2000 6501 -1988
rect 6613 1988 6659 2000
rect 6613 -1988 6619 1988
rect 6653 -1988 6659 1988
rect 6613 -2000 6659 -1988
rect 6771 1988 6817 2000
rect 6771 -1988 6777 1988
rect 6811 -1988 6817 1988
rect 6771 -2000 6817 -1988
rect 6929 1988 6975 2000
rect 6929 -1988 6935 1988
rect 6969 -1988 6975 1988
rect 6929 -2000 6975 -1988
rect 7087 1988 7133 2000
rect 7087 -1988 7093 1988
rect 7127 -1988 7133 1988
rect 7087 -2000 7133 -1988
rect 7245 1988 7291 2000
rect 7245 -1988 7251 1988
rect 7285 -1988 7291 1988
rect 7245 -2000 7291 -1988
rect 7403 1988 7449 2000
rect 7403 -1988 7409 1988
rect 7443 -1988 7449 1988
rect 7403 -2000 7449 -1988
rect 7561 1988 7607 2000
rect 7561 -1988 7567 1988
rect 7601 -1988 7607 1988
rect 7561 -2000 7607 -1988
rect 7719 1988 7765 2000
rect 7719 -1988 7725 1988
rect 7759 -1988 7765 1988
rect 7719 -2000 7765 -1988
rect 7877 1988 7923 2000
rect 7877 -1988 7883 1988
rect 7917 -1988 7923 1988
rect 7877 -2000 7923 -1988
rect 8035 1988 8081 2000
rect 8035 -1988 8041 1988
rect 8075 -1988 8081 1988
rect 8035 -2000 8081 -1988
rect 8193 1988 8239 2000
rect 8193 -1988 8199 1988
rect 8233 -1988 8239 1988
rect 8193 -2000 8239 -1988
rect 8351 1988 8397 2000
rect 8351 -1988 8357 1988
rect 8391 -1988 8397 1988
rect 8351 -2000 8397 -1988
rect 8509 1988 8555 2000
rect 8509 -1988 8515 1988
rect 8549 -1988 8555 1988
rect 8509 -2000 8555 -1988
rect 8667 1988 8713 2000
rect 8667 -1988 8673 1988
rect 8707 -1988 8713 1988
rect 8667 -2000 8713 -1988
rect 8825 1988 8871 2000
rect 8825 -1988 8831 1988
rect 8865 -1988 8871 1988
rect 8825 -2000 8871 -1988
rect 8983 1988 9029 2000
rect 8983 -1988 8989 1988
rect 9023 -1988 9029 1988
rect 8983 -2000 9029 -1988
rect 9141 1988 9187 2000
rect 9141 -1988 9147 1988
rect 9181 -1988 9187 1988
rect 9141 -2000 9187 -1988
rect 9299 1988 9345 2000
rect 9299 -1988 9305 1988
rect 9339 -1988 9345 1988
rect 9299 -2000 9345 -1988
rect 9457 1988 9503 2000
rect 9457 -1988 9463 1988
rect 9497 -1988 9503 1988
rect 9457 -2000 9503 -1988
rect 9615 1988 9661 2000
rect 9615 -1988 9621 1988
rect 9655 -1988 9661 1988
rect 9615 -2000 9661 -1988
rect 9773 1988 9819 2000
rect 9773 -1988 9779 1988
rect 9813 -1988 9819 1988
rect 9773 -2000 9819 -1988
rect 9931 1988 9977 2000
rect 9931 -1988 9937 1988
rect 9971 -1988 9977 1988
rect 9931 -2000 9977 -1988
rect 10089 1988 10135 2000
rect 10089 -1988 10095 1988
rect 10129 -1988 10135 1988
rect 10089 -2000 10135 -1988
rect -10079 -2038 -9987 -2032
rect -10079 -2072 -10067 -2038
rect -9999 -2072 -9987 -2038
rect -10079 -2078 -9987 -2072
rect -9921 -2038 -9829 -2032
rect -9921 -2072 -9909 -2038
rect -9841 -2072 -9829 -2038
rect -9921 -2078 -9829 -2072
rect -9763 -2038 -9671 -2032
rect -9763 -2072 -9751 -2038
rect -9683 -2072 -9671 -2038
rect -9763 -2078 -9671 -2072
rect -9605 -2038 -9513 -2032
rect -9605 -2072 -9593 -2038
rect -9525 -2072 -9513 -2038
rect -9605 -2078 -9513 -2072
rect -9447 -2038 -9355 -2032
rect -9447 -2072 -9435 -2038
rect -9367 -2072 -9355 -2038
rect -9447 -2078 -9355 -2072
rect -9289 -2038 -9197 -2032
rect -9289 -2072 -9277 -2038
rect -9209 -2072 -9197 -2038
rect -9289 -2078 -9197 -2072
rect -9131 -2038 -9039 -2032
rect -9131 -2072 -9119 -2038
rect -9051 -2072 -9039 -2038
rect -9131 -2078 -9039 -2072
rect -8973 -2038 -8881 -2032
rect -8973 -2072 -8961 -2038
rect -8893 -2072 -8881 -2038
rect -8973 -2078 -8881 -2072
rect -8815 -2038 -8723 -2032
rect -8815 -2072 -8803 -2038
rect -8735 -2072 -8723 -2038
rect -8815 -2078 -8723 -2072
rect -8657 -2038 -8565 -2032
rect -8657 -2072 -8645 -2038
rect -8577 -2072 -8565 -2038
rect -8657 -2078 -8565 -2072
rect -8499 -2038 -8407 -2032
rect -8499 -2072 -8487 -2038
rect -8419 -2072 -8407 -2038
rect -8499 -2078 -8407 -2072
rect -8341 -2038 -8249 -2032
rect -8341 -2072 -8329 -2038
rect -8261 -2072 -8249 -2038
rect -8341 -2078 -8249 -2072
rect -8183 -2038 -8091 -2032
rect -8183 -2072 -8171 -2038
rect -8103 -2072 -8091 -2038
rect -8183 -2078 -8091 -2072
rect -8025 -2038 -7933 -2032
rect -8025 -2072 -8013 -2038
rect -7945 -2072 -7933 -2038
rect -8025 -2078 -7933 -2072
rect -7867 -2038 -7775 -2032
rect -7867 -2072 -7855 -2038
rect -7787 -2072 -7775 -2038
rect -7867 -2078 -7775 -2072
rect -7709 -2038 -7617 -2032
rect -7709 -2072 -7697 -2038
rect -7629 -2072 -7617 -2038
rect -7709 -2078 -7617 -2072
rect -7551 -2038 -7459 -2032
rect -7551 -2072 -7539 -2038
rect -7471 -2072 -7459 -2038
rect -7551 -2078 -7459 -2072
rect -7393 -2038 -7301 -2032
rect -7393 -2072 -7381 -2038
rect -7313 -2072 -7301 -2038
rect -7393 -2078 -7301 -2072
rect -7235 -2038 -7143 -2032
rect -7235 -2072 -7223 -2038
rect -7155 -2072 -7143 -2038
rect -7235 -2078 -7143 -2072
rect -7077 -2038 -6985 -2032
rect -7077 -2072 -7065 -2038
rect -6997 -2072 -6985 -2038
rect -7077 -2078 -6985 -2072
rect -6919 -2038 -6827 -2032
rect -6919 -2072 -6907 -2038
rect -6839 -2072 -6827 -2038
rect -6919 -2078 -6827 -2072
rect -6761 -2038 -6669 -2032
rect -6761 -2072 -6749 -2038
rect -6681 -2072 -6669 -2038
rect -6761 -2078 -6669 -2072
rect -6603 -2038 -6511 -2032
rect -6603 -2072 -6591 -2038
rect -6523 -2072 -6511 -2038
rect -6603 -2078 -6511 -2072
rect -6445 -2038 -6353 -2032
rect -6445 -2072 -6433 -2038
rect -6365 -2072 -6353 -2038
rect -6445 -2078 -6353 -2072
rect -6287 -2038 -6195 -2032
rect -6287 -2072 -6275 -2038
rect -6207 -2072 -6195 -2038
rect -6287 -2078 -6195 -2072
rect -6129 -2038 -6037 -2032
rect -6129 -2072 -6117 -2038
rect -6049 -2072 -6037 -2038
rect -6129 -2078 -6037 -2072
rect -5971 -2038 -5879 -2032
rect -5971 -2072 -5959 -2038
rect -5891 -2072 -5879 -2038
rect -5971 -2078 -5879 -2072
rect -5813 -2038 -5721 -2032
rect -5813 -2072 -5801 -2038
rect -5733 -2072 -5721 -2038
rect -5813 -2078 -5721 -2072
rect -5655 -2038 -5563 -2032
rect -5655 -2072 -5643 -2038
rect -5575 -2072 -5563 -2038
rect -5655 -2078 -5563 -2072
rect -5497 -2038 -5405 -2032
rect -5497 -2072 -5485 -2038
rect -5417 -2072 -5405 -2038
rect -5497 -2078 -5405 -2072
rect -5339 -2038 -5247 -2032
rect -5339 -2072 -5327 -2038
rect -5259 -2072 -5247 -2038
rect -5339 -2078 -5247 -2072
rect -5181 -2038 -5089 -2032
rect -5181 -2072 -5169 -2038
rect -5101 -2072 -5089 -2038
rect -5181 -2078 -5089 -2072
rect -5023 -2038 -4931 -2032
rect -5023 -2072 -5011 -2038
rect -4943 -2072 -4931 -2038
rect -5023 -2078 -4931 -2072
rect -4865 -2038 -4773 -2032
rect -4865 -2072 -4853 -2038
rect -4785 -2072 -4773 -2038
rect -4865 -2078 -4773 -2072
rect -4707 -2038 -4615 -2032
rect -4707 -2072 -4695 -2038
rect -4627 -2072 -4615 -2038
rect -4707 -2078 -4615 -2072
rect -4549 -2038 -4457 -2032
rect -4549 -2072 -4537 -2038
rect -4469 -2072 -4457 -2038
rect -4549 -2078 -4457 -2072
rect -4391 -2038 -4299 -2032
rect -4391 -2072 -4379 -2038
rect -4311 -2072 -4299 -2038
rect -4391 -2078 -4299 -2072
rect -4233 -2038 -4141 -2032
rect -4233 -2072 -4221 -2038
rect -4153 -2072 -4141 -2038
rect -4233 -2078 -4141 -2072
rect -4075 -2038 -3983 -2032
rect -4075 -2072 -4063 -2038
rect -3995 -2072 -3983 -2038
rect -4075 -2078 -3983 -2072
rect -3917 -2038 -3825 -2032
rect -3917 -2072 -3905 -2038
rect -3837 -2072 -3825 -2038
rect -3917 -2078 -3825 -2072
rect -3759 -2038 -3667 -2032
rect -3759 -2072 -3747 -2038
rect -3679 -2072 -3667 -2038
rect -3759 -2078 -3667 -2072
rect -3601 -2038 -3509 -2032
rect -3601 -2072 -3589 -2038
rect -3521 -2072 -3509 -2038
rect -3601 -2078 -3509 -2072
rect -3443 -2038 -3351 -2032
rect -3443 -2072 -3431 -2038
rect -3363 -2072 -3351 -2038
rect -3443 -2078 -3351 -2072
rect -3285 -2038 -3193 -2032
rect -3285 -2072 -3273 -2038
rect -3205 -2072 -3193 -2038
rect -3285 -2078 -3193 -2072
rect -3127 -2038 -3035 -2032
rect -3127 -2072 -3115 -2038
rect -3047 -2072 -3035 -2038
rect -3127 -2078 -3035 -2072
rect -2969 -2038 -2877 -2032
rect -2969 -2072 -2957 -2038
rect -2889 -2072 -2877 -2038
rect -2969 -2078 -2877 -2072
rect -2811 -2038 -2719 -2032
rect -2811 -2072 -2799 -2038
rect -2731 -2072 -2719 -2038
rect -2811 -2078 -2719 -2072
rect -2653 -2038 -2561 -2032
rect -2653 -2072 -2641 -2038
rect -2573 -2072 -2561 -2038
rect -2653 -2078 -2561 -2072
rect -2495 -2038 -2403 -2032
rect -2495 -2072 -2483 -2038
rect -2415 -2072 -2403 -2038
rect -2495 -2078 -2403 -2072
rect -2337 -2038 -2245 -2032
rect -2337 -2072 -2325 -2038
rect -2257 -2072 -2245 -2038
rect -2337 -2078 -2245 -2072
rect -2179 -2038 -2087 -2032
rect -2179 -2072 -2167 -2038
rect -2099 -2072 -2087 -2038
rect -2179 -2078 -2087 -2072
rect -2021 -2038 -1929 -2032
rect -2021 -2072 -2009 -2038
rect -1941 -2072 -1929 -2038
rect -2021 -2078 -1929 -2072
rect -1863 -2038 -1771 -2032
rect -1863 -2072 -1851 -2038
rect -1783 -2072 -1771 -2038
rect -1863 -2078 -1771 -2072
rect -1705 -2038 -1613 -2032
rect -1705 -2072 -1693 -2038
rect -1625 -2072 -1613 -2038
rect -1705 -2078 -1613 -2072
rect -1547 -2038 -1455 -2032
rect -1547 -2072 -1535 -2038
rect -1467 -2072 -1455 -2038
rect -1547 -2078 -1455 -2072
rect -1389 -2038 -1297 -2032
rect -1389 -2072 -1377 -2038
rect -1309 -2072 -1297 -2038
rect -1389 -2078 -1297 -2072
rect -1231 -2038 -1139 -2032
rect -1231 -2072 -1219 -2038
rect -1151 -2072 -1139 -2038
rect -1231 -2078 -1139 -2072
rect -1073 -2038 -981 -2032
rect -1073 -2072 -1061 -2038
rect -993 -2072 -981 -2038
rect -1073 -2078 -981 -2072
rect -915 -2038 -823 -2032
rect -915 -2072 -903 -2038
rect -835 -2072 -823 -2038
rect -915 -2078 -823 -2072
rect -757 -2038 -665 -2032
rect -757 -2072 -745 -2038
rect -677 -2072 -665 -2038
rect -757 -2078 -665 -2072
rect -599 -2038 -507 -2032
rect -599 -2072 -587 -2038
rect -519 -2072 -507 -2038
rect -599 -2078 -507 -2072
rect -441 -2038 -349 -2032
rect -441 -2072 -429 -2038
rect -361 -2072 -349 -2038
rect -441 -2078 -349 -2072
rect -283 -2038 -191 -2032
rect -283 -2072 -271 -2038
rect -203 -2072 -191 -2038
rect -283 -2078 -191 -2072
rect -125 -2038 -33 -2032
rect -125 -2072 -113 -2038
rect -45 -2072 -33 -2038
rect -125 -2078 -33 -2072
rect 33 -2038 125 -2032
rect 33 -2072 45 -2038
rect 113 -2072 125 -2038
rect 33 -2078 125 -2072
rect 191 -2038 283 -2032
rect 191 -2072 203 -2038
rect 271 -2072 283 -2038
rect 191 -2078 283 -2072
rect 349 -2038 441 -2032
rect 349 -2072 361 -2038
rect 429 -2072 441 -2038
rect 349 -2078 441 -2072
rect 507 -2038 599 -2032
rect 507 -2072 519 -2038
rect 587 -2072 599 -2038
rect 507 -2078 599 -2072
rect 665 -2038 757 -2032
rect 665 -2072 677 -2038
rect 745 -2072 757 -2038
rect 665 -2078 757 -2072
rect 823 -2038 915 -2032
rect 823 -2072 835 -2038
rect 903 -2072 915 -2038
rect 823 -2078 915 -2072
rect 981 -2038 1073 -2032
rect 981 -2072 993 -2038
rect 1061 -2072 1073 -2038
rect 981 -2078 1073 -2072
rect 1139 -2038 1231 -2032
rect 1139 -2072 1151 -2038
rect 1219 -2072 1231 -2038
rect 1139 -2078 1231 -2072
rect 1297 -2038 1389 -2032
rect 1297 -2072 1309 -2038
rect 1377 -2072 1389 -2038
rect 1297 -2078 1389 -2072
rect 1455 -2038 1547 -2032
rect 1455 -2072 1467 -2038
rect 1535 -2072 1547 -2038
rect 1455 -2078 1547 -2072
rect 1613 -2038 1705 -2032
rect 1613 -2072 1625 -2038
rect 1693 -2072 1705 -2038
rect 1613 -2078 1705 -2072
rect 1771 -2038 1863 -2032
rect 1771 -2072 1783 -2038
rect 1851 -2072 1863 -2038
rect 1771 -2078 1863 -2072
rect 1929 -2038 2021 -2032
rect 1929 -2072 1941 -2038
rect 2009 -2072 2021 -2038
rect 1929 -2078 2021 -2072
rect 2087 -2038 2179 -2032
rect 2087 -2072 2099 -2038
rect 2167 -2072 2179 -2038
rect 2087 -2078 2179 -2072
rect 2245 -2038 2337 -2032
rect 2245 -2072 2257 -2038
rect 2325 -2072 2337 -2038
rect 2245 -2078 2337 -2072
rect 2403 -2038 2495 -2032
rect 2403 -2072 2415 -2038
rect 2483 -2072 2495 -2038
rect 2403 -2078 2495 -2072
rect 2561 -2038 2653 -2032
rect 2561 -2072 2573 -2038
rect 2641 -2072 2653 -2038
rect 2561 -2078 2653 -2072
rect 2719 -2038 2811 -2032
rect 2719 -2072 2731 -2038
rect 2799 -2072 2811 -2038
rect 2719 -2078 2811 -2072
rect 2877 -2038 2969 -2032
rect 2877 -2072 2889 -2038
rect 2957 -2072 2969 -2038
rect 2877 -2078 2969 -2072
rect 3035 -2038 3127 -2032
rect 3035 -2072 3047 -2038
rect 3115 -2072 3127 -2038
rect 3035 -2078 3127 -2072
rect 3193 -2038 3285 -2032
rect 3193 -2072 3205 -2038
rect 3273 -2072 3285 -2038
rect 3193 -2078 3285 -2072
rect 3351 -2038 3443 -2032
rect 3351 -2072 3363 -2038
rect 3431 -2072 3443 -2038
rect 3351 -2078 3443 -2072
rect 3509 -2038 3601 -2032
rect 3509 -2072 3521 -2038
rect 3589 -2072 3601 -2038
rect 3509 -2078 3601 -2072
rect 3667 -2038 3759 -2032
rect 3667 -2072 3679 -2038
rect 3747 -2072 3759 -2038
rect 3667 -2078 3759 -2072
rect 3825 -2038 3917 -2032
rect 3825 -2072 3837 -2038
rect 3905 -2072 3917 -2038
rect 3825 -2078 3917 -2072
rect 3983 -2038 4075 -2032
rect 3983 -2072 3995 -2038
rect 4063 -2072 4075 -2038
rect 3983 -2078 4075 -2072
rect 4141 -2038 4233 -2032
rect 4141 -2072 4153 -2038
rect 4221 -2072 4233 -2038
rect 4141 -2078 4233 -2072
rect 4299 -2038 4391 -2032
rect 4299 -2072 4311 -2038
rect 4379 -2072 4391 -2038
rect 4299 -2078 4391 -2072
rect 4457 -2038 4549 -2032
rect 4457 -2072 4469 -2038
rect 4537 -2072 4549 -2038
rect 4457 -2078 4549 -2072
rect 4615 -2038 4707 -2032
rect 4615 -2072 4627 -2038
rect 4695 -2072 4707 -2038
rect 4615 -2078 4707 -2072
rect 4773 -2038 4865 -2032
rect 4773 -2072 4785 -2038
rect 4853 -2072 4865 -2038
rect 4773 -2078 4865 -2072
rect 4931 -2038 5023 -2032
rect 4931 -2072 4943 -2038
rect 5011 -2072 5023 -2038
rect 4931 -2078 5023 -2072
rect 5089 -2038 5181 -2032
rect 5089 -2072 5101 -2038
rect 5169 -2072 5181 -2038
rect 5089 -2078 5181 -2072
rect 5247 -2038 5339 -2032
rect 5247 -2072 5259 -2038
rect 5327 -2072 5339 -2038
rect 5247 -2078 5339 -2072
rect 5405 -2038 5497 -2032
rect 5405 -2072 5417 -2038
rect 5485 -2072 5497 -2038
rect 5405 -2078 5497 -2072
rect 5563 -2038 5655 -2032
rect 5563 -2072 5575 -2038
rect 5643 -2072 5655 -2038
rect 5563 -2078 5655 -2072
rect 5721 -2038 5813 -2032
rect 5721 -2072 5733 -2038
rect 5801 -2072 5813 -2038
rect 5721 -2078 5813 -2072
rect 5879 -2038 5971 -2032
rect 5879 -2072 5891 -2038
rect 5959 -2072 5971 -2038
rect 5879 -2078 5971 -2072
rect 6037 -2038 6129 -2032
rect 6037 -2072 6049 -2038
rect 6117 -2072 6129 -2038
rect 6037 -2078 6129 -2072
rect 6195 -2038 6287 -2032
rect 6195 -2072 6207 -2038
rect 6275 -2072 6287 -2038
rect 6195 -2078 6287 -2072
rect 6353 -2038 6445 -2032
rect 6353 -2072 6365 -2038
rect 6433 -2072 6445 -2038
rect 6353 -2078 6445 -2072
rect 6511 -2038 6603 -2032
rect 6511 -2072 6523 -2038
rect 6591 -2072 6603 -2038
rect 6511 -2078 6603 -2072
rect 6669 -2038 6761 -2032
rect 6669 -2072 6681 -2038
rect 6749 -2072 6761 -2038
rect 6669 -2078 6761 -2072
rect 6827 -2038 6919 -2032
rect 6827 -2072 6839 -2038
rect 6907 -2072 6919 -2038
rect 6827 -2078 6919 -2072
rect 6985 -2038 7077 -2032
rect 6985 -2072 6997 -2038
rect 7065 -2072 7077 -2038
rect 6985 -2078 7077 -2072
rect 7143 -2038 7235 -2032
rect 7143 -2072 7155 -2038
rect 7223 -2072 7235 -2038
rect 7143 -2078 7235 -2072
rect 7301 -2038 7393 -2032
rect 7301 -2072 7313 -2038
rect 7381 -2072 7393 -2038
rect 7301 -2078 7393 -2072
rect 7459 -2038 7551 -2032
rect 7459 -2072 7471 -2038
rect 7539 -2072 7551 -2038
rect 7459 -2078 7551 -2072
rect 7617 -2038 7709 -2032
rect 7617 -2072 7629 -2038
rect 7697 -2072 7709 -2038
rect 7617 -2078 7709 -2072
rect 7775 -2038 7867 -2032
rect 7775 -2072 7787 -2038
rect 7855 -2072 7867 -2038
rect 7775 -2078 7867 -2072
rect 7933 -2038 8025 -2032
rect 7933 -2072 7945 -2038
rect 8013 -2072 8025 -2038
rect 7933 -2078 8025 -2072
rect 8091 -2038 8183 -2032
rect 8091 -2072 8103 -2038
rect 8171 -2072 8183 -2038
rect 8091 -2078 8183 -2072
rect 8249 -2038 8341 -2032
rect 8249 -2072 8261 -2038
rect 8329 -2072 8341 -2038
rect 8249 -2078 8341 -2072
rect 8407 -2038 8499 -2032
rect 8407 -2072 8419 -2038
rect 8487 -2072 8499 -2038
rect 8407 -2078 8499 -2072
rect 8565 -2038 8657 -2032
rect 8565 -2072 8577 -2038
rect 8645 -2072 8657 -2038
rect 8565 -2078 8657 -2072
rect 8723 -2038 8815 -2032
rect 8723 -2072 8735 -2038
rect 8803 -2072 8815 -2038
rect 8723 -2078 8815 -2072
rect 8881 -2038 8973 -2032
rect 8881 -2072 8893 -2038
rect 8961 -2072 8973 -2038
rect 8881 -2078 8973 -2072
rect 9039 -2038 9131 -2032
rect 9039 -2072 9051 -2038
rect 9119 -2072 9131 -2038
rect 9039 -2078 9131 -2072
rect 9197 -2038 9289 -2032
rect 9197 -2072 9209 -2038
rect 9277 -2072 9289 -2038
rect 9197 -2078 9289 -2072
rect 9355 -2038 9447 -2032
rect 9355 -2072 9367 -2038
rect 9435 -2072 9447 -2038
rect 9355 -2078 9447 -2072
rect 9513 -2038 9605 -2032
rect 9513 -2072 9525 -2038
rect 9593 -2072 9605 -2038
rect 9513 -2078 9605 -2072
rect 9671 -2038 9763 -2032
rect 9671 -2072 9683 -2038
rect 9751 -2072 9763 -2038
rect 9671 -2078 9763 -2072
rect 9829 -2038 9921 -2032
rect 9829 -2072 9841 -2038
rect 9909 -2072 9921 -2038
rect 9829 -2078 9921 -2072
rect 9987 -2038 10079 -2032
rect 9987 -2072 9999 -2038
rect 10067 -2072 10079 -2038
rect 9987 -2078 10079 -2072
<< properties >>
string FIXED_BBOX -10246 -2193 10246 2193
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 20.0 l 0.5 m 1 nf 128 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
