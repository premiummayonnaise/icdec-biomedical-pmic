magic
tech sky130A
magscale 1 2
timestamp 1769135993
<< pwell >>
rect -483 -380 483 380
<< nmos >>
rect -287 -170 -187 170
rect -129 -170 -29 170
rect 29 -170 129 170
rect 187 -170 287 170
<< ndiff >>
rect -345 158 -287 170
rect -345 -158 -333 158
rect -299 -158 -287 158
rect -345 -170 -287 -158
rect -187 158 -129 170
rect -187 -158 -175 158
rect -141 -158 -129 158
rect -187 -170 -129 -158
rect -29 158 29 170
rect -29 -158 -17 158
rect 17 -158 29 158
rect -29 -170 29 -158
rect 129 158 187 170
rect 129 -158 141 158
rect 175 -158 187 158
rect 129 -170 187 -158
rect 287 158 345 170
rect 287 -158 299 158
rect 333 -158 345 158
rect 287 -170 345 -158
<< ndiffc >>
rect -333 -158 -299 158
rect -175 -158 -141 158
rect -17 -158 17 158
rect 141 -158 175 158
rect 299 -158 333 158
<< psubdiff >>
rect -447 310 -351 344
rect 351 310 447 344
rect -447 248 -413 310
rect 413 248 447 310
rect -447 -310 -413 -248
rect 413 -310 447 -248
rect -447 -344 -351 -310
rect 351 -344 447 -310
<< psubdiffcont >>
rect -351 310 351 344
rect -447 -248 -413 248
rect 413 -248 447 248
rect -351 -344 351 -310
<< poly >>
rect -287 242 -187 258
rect -287 208 -271 242
rect -203 208 -187 242
rect -287 170 -187 208
rect -129 242 -29 258
rect -129 208 -113 242
rect -45 208 -29 242
rect -129 170 -29 208
rect 29 242 129 258
rect 29 208 45 242
rect 113 208 129 242
rect 29 170 129 208
rect 187 242 287 258
rect 187 208 203 242
rect 271 208 287 242
rect 187 170 287 208
rect -287 -208 -187 -170
rect -287 -242 -271 -208
rect -203 -242 -187 -208
rect -287 -258 -187 -242
rect -129 -208 -29 -170
rect -129 -242 -113 -208
rect -45 -242 -29 -208
rect -129 -258 -29 -242
rect 29 -208 129 -170
rect 29 -242 45 -208
rect 113 -242 129 -208
rect 29 -258 129 -242
rect 187 -208 287 -170
rect 187 -242 203 -208
rect 271 -242 287 -208
rect 187 -258 287 -242
<< polycont >>
rect -271 208 -203 242
rect -113 208 -45 242
rect 45 208 113 242
rect 203 208 271 242
rect -271 -242 -203 -208
rect -113 -242 -45 -208
rect 45 -242 113 -208
rect 203 -242 271 -208
<< locali >>
rect -447 310 -351 344
rect 351 310 447 344
rect -447 248 -413 310
rect 413 248 447 310
rect -287 208 -271 242
rect -203 208 -187 242
rect -129 208 -113 242
rect -45 208 -29 242
rect 29 208 45 242
rect 113 208 129 242
rect 187 208 203 242
rect 271 208 287 242
rect -333 158 -299 174
rect -333 -174 -299 -158
rect -175 158 -141 174
rect -175 -174 -141 -158
rect -17 158 17 174
rect -17 -174 17 -158
rect 141 158 175 174
rect 141 -174 175 -158
rect 299 158 333 174
rect 299 -174 333 -158
rect -287 -242 -271 -208
rect -203 -242 -187 -208
rect -129 -242 -113 -208
rect -45 -242 -29 -208
rect 29 -242 45 -208
rect 113 -242 129 -208
rect 187 -242 203 -208
rect 271 -242 287 -208
rect -447 -310 -413 -248
rect 413 -310 447 -248
rect -447 -344 -351 -310
rect 351 -344 447 -310
<< viali >>
rect -271 208 -203 242
rect -113 208 -45 242
rect 45 208 113 242
rect 203 208 271 242
rect -333 -158 -299 158
rect -175 -158 -141 158
rect -17 -158 17 158
rect 141 -158 175 158
rect 299 -158 333 158
rect -271 -242 -203 -208
rect -113 -242 -45 -208
rect 45 -242 113 -208
rect 203 -242 271 -208
<< metal1 >>
rect -283 242 -191 248
rect -283 208 -271 242
rect -203 208 -191 242
rect -283 202 -191 208
rect -125 242 -33 248
rect -125 208 -113 242
rect -45 208 -33 242
rect -125 202 -33 208
rect 33 242 125 248
rect 33 208 45 242
rect 113 208 125 242
rect 33 202 125 208
rect 191 242 283 248
rect 191 208 203 242
rect 271 208 283 242
rect 191 202 283 208
rect -339 158 -293 170
rect -339 -158 -333 158
rect -299 -158 -293 158
rect -339 -170 -293 -158
rect -181 158 -135 170
rect -181 -158 -175 158
rect -141 -158 -135 158
rect -181 -170 -135 -158
rect -23 158 23 170
rect -23 -158 -17 158
rect 17 -158 23 158
rect -23 -170 23 -158
rect 135 158 181 170
rect 135 -158 141 158
rect 175 -158 181 158
rect 135 -170 181 -158
rect 293 158 339 170
rect 293 -158 299 158
rect 333 -158 339 158
rect 293 -170 339 -158
rect -283 -208 -191 -202
rect -283 -242 -271 -208
rect -203 -242 -191 -208
rect -283 -248 -191 -242
rect -125 -208 -33 -202
rect -125 -242 -113 -208
rect -45 -242 -33 -208
rect -125 -248 -33 -242
rect 33 -208 125 -202
rect 33 -242 45 -208
rect 113 -242 125 -208
rect 33 -248 125 -242
rect 191 -208 283 -202
rect 191 -242 203 -208
rect 271 -242 283 -208
rect 191 -248 283 -242
<< properties >>
string FIXED_BBOX -430 -327 430 327
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.7 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
