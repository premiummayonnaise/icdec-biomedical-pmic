magic
tech sky130A
magscale 1 2
timestamp 1769400417
<< nwell >>
rect -4993 -408 4993 442
<< pmos >>
rect -4899 -308 -4649 380
rect -4591 -308 -4341 380
rect -4283 -308 -4033 380
rect -3975 -308 -3725 380
rect -3667 -308 -3417 380
rect -3359 -308 -3109 380
rect -3051 -308 -2801 380
rect -2743 -308 -2493 380
rect -2435 -308 -2185 380
rect -2127 -308 -1877 380
rect -1819 -308 -1569 380
rect -1511 -308 -1261 380
rect -1203 -308 -953 380
rect -895 -308 -645 380
rect -587 -308 -337 380
rect -279 -308 -29 380
rect 29 -308 279 380
rect 337 -308 587 380
rect 645 -308 895 380
rect 953 -308 1203 380
rect 1261 -308 1511 380
rect 1569 -308 1819 380
rect 1877 -308 2127 380
rect 2185 -308 2435 380
rect 2493 -308 2743 380
rect 2801 -308 3051 380
rect 3109 -308 3359 380
rect 3417 -308 3667 380
rect 3725 -308 3975 380
rect 4033 -308 4283 380
rect 4341 -308 4591 380
rect 4649 -308 4899 380
<< pdiff >>
rect -4957 368 -4899 380
rect -4957 -296 -4945 368
rect -4911 -296 -4899 368
rect -4957 -308 -4899 -296
rect -4649 368 -4591 380
rect -4649 -296 -4637 368
rect -4603 -296 -4591 368
rect -4649 -308 -4591 -296
rect -4341 368 -4283 380
rect -4341 -296 -4329 368
rect -4295 -296 -4283 368
rect -4341 -308 -4283 -296
rect -4033 368 -3975 380
rect -4033 -296 -4021 368
rect -3987 -296 -3975 368
rect -4033 -308 -3975 -296
rect -3725 368 -3667 380
rect -3725 -296 -3713 368
rect -3679 -296 -3667 368
rect -3725 -308 -3667 -296
rect -3417 368 -3359 380
rect -3417 -296 -3405 368
rect -3371 -296 -3359 368
rect -3417 -308 -3359 -296
rect -3109 368 -3051 380
rect -3109 -296 -3097 368
rect -3063 -296 -3051 368
rect -3109 -308 -3051 -296
rect -2801 368 -2743 380
rect -2801 -296 -2789 368
rect -2755 -296 -2743 368
rect -2801 -308 -2743 -296
rect -2493 368 -2435 380
rect -2493 -296 -2481 368
rect -2447 -296 -2435 368
rect -2493 -308 -2435 -296
rect -2185 368 -2127 380
rect -2185 -296 -2173 368
rect -2139 -296 -2127 368
rect -2185 -308 -2127 -296
rect -1877 368 -1819 380
rect -1877 -296 -1865 368
rect -1831 -296 -1819 368
rect -1877 -308 -1819 -296
rect -1569 368 -1511 380
rect -1569 -296 -1557 368
rect -1523 -296 -1511 368
rect -1569 -308 -1511 -296
rect -1261 368 -1203 380
rect -1261 -296 -1249 368
rect -1215 -296 -1203 368
rect -1261 -308 -1203 -296
rect -953 368 -895 380
rect -953 -296 -941 368
rect -907 -296 -895 368
rect -953 -308 -895 -296
rect -645 368 -587 380
rect -645 -296 -633 368
rect -599 -296 -587 368
rect -645 -308 -587 -296
rect -337 368 -279 380
rect -337 -296 -325 368
rect -291 -296 -279 368
rect -337 -308 -279 -296
rect -29 368 29 380
rect -29 -296 -17 368
rect 17 -296 29 368
rect -29 -308 29 -296
rect 279 368 337 380
rect 279 -296 291 368
rect 325 -296 337 368
rect 279 -308 337 -296
rect 587 368 645 380
rect 587 -296 599 368
rect 633 -296 645 368
rect 587 -308 645 -296
rect 895 368 953 380
rect 895 -296 907 368
rect 941 -296 953 368
rect 895 -308 953 -296
rect 1203 368 1261 380
rect 1203 -296 1215 368
rect 1249 -296 1261 368
rect 1203 -308 1261 -296
rect 1511 368 1569 380
rect 1511 -296 1523 368
rect 1557 -296 1569 368
rect 1511 -308 1569 -296
rect 1819 368 1877 380
rect 1819 -296 1831 368
rect 1865 -296 1877 368
rect 1819 -308 1877 -296
rect 2127 368 2185 380
rect 2127 -296 2139 368
rect 2173 -296 2185 368
rect 2127 -308 2185 -296
rect 2435 368 2493 380
rect 2435 -296 2447 368
rect 2481 -296 2493 368
rect 2435 -308 2493 -296
rect 2743 368 2801 380
rect 2743 -296 2755 368
rect 2789 -296 2801 368
rect 2743 -308 2801 -296
rect 3051 368 3109 380
rect 3051 -296 3063 368
rect 3097 -296 3109 368
rect 3051 -308 3109 -296
rect 3359 368 3417 380
rect 3359 -296 3371 368
rect 3405 -296 3417 368
rect 3359 -308 3417 -296
rect 3667 368 3725 380
rect 3667 -296 3679 368
rect 3713 -296 3725 368
rect 3667 -308 3725 -296
rect 3975 368 4033 380
rect 3975 -296 3987 368
rect 4021 -296 4033 368
rect 3975 -308 4033 -296
rect 4283 368 4341 380
rect 4283 -296 4295 368
rect 4329 -296 4341 368
rect 4283 -308 4341 -296
rect 4591 368 4649 380
rect 4591 -296 4603 368
rect 4637 -296 4649 368
rect 4591 -308 4649 -296
rect 4899 368 4957 380
rect 4899 -296 4911 368
rect 4945 -296 4957 368
rect 4899 -308 4957 -296
<< pdiffc >>
rect -4945 -296 -4911 368
rect -4637 -296 -4603 368
rect -4329 -296 -4295 368
rect -4021 -296 -3987 368
rect -3713 -296 -3679 368
rect -3405 -296 -3371 368
rect -3097 -296 -3063 368
rect -2789 -296 -2755 368
rect -2481 -296 -2447 368
rect -2173 -296 -2139 368
rect -1865 -296 -1831 368
rect -1557 -296 -1523 368
rect -1249 -296 -1215 368
rect -941 -296 -907 368
rect -633 -296 -599 368
rect -325 -296 -291 368
rect -17 -296 17 368
rect 291 -296 325 368
rect 599 -296 633 368
rect 907 -296 941 368
rect 1215 -296 1249 368
rect 1523 -296 1557 368
rect 1831 -296 1865 368
rect 2139 -296 2173 368
rect 2447 -296 2481 368
rect 2755 -296 2789 368
rect 3063 -296 3097 368
rect 3371 -296 3405 368
rect 3679 -296 3713 368
rect 3987 -296 4021 368
rect 4295 -296 4329 368
rect 4603 -296 4637 368
rect 4911 -296 4945 368
<< poly >>
rect -4899 380 -4649 406
rect -4591 380 -4341 406
rect -4283 380 -4033 406
rect -3975 380 -3725 406
rect -3667 380 -3417 406
rect -3359 380 -3109 406
rect -3051 380 -2801 406
rect -2743 380 -2493 406
rect -2435 380 -2185 406
rect -2127 380 -1877 406
rect -1819 380 -1569 406
rect -1511 380 -1261 406
rect -1203 380 -953 406
rect -895 380 -645 406
rect -587 380 -337 406
rect -279 380 -29 406
rect 29 380 279 406
rect 337 380 587 406
rect 645 380 895 406
rect 953 380 1203 406
rect 1261 380 1511 406
rect 1569 380 1819 406
rect 1877 380 2127 406
rect 2185 380 2435 406
rect 2493 380 2743 406
rect 2801 380 3051 406
rect 3109 380 3359 406
rect 3417 380 3667 406
rect 3725 380 3975 406
rect 4033 380 4283 406
rect 4341 380 4591 406
rect 4649 380 4899 406
rect -4899 -355 -4649 -308
rect -4899 -389 -4883 -355
rect -4665 -389 -4649 -355
rect -4899 -405 -4649 -389
rect -4591 -355 -4341 -308
rect -4591 -389 -4575 -355
rect -4357 -389 -4341 -355
rect -4591 -405 -4341 -389
rect -4283 -355 -4033 -308
rect -4283 -389 -4267 -355
rect -4049 -389 -4033 -355
rect -4283 -405 -4033 -389
rect -3975 -355 -3725 -308
rect -3975 -389 -3959 -355
rect -3741 -389 -3725 -355
rect -3975 -405 -3725 -389
rect -3667 -355 -3417 -308
rect -3667 -389 -3651 -355
rect -3433 -389 -3417 -355
rect -3667 -405 -3417 -389
rect -3359 -355 -3109 -308
rect -3359 -389 -3343 -355
rect -3125 -389 -3109 -355
rect -3359 -405 -3109 -389
rect -3051 -355 -2801 -308
rect -3051 -389 -3035 -355
rect -2817 -389 -2801 -355
rect -3051 -405 -2801 -389
rect -2743 -355 -2493 -308
rect -2743 -389 -2727 -355
rect -2509 -389 -2493 -355
rect -2743 -405 -2493 -389
rect -2435 -355 -2185 -308
rect -2435 -389 -2419 -355
rect -2201 -389 -2185 -355
rect -2435 -405 -2185 -389
rect -2127 -355 -1877 -308
rect -2127 -389 -2111 -355
rect -1893 -389 -1877 -355
rect -2127 -405 -1877 -389
rect -1819 -355 -1569 -308
rect -1819 -389 -1803 -355
rect -1585 -389 -1569 -355
rect -1819 -405 -1569 -389
rect -1511 -355 -1261 -308
rect -1511 -389 -1495 -355
rect -1277 -389 -1261 -355
rect -1511 -405 -1261 -389
rect -1203 -355 -953 -308
rect -1203 -389 -1187 -355
rect -969 -389 -953 -355
rect -1203 -405 -953 -389
rect -895 -355 -645 -308
rect -895 -389 -879 -355
rect -661 -389 -645 -355
rect -895 -405 -645 -389
rect -587 -355 -337 -308
rect -587 -389 -571 -355
rect -353 -389 -337 -355
rect -587 -405 -337 -389
rect -279 -355 -29 -308
rect -279 -389 -263 -355
rect -45 -389 -29 -355
rect -279 -405 -29 -389
rect 29 -355 279 -308
rect 29 -389 45 -355
rect 263 -389 279 -355
rect 29 -405 279 -389
rect 337 -355 587 -308
rect 337 -389 353 -355
rect 571 -389 587 -355
rect 337 -405 587 -389
rect 645 -355 895 -308
rect 645 -389 661 -355
rect 879 -389 895 -355
rect 645 -405 895 -389
rect 953 -355 1203 -308
rect 953 -389 969 -355
rect 1187 -389 1203 -355
rect 953 -405 1203 -389
rect 1261 -355 1511 -308
rect 1261 -389 1277 -355
rect 1495 -389 1511 -355
rect 1261 -405 1511 -389
rect 1569 -355 1819 -308
rect 1569 -389 1585 -355
rect 1803 -389 1819 -355
rect 1569 -405 1819 -389
rect 1877 -355 2127 -308
rect 1877 -389 1893 -355
rect 2111 -389 2127 -355
rect 1877 -405 2127 -389
rect 2185 -355 2435 -308
rect 2185 -389 2201 -355
rect 2419 -389 2435 -355
rect 2185 -405 2435 -389
rect 2493 -355 2743 -308
rect 2493 -389 2509 -355
rect 2727 -389 2743 -355
rect 2493 -405 2743 -389
rect 2801 -355 3051 -308
rect 2801 -389 2817 -355
rect 3035 -389 3051 -355
rect 2801 -405 3051 -389
rect 3109 -355 3359 -308
rect 3109 -389 3125 -355
rect 3343 -389 3359 -355
rect 3109 -405 3359 -389
rect 3417 -355 3667 -308
rect 3417 -389 3433 -355
rect 3651 -389 3667 -355
rect 3417 -405 3667 -389
rect 3725 -355 3975 -308
rect 3725 -389 3741 -355
rect 3959 -389 3975 -355
rect 3725 -405 3975 -389
rect 4033 -355 4283 -308
rect 4033 -389 4049 -355
rect 4267 -389 4283 -355
rect 4033 -405 4283 -389
rect 4341 -355 4591 -308
rect 4341 -389 4357 -355
rect 4575 -389 4591 -355
rect 4341 -405 4591 -389
rect 4649 -355 4899 -308
rect 4649 -389 4665 -355
rect 4883 -389 4899 -355
rect 4649 -405 4899 -389
<< polycont >>
rect -4883 -389 -4665 -355
rect -4575 -389 -4357 -355
rect -4267 -389 -4049 -355
rect -3959 -389 -3741 -355
rect -3651 -389 -3433 -355
rect -3343 -389 -3125 -355
rect -3035 -389 -2817 -355
rect -2727 -389 -2509 -355
rect -2419 -389 -2201 -355
rect -2111 -389 -1893 -355
rect -1803 -389 -1585 -355
rect -1495 -389 -1277 -355
rect -1187 -389 -969 -355
rect -879 -389 -661 -355
rect -571 -389 -353 -355
rect -263 -389 -45 -355
rect 45 -389 263 -355
rect 353 -389 571 -355
rect 661 -389 879 -355
rect 969 -389 1187 -355
rect 1277 -389 1495 -355
rect 1585 -389 1803 -355
rect 1893 -389 2111 -355
rect 2201 -389 2419 -355
rect 2509 -389 2727 -355
rect 2817 -389 3035 -355
rect 3125 -389 3343 -355
rect 3433 -389 3651 -355
rect 3741 -389 3959 -355
rect 4049 -389 4267 -355
rect 4357 -389 4575 -355
rect 4665 -389 4883 -355
<< locali >>
rect -4945 368 -4911 384
rect -4945 -312 -4911 -296
rect -4637 368 -4603 384
rect -4637 -312 -4603 -296
rect -4329 368 -4295 384
rect -4329 -312 -4295 -296
rect -4021 368 -3987 384
rect -4021 -312 -3987 -296
rect -3713 368 -3679 384
rect -3713 -312 -3679 -296
rect -3405 368 -3371 384
rect -3405 -312 -3371 -296
rect -3097 368 -3063 384
rect -3097 -312 -3063 -296
rect -2789 368 -2755 384
rect -2789 -312 -2755 -296
rect -2481 368 -2447 384
rect -2481 -312 -2447 -296
rect -2173 368 -2139 384
rect -2173 -312 -2139 -296
rect -1865 368 -1831 384
rect -1865 -312 -1831 -296
rect -1557 368 -1523 384
rect -1557 -312 -1523 -296
rect -1249 368 -1215 384
rect -1249 -312 -1215 -296
rect -941 368 -907 384
rect -941 -312 -907 -296
rect -633 368 -599 384
rect -633 -312 -599 -296
rect -325 368 -291 384
rect -325 -312 -291 -296
rect -17 368 17 384
rect -17 -312 17 -296
rect 291 368 325 384
rect 291 -312 325 -296
rect 599 368 633 384
rect 599 -312 633 -296
rect 907 368 941 384
rect 907 -312 941 -296
rect 1215 368 1249 384
rect 1215 -312 1249 -296
rect 1523 368 1557 384
rect 1523 -312 1557 -296
rect 1831 368 1865 384
rect 1831 -312 1865 -296
rect 2139 368 2173 384
rect 2139 -312 2173 -296
rect 2447 368 2481 384
rect 2447 -312 2481 -296
rect 2755 368 2789 384
rect 2755 -312 2789 -296
rect 3063 368 3097 384
rect 3063 -312 3097 -296
rect 3371 368 3405 384
rect 3371 -312 3405 -296
rect 3679 368 3713 384
rect 3679 -312 3713 -296
rect 3987 368 4021 384
rect 3987 -312 4021 -296
rect 4295 368 4329 384
rect 4295 -312 4329 -296
rect 4603 368 4637 384
rect 4603 -312 4637 -296
rect 4911 368 4945 384
rect 4911 -312 4945 -296
rect -4899 -389 -4883 -355
rect -4665 -389 -4649 -355
rect -4591 -389 -4575 -355
rect -4357 -389 -4341 -355
rect -4283 -389 -4267 -355
rect -4049 -389 -4033 -355
rect -3975 -389 -3959 -355
rect -3741 -389 -3725 -355
rect -3667 -389 -3651 -355
rect -3433 -389 -3417 -355
rect -3359 -389 -3343 -355
rect -3125 -389 -3109 -355
rect -3051 -389 -3035 -355
rect -2817 -389 -2801 -355
rect -2743 -389 -2727 -355
rect -2509 -389 -2493 -355
rect -2435 -389 -2419 -355
rect -2201 -389 -2185 -355
rect -2127 -389 -2111 -355
rect -1893 -389 -1877 -355
rect -1819 -389 -1803 -355
rect -1585 -389 -1569 -355
rect -1511 -389 -1495 -355
rect -1277 -389 -1261 -355
rect -1203 -389 -1187 -355
rect -969 -389 -953 -355
rect -895 -389 -879 -355
rect -661 -389 -645 -355
rect -587 -389 -571 -355
rect -353 -389 -337 -355
rect -279 -389 -263 -355
rect -45 -389 -29 -355
rect 29 -389 45 -355
rect 263 -389 279 -355
rect 337 -389 353 -355
rect 571 -389 587 -355
rect 645 -389 661 -355
rect 879 -389 895 -355
rect 953 -389 969 -355
rect 1187 -389 1203 -355
rect 1261 -389 1277 -355
rect 1495 -389 1511 -355
rect 1569 -389 1585 -355
rect 1803 -389 1819 -355
rect 1877 -389 1893 -355
rect 2111 -389 2127 -355
rect 2185 -389 2201 -355
rect 2419 -389 2435 -355
rect 2493 -389 2509 -355
rect 2727 -389 2743 -355
rect 2801 -389 2817 -355
rect 3035 -389 3051 -355
rect 3109 -389 3125 -355
rect 3343 -389 3359 -355
rect 3417 -389 3433 -355
rect 3651 -389 3667 -355
rect 3725 -389 3741 -355
rect 3959 -389 3975 -355
rect 4033 -389 4049 -355
rect 4267 -389 4283 -355
rect 4341 -389 4357 -355
rect 4575 -389 4591 -355
rect 4649 -389 4665 -355
rect 4883 -389 4899 -355
<< viali >>
rect -4945 -296 -4911 368
rect -4637 -296 -4603 368
rect -4329 -296 -4295 368
rect -4021 -296 -3987 368
rect -3713 -296 -3679 368
rect -3405 -296 -3371 368
rect -3097 -296 -3063 368
rect -2789 -296 -2755 368
rect -2481 -296 -2447 368
rect -2173 -296 -2139 368
rect -1865 -296 -1831 368
rect -1557 -296 -1523 368
rect -1249 -296 -1215 368
rect -941 -296 -907 368
rect -633 -296 -599 368
rect -325 -296 -291 368
rect -17 -296 17 368
rect 291 -296 325 368
rect 599 -296 633 368
rect 907 -296 941 368
rect 1215 -296 1249 368
rect 1523 -296 1557 368
rect 1831 -296 1865 368
rect 2139 -296 2173 368
rect 2447 -296 2481 368
rect 2755 -296 2789 368
rect 3063 -296 3097 368
rect 3371 -296 3405 368
rect 3679 -296 3713 368
rect 3987 -296 4021 368
rect 4295 -296 4329 368
rect 4603 -296 4637 368
rect 4911 -296 4945 368
rect -4883 -389 -4665 -355
rect -4575 -389 -4357 -355
rect -4267 -389 -4049 -355
rect -3959 -389 -3741 -355
rect -3651 -389 -3433 -355
rect -3343 -389 -3125 -355
rect -3035 -389 -2817 -355
rect -2727 -389 -2509 -355
rect -2419 -389 -2201 -355
rect -2111 -389 -1893 -355
rect -1803 -389 -1585 -355
rect -1495 -389 -1277 -355
rect -1187 -389 -969 -355
rect -879 -389 -661 -355
rect -571 -389 -353 -355
rect -263 -389 -45 -355
rect 45 -389 263 -355
rect 353 -389 571 -355
rect 661 -389 879 -355
rect 969 -389 1187 -355
rect 1277 -389 1495 -355
rect 1585 -389 1803 -355
rect 1893 -389 2111 -355
rect 2201 -389 2419 -355
rect 2509 -389 2727 -355
rect 2817 -389 3035 -355
rect 3125 -389 3343 -355
rect 3433 -389 3651 -355
rect 3741 -389 3959 -355
rect 4049 -389 4267 -355
rect 4357 -389 4575 -355
rect 4665 -389 4883 -355
<< metal1 >>
rect -4951 368 -4905 380
rect -4951 -296 -4945 368
rect -4911 -296 -4905 368
rect -4951 -308 -4905 -296
rect -4643 368 -4597 380
rect -4643 -296 -4637 368
rect -4603 -296 -4597 368
rect -4643 -308 -4597 -296
rect -4335 368 -4289 380
rect -4335 -296 -4329 368
rect -4295 -296 -4289 368
rect -4335 -308 -4289 -296
rect -4027 368 -3981 380
rect -4027 -296 -4021 368
rect -3987 -296 -3981 368
rect -4027 -308 -3981 -296
rect -3719 368 -3673 380
rect -3719 -296 -3713 368
rect -3679 -296 -3673 368
rect -3719 -308 -3673 -296
rect -3411 368 -3365 380
rect -3411 -296 -3405 368
rect -3371 -296 -3365 368
rect -3411 -308 -3365 -296
rect -3103 368 -3057 380
rect -3103 -296 -3097 368
rect -3063 -296 -3057 368
rect -3103 -308 -3057 -296
rect -2795 368 -2749 380
rect -2795 -296 -2789 368
rect -2755 -296 -2749 368
rect -2795 -308 -2749 -296
rect -2487 368 -2441 380
rect -2487 -296 -2481 368
rect -2447 -296 -2441 368
rect -2487 -308 -2441 -296
rect -2179 368 -2133 380
rect -2179 -296 -2173 368
rect -2139 -296 -2133 368
rect -2179 -308 -2133 -296
rect -1871 368 -1825 380
rect -1871 -296 -1865 368
rect -1831 -296 -1825 368
rect -1871 -308 -1825 -296
rect -1563 368 -1517 380
rect -1563 -296 -1557 368
rect -1523 -296 -1517 368
rect -1563 -308 -1517 -296
rect -1255 368 -1209 380
rect -1255 -296 -1249 368
rect -1215 -296 -1209 368
rect -1255 -308 -1209 -296
rect -947 368 -901 380
rect -947 -296 -941 368
rect -907 -296 -901 368
rect -947 -308 -901 -296
rect -639 368 -593 380
rect -639 -296 -633 368
rect -599 -296 -593 368
rect -639 -308 -593 -296
rect -331 368 -285 380
rect -331 -296 -325 368
rect -291 -296 -285 368
rect -331 -308 -285 -296
rect -23 368 23 380
rect -23 -296 -17 368
rect 17 -296 23 368
rect -23 -308 23 -296
rect 285 368 331 380
rect 285 -296 291 368
rect 325 -296 331 368
rect 285 -308 331 -296
rect 593 368 639 380
rect 593 -296 599 368
rect 633 -296 639 368
rect 593 -308 639 -296
rect 901 368 947 380
rect 901 -296 907 368
rect 941 -296 947 368
rect 901 -308 947 -296
rect 1209 368 1255 380
rect 1209 -296 1215 368
rect 1249 -296 1255 368
rect 1209 -308 1255 -296
rect 1517 368 1563 380
rect 1517 -296 1523 368
rect 1557 -296 1563 368
rect 1517 -308 1563 -296
rect 1825 368 1871 380
rect 1825 -296 1831 368
rect 1865 -296 1871 368
rect 1825 -308 1871 -296
rect 2133 368 2179 380
rect 2133 -296 2139 368
rect 2173 -296 2179 368
rect 2133 -308 2179 -296
rect 2441 368 2487 380
rect 2441 -296 2447 368
rect 2481 -296 2487 368
rect 2441 -308 2487 -296
rect 2749 368 2795 380
rect 2749 -296 2755 368
rect 2789 -296 2795 368
rect 2749 -308 2795 -296
rect 3057 368 3103 380
rect 3057 -296 3063 368
rect 3097 -296 3103 368
rect 3057 -308 3103 -296
rect 3365 368 3411 380
rect 3365 -296 3371 368
rect 3405 -296 3411 368
rect 3365 -308 3411 -296
rect 3673 368 3719 380
rect 3673 -296 3679 368
rect 3713 -296 3719 368
rect 3673 -308 3719 -296
rect 3981 368 4027 380
rect 3981 -296 3987 368
rect 4021 -296 4027 368
rect 3981 -308 4027 -296
rect 4289 368 4335 380
rect 4289 -296 4295 368
rect 4329 -296 4335 368
rect 4289 -308 4335 -296
rect 4597 368 4643 380
rect 4597 -296 4603 368
rect 4637 -296 4643 368
rect 4597 -308 4643 -296
rect 4905 368 4951 380
rect 4905 -296 4911 368
rect 4945 -296 4951 368
rect 4905 -308 4951 -296
rect -4895 -355 -4653 -349
rect -4895 -389 -4883 -355
rect -4665 -389 -4653 -355
rect -4895 -395 -4653 -389
rect -4587 -355 -4345 -349
rect -4587 -389 -4575 -355
rect -4357 -389 -4345 -355
rect -4587 -395 -4345 -389
rect -4279 -355 -4037 -349
rect -4279 -389 -4267 -355
rect -4049 -389 -4037 -355
rect -4279 -395 -4037 -389
rect -3971 -355 -3729 -349
rect -3971 -389 -3959 -355
rect -3741 -389 -3729 -355
rect -3971 -395 -3729 -389
rect -3663 -355 -3421 -349
rect -3663 -389 -3651 -355
rect -3433 -389 -3421 -355
rect -3663 -395 -3421 -389
rect -3355 -355 -3113 -349
rect -3355 -389 -3343 -355
rect -3125 -389 -3113 -355
rect -3355 -395 -3113 -389
rect -3047 -355 -2805 -349
rect -3047 -389 -3035 -355
rect -2817 -389 -2805 -355
rect -3047 -395 -2805 -389
rect -2739 -355 -2497 -349
rect -2739 -389 -2727 -355
rect -2509 -389 -2497 -355
rect -2739 -395 -2497 -389
rect -2431 -355 -2189 -349
rect -2431 -389 -2419 -355
rect -2201 -389 -2189 -355
rect -2431 -395 -2189 -389
rect -2123 -355 -1881 -349
rect -2123 -389 -2111 -355
rect -1893 -389 -1881 -355
rect -2123 -395 -1881 -389
rect -1815 -355 -1573 -349
rect -1815 -389 -1803 -355
rect -1585 -389 -1573 -355
rect -1815 -395 -1573 -389
rect -1507 -355 -1265 -349
rect -1507 -389 -1495 -355
rect -1277 -389 -1265 -355
rect -1507 -395 -1265 -389
rect -1199 -355 -957 -349
rect -1199 -389 -1187 -355
rect -969 -389 -957 -355
rect -1199 -395 -957 -389
rect -891 -355 -649 -349
rect -891 -389 -879 -355
rect -661 -389 -649 -355
rect -891 -395 -649 -389
rect -583 -355 -341 -349
rect -583 -389 -571 -355
rect -353 -389 -341 -355
rect -583 -395 -341 -389
rect -275 -355 -33 -349
rect -275 -389 -263 -355
rect -45 -389 -33 -355
rect -275 -395 -33 -389
rect 33 -355 275 -349
rect 33 -389 45 -355
rect 263 -389 275 -355
rect 33 -395 275 -389
rect 341 -355 583 -349
rect 341 -389 353 -355
rect 571 -389 583 -355
rect 341 -395 583 -389
rect 649 -355 891 -349
rect 649 -389 661 -355
rect 879 -389 891 -355
rect 649 -395 891 -389
rect 957 -355 1199 -349
rect 957 -389 969 -355
rect 1187 -389 1199 -355
rect 957 -395 1199 -389
rect 1265 -355 1507 -349
rect 1265 -389 1277 -355
rect 1495 -389 1507 -355
rect 1265 -395 1507 -389
rect 1573 -355 1815 -349
rect 1573 -389 1585 -355
rect 1803 -389 1815 -355
rect 1573 -395 1815 -389
rect 1881 -355 2123 -349
rect 1881 -389 1893 -355
rect 2111 -389 2123 -355
rect 1881 -395 2123 -389
rect 2189 -355 2431 -349
rect 2189 -389 2201 -355
rect 2419 -389 2431 -355
rect 2189 -395 2431 -389
rect 2497 -355 2739 -349
rect 2497 -389 2509 -355
rect 2727 -389 2739 -355
rect 2497 -395 2739 -389
rect 2805 -355 3047 -349
rect 2805 -389 2817 -355
rect 3035 -389 3047 -355
rect 2805 -395 3047 -389
rect 3113 -355 3355 -349
rect 3113 -389 3125 -355
rect 3343 -389 3355 -355
rect 3113 -395 3355 -389
rect 3421 -355 3663 -349
rect 3421 -389 3433 -355
rect 3651 -389 3663 -355
rect 3421 -395 3663 -389
rect 3729 -355 3971 -349
rect 3729 -389 3741 -355
rect 3959 -389 3971 -355
rect 3729 -395 3971 -389
rect 4037 -355 4279 -349
rect 4037 -389 4049 -355
rect 4267 -389 4279 -355
rect 4037 -395 4279 -389
rect 4345 -355 4587 -349
rect 4345 -389 4357 -355
rect 4575 -389 4587 -355
rect 4345 -395 4587 -389
rect 4653 -355 4895 -349
rect 4653 -389 4665 -355
rect 4883 -389 4895 -355
rect 4653 -395 4895 -389
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.4375 l 1.25 m 1 nf 32 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
