magic
tech sky130A
magscale 1 2
timestamp 1770023980
<< error_p >>
rect -2559 1038 2559 1042
rect -2559 -970 -2529 1038
rect -2493 972 2493 976
rect -2493 -904 -2463 972
rect 2463 -904 2493 972
rect -2344 -951 -2276 -945
rect -2036 -951 -1968 -945
rect -1728 -951 -1660 -945
rect -1420 -951 -1352 -945
rect -1112 -951 -1044 -945
rect -804 -951 -736 -945
rect -496 -951 -428 -945
rect -188 -951 -120 -945
rect 120 -951 188 -945
rect 428 -951 496 -945
rect 736 -951 804 -945
rect 1044 -951 1112 -945
rect 1352 -951 1420 -945
rect 1660 -951 1728 -945
rect 1968 -951 2036 -945
rect 2276 -951 2344 -945
rect -2344 -985 -2332 -951
rect -2036 -985 -2024 -951
rect -1728 -985 -1716 -951
rect -1420 -985 -1408 -951
rect -1112 -985 -1100 -951
rect -804 -985 -792 -951
rect -496 -985 -484 -951
rect -188 -985 -176 -951
rect 120 -972 132 -951
rect -2344 -991 -2276 -985
rect -2036 -991 -1968 -985
rect -1728 -991 -1660 -985
rect -1420 -991 -1352 -985
rect -1112 -991 -1044 -985
rect -804 -991 -736 -985
rect -496 -991 -428 -985
rect -188 -991 -120 -985
rect 120 -991 188 -972
rect 428 -985 440 -951
rect 736 -985 748 -951
rect 1044 -985 1056 -951
rect 1352 -985 1364 -951
rect 1660 -985 1672 -951
rect 1968 -985 1980 -951
rect 2276 -985 2288 -951
rect 2529 -970 2559 1038
rect 428 -991 496 -985
rect 736 -991 804 -985
rect 1044 -991 1112 -985
rect 1352 -991 1420 -985
rect 1660 -991 1728 -985
rect 1968 -991 2036 -985
rect 2276 -991 2344 -985
rect 92 -1019 200 -1000
<< nwell >>
rect -2529 -1004 2529 1038
<< mvpmos >>
rect -2435 -904 -2185 976
rect -2127 -904 -1877 976
rect -1819 -904 -1569 976
rect -1511 -904 -1261 976
rect -1203 -904 -953 976
rect -895 -904 -645 976
rect -587 -904 -337 976
rect -279 -904 -29 976
rect 29 -904 279 976
rect 337 -904 587 976
rect 645 -904 895 976
rect 953 -904 1203 976
rect 1261 -904 1511 976
rect 1569 -904 1819 976
rect 1877 -904 2127 976
rect 2185 -904 2435 976
<< mvpdiff >>
rect -2493 964 -2435 976
rect -2493 -892 -2481 964
rect -2447 -892 -2435 964
rect -2493 -904 -2435 -892
rect -2185 964 -2127 976
rect -2185 -892 -2173 964
rect -2139 -892 -2127 964
rect -2185 -904 -2127 -892
rect -1877 964 -1819 976
rect -1877 -892 -1865 964
rect -1831 -892 -1819 964
rect -1877 -904 -1819 -892
rect -1569 964 -1511 976
rect -1569 -892 -1557 964
rect -1523 -892 -1511 964
rect -1569 -904 -1511 -892
rect -1261 964 -1203 976
rect -1261 -892 -1249 964
rect -1215 -892 -1203 964
rect -1261 -904 -1203 -892
rect -953 964 -895 976
rect -953 -892 -941 964
rect -907 -892 -895 964
rect -953 -904 -895 -892
rect -645 964 -587 976
rect -645 -892 -633 964
rect -599 -892 -587 964
rect -645 -904 -587 -892
rect -337 964 -279 976
rect -337 -892 -325 964
rect -291 -892 -279 964
rect -337 -904 -279 -892
rect -29 964 29 976
rect -29 -892 -17 964
rect 17 -892 29 964
rect -29 -904 29 -892
rect 279 964 337 976
rect 279 -892 291 964
rect 325 -892 337 964
rect 279 -904 337 -892
rect 587 964 645 976
rect 587 -892 599 964
rect 633 -892 645 964
rect 587 -904 645 -892
rect 895 964 953 976
rect 895 -892 907 964
rect 941 -892 953 964
rect 895 -904 953 -892
rect 1203 964 1261 976
rect 1203 -892 1215 964
rect 1249 -892 1261 964
rect 1203 -904 1261 -892
rect 1511 964 1569 976
rect 1511 -892 1523 964
rect 1557 -892 1569 964
rect 1511 -904 1569 -892
rect 1819 964 1877 976
rect 1819 -892 1831 964
rect 1865 -892 1877 964
rect 1819 -904 1877 -892
rect 2127 964 2185 976
rect 2127 -892 2139 964
rect 2173 -892 2185 964
rect 2127 -904 2185 -892
rect 2435 964 2493 976
rect 2435 -892 2447 964
rect 2481 -892 2493 964
rect 2435 -904 2493 -892
<< mvpdiffc >>
rect -2481 -892 -2447 964
rect -2173 -892 -2139 964
rect -1865 -892 -1831 964
rect -1557 -892 -1523 964
rect -1249 -892 -1215 964
rect -941 -892 -907 964
rect -633 -892 -599 964
rect -325 -892 -291 964
rect -17 -892 17 964
rect 291 -892 325 964
rect 599 -892 633 964
rect 907 -892 941 964
rect 1215 -892 1249 964
rect 1523 -892 1557 964
rect 1831 -892 1865 964
rect 2139 -892 2173 964
rect 2447 -892 2481 964
<< poly >>
rect -2435 976 -2185 1002
rect -2127 976 -1877 1002
rect -1819 976 -1569 1002
rect -1511 976 -1261 1002
rect -1203 976 -953 1002
rect -895 976 -645 1002
rect -587 976 -337 1002
rect -279 976 -29 1002
rect 29 976 279 1002
rect 337 976 587 1002
rect 645 976 895 1002
rect 953 976 1203 1002
rect 1261 976 1511 1002
rect 1569 976 1819 1002
rect 1877 976 2127 1002
rect 2185 976 2435 1002
rect -2435 -951 -2185 -904
rect -2435 -968 -2332 -951
rect -2348 -985 -2332 -968
rect -2288 -968 -2185 -951
rect -2127 -951 -1877 -904
rect -2127 -968 -2024 -951
rect -2288 -985 -2272 -968
rect -2348 -1001 -2272 -985
rect -2040 -985 -2024 -968
rect -1980 -968 -1877 -951
rect -1819 -951 -1569 -904
rect -1819 -968 -1716 -951
rect -1980 -985 -1964 -968
rect -2040 -1001 -1964 -985
rect -1732 -985 -1716 -968
rect -1672 -968 -1569 -951
rect -1511 -951 -1261 -904
rect -1511 -968 -1408 -951
rect -1672 -985 -1656 -968
rect -1732 -1001 -1656 -985
rect -1424 -985 -1408 -968
rect -1364 -968 -1261 -951
rect -1203 -951 -953 -904
rect -1203 -968 -1100 -951
rect -1364 -985 -1348 -968
rect -1424 -1001 -1348 -985
rect -1116 -985 -1100 -968
rect -1056 -968 -953 -951
rect -895 -951 -645 -904
rect -895 -968 -792 -951
rect -1056 -985 -1040 -968
rect -1116 -1001 -1040 -985
rect -808 -985 -792 -968
rect -748 -968 -645 -951
rect -587 -951 -337 -904
rect -587 -968 -484 -951
rect -748 -985 -732 -968
rect -808 -1001 -732 -985
rect -500 -985 -484 -968
rect -440 -968 -337 -951
rect -279 -951 -29 -904
rect -279 -968 -176 -951
rect -440 -985 -424 -968
rect -500 -1001 -424 -985
rect -192 -985 -176 -968
rect -132 -968 -29 -951
rect 29 -951 279 -904
rect 29 -968 132 -951
rect -132 -985 -116 -968
rect -192 -1001 -116 -985
rect 116 -985 132 -968
rect 176 -968 279 -951
rect 337 -951 587 -904
rect 337 -968 440 -951
rect 176 -985 192 -968
rect 116 -1001 192 -985
rect 424 -985 440 -968
rect 484 -968 587 -951
rect 645 -951 895 -904
rect 645 -968 748 -951
rect 484 -985 500 -968
rect 424 -1001 500 -985
rect 732 -985 748 -968
rect 792 -968 895 -951
rect 953 -951 1203 -904
rect 953 -968 1056 -951
rect 792 -985 808 -968
rect 732 -1001 808 -985
rect 1040 -985 1056 -968
rect 1100 -968 1203 -951
rect 1261 -951 1511 -904
rect 1261 -968 1364 -951
rect 1100 -985 1116 -968
rect 1040 -1001 1116 -985
rect 1348 -985 1364 -968
rect 1408 -968 1511 -951
rect 1569 -951 1819 -904
rect 1569 -968 1672 -951
rect 1408 -985 1424 -968
rect 1348 -1001 1424 -985
rect 1656 -985 1672 -968
rect 1716 -968 1819 -951
rect 1877 -951 2127 -904
rect 1877 -968 1980 -951
rect 1716 -985 1732 -968
rect 1656 -1001 1732 -985
rect 1964 -985 1980 -968
rect 2024 -968 2127 -951
rect 2185 -951 2435 -904
rect 2185 -968 2288 -951
rect 2024 -985 2040 -968
rect 1964 -1001 2040 -985
rect 2272 -985 2288 -968
rect 2332 -968 2435 -951
rect 2332 -985 2348 -968
rect 2272 -1001 2348 -985
<< polycont >>
rect -2332 -985 -2288 -951
rect -2024 -985 -1980 -951
rect -1716 -985 -1672 -951
rect -1408 -985 -1364 -951
rect -1100 -985 -1056 -951
rect -792 -985 -748 -951
rect -484 -985 -440 -951
rect -176 -985 -132 -951
rect 132 -985 176 -951
rect 440 -985 484 -951
rect 748 -985 792 -951
rect 1056 -985 1100 -951
rect 1364 -985 1408 -951
rect 1672 -985 1716 -951
rect 1980 -985 2024 -951
rect 2288 -985 2332 -951
<< locali >>
rect -2481 964 -2447 980
rect -2481 -908 -2447 -892
rect -2173 964 -2139 980
rect -2173 -908 -2139 -892
rect -1865 964 -1831 980
rect -1865 -908 -1831 -892
rect -1557 964 -1523 980
rect -1557 -908 -1523 -892
rect -1249 964 -1215 980
rect -1249 -908 -1215 -892
rect -941 964 -907 980
rect -941 -908 -907 -892
rect -633 964 -599 980
rect -633 -908 -599 -892
rect -325 964 -291 980
rect -325 -908 -291 -892
rect -17 964 17 980
rect -17 -908 17 -892
rect 291 964 325 980
rect 291 -908 325 -892
rect 599 964 633 980
rect 599 -908 633 -892
rect 907 964 941 980
rect 907 -908 941 -892
rect 1215 964 1249 980
rect 1215 -908 1249 -892
rect 1523 964 1557 980
rect 1523 -908 1557 -892
rect 1831 964 1865 980
rect 1831 -908 1865 -892
rect 2139 964 2173 980
rect 2139 -908 2173 -892
rect 2447 964 2481 980
rect 2447 -908 2481 -892
rect -2348 -985 -2332 -951
rect -2288 -985 -2272 -951
rect -2040 -985 -2024 -951
rect -1980 -985 -1964 -951
rect -1732 -985 -1716 -951
rect -1672 -985 -1656 -951
rect -1424 -985 -1408 -951
rect -1364 -985 -1348 -951
rect -1116 -985 -1100 -951
rect -1056 -985 -1040 -951
rect -808 -985 -792 -951
rect -748 -985 -732 -951
rect -500 -985 -484 -951
rect -440 -985 -424 -951
rect -192 -985 -176 -951
rect -132 -985 -116 -951
rect 116 -985 132 -951
rect 176 -985 192 -951
rect 424 -985 440 -951
rect 484 -985 500 -951
rect 732 -985 748 -951
rect 792 -985 808 -951
rect 1040 -985 1056 -951
rect 1100 -985 1116 -951
rect 1348 -985 1364 -951
rect 1408 -985 1424 -951
rect 1656 -985 1672 -951
rect 1716 -985 1732 -951
rect 1964 -985 1980 -951
rect 2024 -985 2040 -951
rect 2272 -985 2288 -951
rect 2332 -985 2348 -951
<< viali >>
rect -2481 -892 -2447 964
rect -2173 -892 -2139 964
rect -1865 -892 -1831 964
rect -1557 -892 -1523 964
rect -1249 -892 -1215 964
rect -941 -892 -907 964
rect -633 -892 -599 964
rect -325 -892 -291 964
rect -17 -892 17 964
rect 291 -892 325 964
rect 599 -892 633 964
rect 907 -892 941 964
rect 1215 -892 1249 964
rect 1523 -892 1557 964
rect 1831 -892 1865 964
rect 2139 -892 2173 964
rect 2447 -892 2481 964
rect -2332 -985 -2288 -951
rect -2024 -985 -1980 -951
rect -1716 -985 -1672 -951
rect -1408 -985 -1364 -951
rect -1100 -985 -1056 -951
rect -792 -985 -748 -951
rect -484 -985 -440 -951
rect -176 -985 -132 -951
rect 132 -985 176 -951
rect 440 -985 484 -951
rect 748 -985 792 -951
rect 1056 -985 1100 -951
rect 1364 -985 1408 -951
rect 1672 -985 1716 -951
rect 1980 -985 2024 -951
rect 2288 -985 2332 -951
<< metal1 >>
rect -2487 964 -2441 976
rect -2487 -892 -2481 964
rect -2447 -892 -2441 964
rect -2487 -904 -2441 -892
rect -2179 964 -2133 976
rect -2179 -892 -2173 964
rect -2139 -892 -2133 964
rect -2179 -904 -2133 -892
rect -1871 964 -1825 976
rect -1871 -892 -1865 964
rect -1831 -892 -1825 964
rect -1871 -904 -1825 -892
rect -1563 964 -1517 976
rect -1563 -892 -1557 964
rect -1523 -892 -1517 964
rect -1563 -904 -1517 -892
rect -1255 964 -1209 976
rect -1255 -892 -1249 964
rect -1215 -892 -1209 964
rect -1255 -904 -1209 -892
rect -947 964 -901 976
rect -947 -892 -941 964
rect -907 -892 -901 964
rect -947 -904 -901 -892
rect -639 964 -593 976
rect -639 -892 -633 964
rect -599 -892 -593 964
rect -639 -904 -593 -892
rect -331 964 -285 976
rect -331 -892 -325 964
rect -291 -892 -285 964
rect -331 -904 -285 -892
rect -23 964 23 976
rect -23 -892 -17 964
rect 17 200 23 964
rect 285 964 331 976
rect 17 0 200 200
rect 17 -200 23 0
rect 17 -400 200 -200
rect 17 -600 23 -400
rect 17 -800 200 -600
rect 17 -892 23 -800
rect -23 -904 23 -892
rect 285 -892 291 964
rect 325 -892 331 964
rect 285 -904 331 -892
rect 593 964 639 976
rect 593 -892 599 964
rect 633 -892 639 964
rect 593 -904 639 -892
rect 901 964 947 976
rect 901 -892 907 964
rect 941 -892 947 964
rect 901 -904 947 -892
rect 1209 964 1255 976
rect 1209 -892 1215 964
rect 1249 -892 1255 964
rect 1209 -904 1255 -892
rect 1517 964 1563 976
rect 1517 -892 1523 964
rect 1557 -892 1563 964
rect 1517 -904 1563 -892
rect 1825 964 1871 976
rect 1825 -892 1831 964
rect 1865 -892 1871 964
rect 1825 -904 1871 -892
rect 2133 964 2179 976
rect 2133 -892 2139 964
rect 2173 -892 2179 964
rect 2133 -904 2179 -892
rect 2441 964 2487 976
rect 2441 -892 2447 964
rect 2481 -892 2487 964
rect 2441 -904 2487 -892
rect -2344 -951 -2276 -945
rect -2344 -985 -2332 -951
rect -2288 -985 -2276 -951
rect -2344 -991 -2276 -985
rect -2036 -951 -1968 -945
rect -2036 -985 -2024 -951
rect -1980 -985 -1968 -951
rect -2036 -991 -1968 -985
rect -1728 -951 -1660 -945
rect -1728 -985 -1716 -951
rect -1672 -985 -1660 -951
rect -1728 -991 -1660 -985
rect -1420 -951 -1352 -945
rect -1420 -985 -1408 -951
rect -1364 -985 -1352 -951
rect -1420 -991 -1352 -985
rect -1112 -951 -1044 -945
rect -1112 -985 -1100 -951
rect -1056 -985 -1044 -951
rect -1112 -991 -1044 -985
rect -804 -951 -736 -945
rect -804 -985 -792 -951
rect -748 -985 -736 -951
rect -804 -991 -736 -985
rect -496 -951 -428 -945
rect -496 -985 -484 -951
rect -440 -985 -428 -951
rect -496 -991 -428 -985
rect -188 -951 -120 -945
rect -188 -985 -176 -951
rect -132 -985 -120 -951
rect -188 -991 -120 -985
rect 120 -951 188 -945
rect 120 -985 132 -951
rect 176 -985 188 -951
rect 120 -991 188 -985
rect 428 -951 496 -945
rect 428 -985 440 -951
rect 484 -985 496 -951
rect 428 -991 496 -985
rect 736 -951 804 -945
rect 736 -985 748 -951
rect 792 -985 804 -951
rect 736 -991 804 -985
rect 1044 -951 1112 -945
rect 1044 -985 1056 -951
rect 1100 -985 1112 -951
rect 1044 -991 1112 -985
rect 1352 -951 1420 -945
rect 1352 -985 1364 -951
rect 1408 -985 1420 -951
rect 1352 -991 1420 -985
rect 1660 -951 1728 -945
rect 1660 -985 1672 -951
rect 1716 -985 1728 -951
rect 1660 -991 1728 -985
rect 1968 -951 2036 -945
rect 1968 -985 1980 -951
rect 2024 -985 2036 -951
rect 1968 -991 2036 -985
rect 2276 -951 2344 -945
rect 2276 -985 2288 -951
rect 2332 -985 2344 -951
rect 2276 -991 2344 -985
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
rect 0 -8800 200 -8600
rect 0 -9200 200 -9000
rect 0 -9600 200 -9400
rect 0 -10000 200 -9800
rect 0 -10400 200 -10200
rect 0 -10800 200 -10600
rect 0 -11200 200 -11000
rect 0 -11600 200 -11400
rect 0 -12000 200 -11800
rect 0 -12400 200 -12200
rect 0 -12800 200 -12600
rect 0 -13200 200 -13000
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X0
timestamp 0
transform 1 0 -2271 0 1 -12058
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X1
timestamp 0
transform 1 0 -1600 0 1 -12153
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X2
timestamp 0
transform 1 0 -929 0 1 -12248
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X3
timestamp 0
transform 1 0 -258 0 1 -12343
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X4
timestamp 0
transform 1 0 413 0 1 -12438
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X5
timestamp 0
transform 1 0 1084 0 1 -12533
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_QQM44N  X6
timestamp 0
transform 1 0 1755 0 1 -12628
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X7
timestamp 0
transform 1 0 2426 0 1 -12723
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X8
timestamp 0
transform 1 0 3097 0 1 -12818
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_NDJLD9  X9
timestamp 0
transform 1 0 3768 0 1 -12913
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X10
timestamp 0
transform 1 0 4439 0 1 -13008
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X11
timestamp 0
transform 1 0 5110 0 1 -13103
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X12
timestamp 0
transform 1 0 5781 0 1 -13198
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X13
timestamp 0
transform 1 0 6452 0 1 -13293
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X14
timestamp 0
transform 1 0 7123 0 1 -13388
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_W34X5V  X15
timestamp 0
transform 1 0 7794 0 1 -13483
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 a_n337_n904#
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 a_n587_n968#
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 a_n953_n904#
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 {}
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 a_645_n968#
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 a_29_n968#
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 a_1261_n968#
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 a_1569_n968#
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 w_n2529_n1004#
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 a_n2185_n904#
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 a_2435_n904#
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 a_n2435_n968#
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 a_279_n904#
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 a_895_n904#
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 a_1511_n904#
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 a_n1261_n904#
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 a_n1569_n904#
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 a_n1511_n968#
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 {}
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 a_n1819_n968#
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 256 0 0 0 a_n279_n968#
port 21 nsew
flabel metal1 0 -8800 200 -8600 0 FreeSans 256 0 0 0 a_n29_n904#
port 22 nsew
flabel metal1 0 -9200 200 -9000 0 FreeSans 256 0 0 0 a_n895_n968#
port 23 nsew
flabel metal1 0 -9600 200 -9400 0 FreeSans 256 0 0 0 a_337_n968#
port 24 nsew
flabel metal1 0 -10000 200 -9800 0 FreeSans 256 0 0 0 a_953_n968#
port 25 nsew
flabel metal1 0 -10400 200 -10200 0 FreeSans 256 0 0 0 a_2127_n904#
port 26 nsew
flabel metal1 0 -10800 200 -10600 0 FreeSans 256 0 0 0 {}
port 27 nsew
flabel metal1 0 -11200 200 -11000 0 FreeSans 256 0 0 0 a_1877_n968#
port 28 nsew
flabel metal1 0 -11600 200 -11400 0 FreeSans 256 0 0 0 a_n2493_n904#
port 29 nsew
flabel metal1 0 -12000 200 -11800 0 FreeSans 256 0 0 0 a_n2127_n968#
port 30 nsew
flabel metal1 0 -12400 200 -12200 0 FreeSans 256 0 0 0 a_1203_n904#
port 31 nsew
flabel metal1 0 -12800 200 -12600 0 FreeSans 256 0 0 0 a_n1203_n968#
port 32 nsew
flabel metal1 0 -13200 200 -13000 0 FreeSans 256 0 0 0 a_2185_n968#
port 33 nsew
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9.4 l 1.25 m 1 nf 16 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
