magic
tech sky130A
magscale 1 2
timestamp 1769402310
<< error_p >>
rect -377 166 -319 172
rect -145 166 -87 172
rect 87 166 145 172
rect 319 166 377 172
rect -377 132 -365 166
rect -145 132 -133 166
rect 87 132 99 166
rect 319 132 331 166
rect -377 126 -319 132
rect -145 126 -87 132
rect 87 126 145 132
rect 319 126 377 132
<< nmos >>
rect -378 -156 -318 94
rect -146 -156 -86 94
rect 86 -156 146 94
rect 318 -156 378 94
<< ndiff >>
rect -436 82 -378 94
rect -436 -144 -424 82
rect -390 -144 -378 82
rect -436 -156 -378 -144
rect -318 82 -260 94
rect -318 -144 -306 82
rect -272 -144 -260 82
rect -318 -156 -260 -144
rect -204 82 -146 94
rect -204 -144 -192 82
rect -158 -144 -146 82
rect -204 -156 -146 -144
rect -86 82 -28 94
rect -86 -144 -74 82
rect -40 -144 -28 82
rect -86 -156 -28 -144
rect 28 82 86 94
rect 28 -144 40 82
rect 74 -144 86 82
rect 28 -156 86 -144
rect 146 82 204 94
rect 146 -144 158 82
rect 192 -144 204 82
rect 146 -156 204 -144
rect 260 82 318 94
rect 260 -144 272 82
rect 306 -144 318 82
rect 260 -156 318 -144
rect 378 82 436 94
rect 378 -144 390 82
rect 424 -144 436 82
rect 378 -156 436 -144
<< ndiffc >>
rect -424 -144 -390 82
rect -306 -144 -272 82
rect -192 -144 -158 82
rect -74 -144 -40 82
rect 40 -144 74 82
rect 158 -144 192 82
rect 272 -144 306 82
rect 390 -144 424 82
<< poly >>
rect -381 166 -315 182
rect -381 132 -365 166
rect -331 132 -315 166
rect -381 116 -315 132
rect -149 166 -83 182
rect -149 132 -133 166
rect -99 132 -83 166
rect -149 116 -83 132
rect 83 166 149 182
rect 83 132 99 166
rect 133 132 149 166
rect 83 116 149 132
rect 315 166 381 182
rect 315 132 331 166
rect 365 132 381 166
rect 315 116 381 132
rect -378 94 -318 116
rect -146 94 -86 116
rect 86 94 146 116
rect 318 94 378 116
rect -378 -182 -318 -156
rect -146 -182 -86 -156
rect 86 -182 146 -156
rect 318 -182 378 -156
<< polycont >>
rect -365 132 -331 166
rect -133 132 -99 166
rect 99 132 133 166
rect 331 132 365 166
<< locali >>
rect -381 132 -365 166
rect -331 132 -315 166
rect -149 132 -133 166
rect -99 132 -83 166
rect 83 132 99 166
rect 133 132 149 166
rect 315 132 331 166
rect 365 132 381 166
rect -424 82 -390 98
rect -424 -160 -390 -144
rect -306 82 -272 98
rect -306 -160 -272 -144
rect -192 82 -158 98
rect -192 -160 -158 -144
rect -74 82 -40 98
rect -74 -160 -40 -144
rect 40 82 74 98
rect 40 -160 74 -144
rect 158 82 192 98
rect 158 -160 192 -144
rect 272 82 306 98
rect 272 -160 306 -144
rect 390 82 424 98
rect 390 -160 424 -144
<< viali >>
rect -365 132 -331 166
rect -133 132 -99 166
rect 99 132 133 166
rect 331 132 365 166
rect -424 -144 -390 82
rect -306 -144 -272 82
rect -192 -144 -158 82
rect -74 -144 -40 82
rect 40 -144 74 82
rect 158 -144 192 82
rect 272 -144 306 82
rect 390 -144 424 82
<< metal1 >>
rect -377 166 -319 172
rect -377 132 -365 166
rect -331 132 -319 166
rect -377 126 -319 132
rect -145 166 -87 172
rect -145 132 -133 166
rect -99 132 -87 166
rect -145 126 -87 132
rect 87 166 145 172
rect 87 132 99 166
rect 133 132 145 166
rect 87 126 145 132
rect 319 166 377 172
rect 319 132 331 166
rect 365 132 377 166
rect 319 126 377 132
rect -430 82 -384 94
rect -430 -144 -424 82
rect -390 -144 -384 82
rect -430 -156 -384 -144
rect -312 82 -266 94
rect -312 -144 -306 82
rect -272 -144 -266 82
rect -312 -156 -266 -144
rect -198 82 -152 94
rect -198 -144 -192 82
rect -158 -144 -152 82
rect -198 -156 -152 -144
rect -80 82 -34 94
rect -80 -144 -74 82
rect -40 -144 -34 82
rect -80 -156 -34 -144
rect 34 82 80 94
rect 34 -144 40 82
rect 74 -144 80 82
rect 34 -156 80 -144
rect 152 82 198 94
rect 152 -144 158 82
rect 192 -144 198 82
rect 152 -156 198 -144
rect 266 82 312 94
rect 266 -144 272 82
rect 306 -144 312 82
rect 266 -156 312 -144
rect 384 82 430 94
rect 384 -144 390 82
rect 424 -144 430 82
rect 384 -156 430 -144
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.25 l 0.3 m 1 nf 4 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
