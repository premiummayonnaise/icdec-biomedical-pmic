* NGSPICE file created from two-stage-miller.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_V6JW4R a_n267_n536# a_29_n562# a_209_n536# a_n29_n536#
+ w_n467_n762# a_n209_n562#
X0 a_n29_n536# a_n209_n562# a_n267_n536# w_n467_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.9
X1 a_209_n536# a_29_n562# a_n29_n536# w_n467_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.9
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_RFPNS8 a_587_n964# a_1203_n964# a_337_n1061#
+ a_n279_n1061# a_953_n1061# a_n895_n1061# a_n1203_n1061# a_n337_n964# a_n953_n964#
+ a_29_n1061# a_279_n964# a_895_n964# w_n1461_n1262# a_n1261_n964# a_645_n1061# a_n587_n1061#
+ a_n645_n964# a_n29_n964#
X0 a_895_n964# a_645_n1061# a_587_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X1 a_n645_n964# a_n895_n1061# a_n953_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X2 a_n29_n964# a_n279_n1061# a_n337_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X3 a_n953_n964# a_n1203_n1061# a_n1261_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1.25
X4 a_1203_n964# a_953_n1061# a_895_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1.25
X5 a_587_n964# a_337_n1061# a_279_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X6 a_n337_n964# a_n587_n1061# a_n645_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
X7 a_279_n964# a_29_n1061# a_n29_n964# w_n1461_n1262# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1.25
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_S5VYLR a_n337_n904# a_n587_n968# a_n953_n904#
+ a_645_n968# a_29_n968# a_1261_n968# a_1569_n968# a_n2185_n904# a_2435_n904# a_n2435_n968#
+ a_279_n904# a_895_n904# a_1511_n904# a_n1261_n904# a_n1569_n904# a_n1511_n968# a_1819_n904#
+ a_n1819_n968# a_n279_n968# a_n29_n904# a_n645_n904# a_n895_n968# a_337_n968# a_953_n968#
+ w_n2693_n1202# a_2127_n904# a_1877_n968# a_n2493_n904# a_n2127_n968# a_587_n904#
+ a_1203_n904# a_n1203_n968# a_n1877_n904# a_2185_n968#
X0 a_n1877_n904# a_n2127_n968# a_n2185_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X1 a_895_n904# a_645_n968# a_587_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X2 a_n1569_n904# a_n1819_n968# a_n1877_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X3 a_n645_n904# a_n895_n968# a_n953_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X4 a_1819_n904# a_1569_n968# a_1511_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X5 a_n29_n904# a_n279_n968# a_n337_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X6 a_n2185_n904# a_n2435_n968# a_n2493_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=2.726 ps=19.38 w=9.4 l=1.25
X7 a_n953_n904# a_n1203_n968# a_n1261_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X8 a_1203_n904# a_953_n968# a_895_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X9 a_2435_n904# a_2185_n968# a_2127_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=2.726 pd=19.38 as=1.363 ps=9.69 w=9.4 l=1.25
X10 a_587_n904# a_337_n968# a_279_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X11 a_2127_n904# a_1877_n968# a_1819_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X12 a_n337_n904# a_n587_n968# a_n645_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X13 a_279_n904# a_29_n968# a_n29_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X14 a_n1261_n904# a_n1511_n968# a_n1569_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
X15 a_1511_n904# a_1261_n968# a_1203_n904# w_n2693_n1202# sky130_fd_pr__pfet_g5v0d10v5 ad=1.363 pd=9.69 as=1.363 ps=9.69 w=9.4 l=1.25
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DC2CKB a_n29_n440# a_29_n495# a_n187_n440# a_n129_n495#
+ a_187_n495# a_n287_n495# a_n345_n440# a_129_n440# a_287_n440# a_n479_n662#
X0 a_n187_n440# a_n287_n495# a_n345_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=1.3659 ps=10 w=4.71 l=0.5
X1 a_287_n440# a_187_n495# a_129_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3659 pd=10 as=0.68295 ps=5 w=4.71 l=0.5
X2 a_129_n440# a_29_n495# a_n29_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X3 a_n29_n440# a_n129_n495# a_n187_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2899RY a_n953_n781# a_2185_n807# a_n587_n807#
+ a_645_n807# a_29_n807# a_2435_n781# a_n2185_n781# a_1261_n807# a_1569_n807# a_279_n781#
+ a_895_n781# a_n2435_n807# a_n1261_n781# a_1511_n781# a_1819_n781# a_n1569_n781#
+ a_n29_n781# a_n645_n781# a_n1511_n807# a_n279_n807# a_n1819_n807# a_n895_n807# a_337_n807#
+ a_953_n807# a_2127_n781# a_n2493_n781# a_587_n781# a_1877_n807# a_n2627_n941# a_n2127_n807#
+ a_1203_n781# a_n1877_n781# a_n337_n781# a_n1203_n807#
X0 a_1511_n781# a_1261_n807# a_1203_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X1 a_n1261_n781# a_n1511_n807# a_n1569_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X2 a_n1877_n781# a_n2127_n807# a_n2185_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X3 a_895_n781# a_645_n807# a_587_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X4 a_n1569_n781# a_n1819_n807# a_n1877_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X5 a_n645_n781# a_n895_n807# a_n953_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X6 a_1819_n781# a_1569_n807# a_1511_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X7 a_n29_n781# a_n279_n807# a_n337_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X8 a_n953_n781# a_n1203_n807# a_n1261_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X9 a_2435_n781# a_2185_n807# a_2127_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=1.25
X10 a_n2185_n781# a_n2435_n807# a_n2493_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=1.25
X11 a_1203_n781# a_953_n807# a_895_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X12 a_587_n781# a_337_n807# a_279_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X13 a_2127_n781# a_1877_n807# a_1819_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X14 a_n337_n781# a_n587_n807# a_n645_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X15 a_279_n781# a_29_n807# a_n29_n781# a_n2627_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_A8KA9K a_n29_n440# a_29_n495# a_n187_n440# a_n129_n495#
+ a_187_n495# a_n287_n495# a_n345_n440# a_129_n440# a_287_n440# a_n479_n662#
X0 a_n187_n440# a_n287_n495# a_n345_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=1.3659 ps=10 w=4.71 l=0.5
X1 a_287_n440# a_187_n495# a_129_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3659 pd=10 as=0.68295 ps=5 w=4.71 l=0.5
X2 a_129_n440# a_29_n495# a_n29_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X3 a_n29_n440# a_n129_n495# a_n187_n440# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_N5GNFR a_n587_n807# a_29_n807# a_279_n781# a_n29_n781#
+ a_n645_n781# a_n779_n941# a_n279_n807# a_337_n807# a_587_n781# a_n337_n781#
X0 a_n29_n781# a_n279_n807# a_n337_n781# a_n779_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
X1 a_587_n781# a_337_n807# a_279_n781# a_n779_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=2.175 pd=15.58 as=1.0875 ps=7.79 w=7.5 l=1.25
X2 a_n337_n781# a_n587_n807# a_n645_n781# a_n779_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=2.175 ps=15.58 w=7.5 l=1.25
X3 a_279_n781# a_29_n807# a_n29_n781# a_n779_n941# sky130_fd_pr__nfet_g5v0d10v5 ad=1.0875 pd=7.79 as=1.0875 ps=7.79 w=7.5 l=1.25
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_X6KG9Z a_n345_n502# a_129_n502# a_29_n528# a_n129_n528#
+ a_287_n502# a_187_n528# a_n287_n528# a_n29_n502# a_n479_n662# a_n187_n502#
X0 a_287_n502# a_187_n528# a_129_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3659 pd=10 as=0.68295 ps=5 w=4.71 l=0.5
X1 a_129_n502# a_29_n528# a_n29_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X2 a_n29_n502# a_n129_n528# a_n187_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X3 a_n187_n502# a_n287_n528# a_n345_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=1.3659 ps=10 w=4.71 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_R7S84X m3_n2686_n21160# c1_n2646_n21120#
X0 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X1 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X2 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X3 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X4 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X5 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X6 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X7 c1_n2646_n21120# m3_n2686_n21160# sky130_fd_pr__cap_mim_m3_1 l=25 w=25
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PBQQNH a_n345_n502# a_129_n502# a_29_n528# a_n129_n528#
+ a_287_n502# a_187_n528# a_n287_n528# a_n29_n502# a_n479_n662# a_n187_n502#
X0 a_287_n502# a_187_n528# a_129_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3659 pd=10 as=0.68295 ps=5 w=4.71 l=0.5
X1 a_129_n502# a_29_n528# a_n29_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X2 a_n29_n502# a_n129_n528# a_n187_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=0.68295 ps=5 w=4.71 l=0.5
X3 a_n187_n502# a_n287_n528# a_n345_n502# a_n479_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.68295 pd=5 as=1.3659 ps=10 w=4.71 l=0.5
.ends

.subckt two-stage-miller VDD OUT VP VN IBIAS VSS
Xsky130_fd_pr__pfet_g5v0d10v5_V6JW4R_1 OUT VSS OUT m1_n2200_3200# VDD VSS sky130_fd_pr__pfet_g5v0d10v5_V6JW4R
Xsky130_fd_pr__pfet_g5v0d10v5_RFPNS8_0 OUT OUT m1_n1120_1120# m1_n1120_1120# m1_n1120_1120#
+ m1_n1120_1120# m1_n1120_1120# VDD VDD m1_n1120_1120# VDD VDD VDD OUT m1_n1120_1120#
+ m1_n1120_1120# OUT OUT sky130_fd_pr__pfet_g5v0d10v5_RFPNS8
XXM2 VDD m1_2160_1440# VDD m1_2160_1440# m1_2160_1440# m1_2160_1440# m1_2160_1440#
+ VDD m1_2160_1440# m1_2160_1440# VDD VDD VDD m1_2160_1440# VDD m1_2160_1440# m1_n1120_1120#
+ m1_2160_1440# m1_2160_1440# m1_2160_1440# m1_n1120_1120# m1_2160_1440# m1_2160_1440#
+ m1_2160_1440# VDD VDD m1_2160_1440# m1_2160_1440# m1_2160_1440# m1_n1120_1120# m1_2160_1440#
+ m1_2160_1440# m1_n1120_1120# m1_2160_1440# sky130_fd_pr__pfet_g5v0d10v5_S5VYLR
XXM3 m1_2160_1440# VP m1_2740_n3440# VP VP VP m1_2160_1440# m1_2740_n3440# m1_2160_1440#
+ VSS sky130_fd_pr__nfet_g5v0d10v5_DC2CKB
XXM5 VSS IBIAS IBIAS IBIAS IBIAS IBIAS VSS IBIAS IBIAS VSS VSS IBIAS IBIAS VSS m1_2740_n3440#
+ VSS IBIAS m1_2740_n3440# IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS VSS IBIAS m1_2740_n3440#
+ IBIAS VSS IBIAS IBIAS m1_2740_n3440# VSS IBIAS sky130_fd_pr__nfet_g5v0d10v5_2899RY
Xsky130_fd_pr__nfet_g5v0d10v5_A8KA9K_0 m1_n1120_1120# VN m1_2740_n3440# VN VN VN m1_n1120_1120#
+ m1_2740_n3440# m1_n1120_1120# VSS sky130_fd_pr__nfet_g5v0d10v5_A8KA9K
XXM7 OUT OUT m1_n1120_1120# m1_n1120_1120# m1_n1120_1120# m1_n1120_1120# m1_n1120_1120#
+ VDD VDD m1_n1120_1120# VDD VDD VDD OUT m1_n1120_1120# m1_n1120_1120# OUT OUT sky130_fd_pr__pfet_g5v0d10v5_RFPNS8
XXM8 IBIAS IBIAS VSS OUT OUT VSS IBIAS IBIAS OUT VSS sky130_fd_pr__nfet_g5v0d10v5_N5GNFR
Xsky130_fd_pr__nfet_g5v0d10v5_X6KG9Z_0 m1_2160_1440# m1_2740_n3440# VP VP m1_2160_1440#
+ VP VP m1_2160_1440# VSS m1_2740_n3440# sky130_fd_pr__nfet_g5v0d10v5_X6KG9Z
Xsky130_fd_pr__cap_mim_m3_1_R7S84X_0 m1_n1120_1120# m1_n2200_3200# sky130_fd_pr__cap_mim_m3_1_R7S84X
Xsky130_fd_pr__nfet_g5v0d10v5_N5GNFR_0 IBIAS IBIAS VSS OUT OUT VSS IBIAS IBIAS OUT
+ VSS sky130_fd_pr__nfet_g5v0d10v5_N5GNFR
Xsky130_fd_pr__nfet_g5v0d10v5_PBQQNH_0 m1_n1120_1120# m1_2740_n3440# VN VN m1_n1120_1120#
+ VN VN m1_n1120_1120# VSS m1_2740_n3440# sky130_fd_pr__nfet_g5v0d10v5_PBQQNH
Xsky130_fd_pr__pfet_g5v0d10v5_V6JW4R_0 OUT VSS OUT m1_n2200_3200# VDD VSS sky130_fd_pr__pfet_g5v0d10v5_V6JW4R
.ends

