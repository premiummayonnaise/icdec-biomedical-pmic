magic
tech sky130A
magscale 1 2
timestamp 1769952370
<< pwell >>
rect 1300 -300 6900 3600
<< psubdiff >>
rect 1300 3580 6900 3600
rect 1300 3520 1410 3580
rect 6810 3520 6900 3580
rect 1300 3500 6900 3520
rect 1300 3490 1400 3500
rect 1300 -190 1320 3490
rect 1380 -190 1400 3490
rect 6800 3480 6900 3500
rect 1600 3370 2700 3400
rect 1600 3330 1620 3370
rect 2680 3330 2700 3370
rect 1600 3300 2700 3330
rect 1600 2000 1700 3300
rect 2600 2000 2700 3300
rect 1600 1900 2700 2000
rect 2800 3370 3900 3400
rect 2800 3330 2820 3370
rect 3880 3330 3900 3370
rect 2800 3300 3900 3330
rect 2800 2000 2900 3300
rect 3800 2000 3900 3300
rect 2800 1900 3900 2000
rect 4300 3370 5400 3400
rect 4300 3330 4320 3370
rect 5380 3330 5400 3370
rect 4300 3300 5400 3330
rect 4300 2000 4400 3300
rect 5300 2000 5400 3300
rect 4300 1900 5400 2000
rect 5500 3370 6600 3400
rect 5500 3330 5520 3370
rect 6580 3330 6600 3370
rect 5500 3300 6600 3330
rect 5500 2000 5600 3300
rect 6500 2000 6600 3300
rect 5500 1900 6600 2000
rect 1600 1300 2700 1400
rect 1600 0 1700 1300
rect 2600 0 2700 1300
rect 1600 -30 2700 0
rect 1600 -70 1620 -30
rect 2680 -70 2700 -30
rect 1600 -100 2700 -70
rect 2800 1300 3900 1400
rect 2800 0 2900 1300
rect 3800 0 3900 1300
rect 2800 -30 3900 0
rect 2800 -70 2820 -30
rect 3880 -70 3900 -30
rect 2800 -100 3900 -70
rect 4300 1300 5400 1400
rect 4300 0 4400 1300
rect 5300 0 5400 1300
rect 4300 -30 5400 0
rect 4300 -70 4320 -30
rect 5380 -70 5400 -30
rect 4300 -100 5400 -70
rect 5500 1300 6600 1400
rect 5500 0 5600 1300
rect 6500 0 6600 1300
rect 5500 -30 6600 0
rect 5500 -70 5520 -30
rect 6580 -70 6600 -30
rect 5500 -100 6600 -70
rect 1300 -200 1400 -190
rect 6800 -190 6820 3480
rect 6880 -190 6900 3480
rect 6800 -200 6900 -190
rect 1300 -220 6900 -200
rect 1300 -280 1400 -220
rect 6800 -280 6900 -220
rect 1300 -300 6900 -280
<< psubdiffcont >>
rect 1410 3520 6810 3580
rect 1320 -190 1380 3490
rect 1620 3330 2680 3370
rect 2820 3330 3880 3370
rect 4320 3330 5380 3370
rect 5520 3330 6580 3370
rect 1620 -70 2680 -30
rect 2820 -70 3880 -30
rect 4320 -70 5380 -30
rect 5520 -70 6580 -30
rect 6820 -190 6880 3480
rect 1400 -280 6800 -220
<< poly >>
rect 1720 2100 1780 3120
rect 2510 2100 2570 3120
rect 2920 2100 2980 3120
rect 3710 2090 3770 3110
rect 4420 2100 4480 3120
rect 5210 2100 5270 3120
rect 5620 2100 5680 3120
rect 6410 2100 6470 3120
rect 1720 200 1780 1220
rect 2510 200 2570 1220
rect 2920 200 2980 1220
rect 3720 200 3780 1220
rect 4420 200 4480 1200
rect 5210 200 5270 1200
rect 5620 200 5680 1200
rect 6410 210 6470 1210
<< locali >>
rect 1300 3580 6900 3600
rect 1300 3520 1410 3580
rect 6810 3520 6900 3580
rect 1300 3500 6900 3520
rect 1300 3490 1400 3500
rect 1300 -190 1320 3490
rect 1380 3402 1400 3490
rect 6800 3480 6900 3500
rect 6800 3402 6820 3480
rect 1380 3400 1720 3402
rect 6480 3400 6820 3402
rect 1380 3370 3900 3400
rect 1380 3330 1620 3370
rect 2680 3330 2820 3370
rect 3880 3330 3900 3370
rect 1380 3300 3900 3330
rect 3960 3360 4240 3400
rect 3960 3300 4020 3360
rect 4080 3300 4120 3360
rect 4180 3300 4240 3360
rect 4300 3370 6820 3400
rect 4300 3330 4320 3370
rect 5380 3330 5520 3370
rect 6580 3330 6820 3370
rect 4300 3300 6820 3330
rect 1380 0 1400 3300
rect 3960 3260 4240 3300
rect 3000 3200 4020 3260
rect 4080 3200 4120 3260
rect 4180 3200 5200 3260
rect 3000 3160 5200 3200
rect 2080 1800 2200 3020
rect 3280 2200 3400 3160
rect 3900 3100 4020 3160
rect 4080 3100 4120 3160
rect 4180 3100 4300 3160
rect 3900 3060 4300 3100
rect 3900 3000 4020 3060
rect 4080 3000 4120 3060
rect 4180 3000 4300 3060
rect 3900 2960 4300 3000
rect 3900 2900 4020 2960
rect 4080 2900 4120 2960
rect 4180 2900 4300 2960
rect 3900 2860 4300 2900
rect 3900 2800 4020 2860
rect 4080 2800 4120 2860
rect 4180 2800 4300 2860
rect 3900 2760 4300 2800
rect 3900 2700 4020 2760
rect 4080 2700 4120 2760
rect 4180 2700 4300 2760
rect 3900 2660 4300 2700
rect 3900 2600 4020 2660
rect 4080 2600 4120 2660
rect 4180 2600 4300 2660
rect 3900 2560 4300 2600
rect 3900 2500 4020 2560
rect 4080 2500 4120 2560
rect 4180 2500 4300 2560
rect 3900 2460 4300 2500
rect 3900 2400 4020 2460
rect 4080 2400 4120 2460
rect 4180 2400 4300 2460
rect 3900 2360 4300 2400
rect 3900 2300 4020 2360
rect 4080 2300 4120 2360
rect 4180 2300 4300 2360
rect 3900 2260 4300 2300
rect 3900 2200 4020 2260
rect 4080 2200 4120 2260
rect 4180 2200 4300 2260
rect 4780 2200 4900 3160
rect 3900 2160 4300 2200
rect 3900 2100 4020 2160
rect 4080 2100 4120 2160
rect 4180 2100 4300 2160
rect 3900 1800 4300 2100
rect 5980 1800 6100 3020
rect 1500 1740 6700 1800
rect 1500 1680 1520 1740
rect 1580 1680 1620 1740
rect 1680 1680 1720 1740
rect 1780 1680 1820 1740
rect 1880 1680 1920 1740
rect 1980 1680 2020 1740
rect 2080 1680 2120 1740
rect 2180 1680 2220 1740
rect 2280 1680 2320 1740
rect 2380 1680 2420 1740
rect 2480 1680 2520 1740
rect 2580 1680 2620 1740
rect 2680 1680 2720 1740
rect 2780 1680 2820 1740
rect 2880 1680 2920 1740
rect 2980 1680 3020 1740
rect 3080 1680 3120 1740
rect 3180 1680 3220 1740
rect 3280 1680 3320 1740
rect 3380 1680 3420 1740
rect 3480 1680 3520 1740
rect 3580 1680 3620 1740
rect 3680 1680 3720 1740
rect 3780 1680 3820 1740
rect 3880 1680 3920 1740
rect 3980 1680 4020 1740
rect 4080 1680 4120 1740
rect 4180 1680 4220 1740
rect 4280 1680 4320 1740
rect 4380 1680 4420 1740
rect 4480 1680 4520 1740
rect 4580 1680 4620 1740
rect 4680 1680 4720 1740
rect 4780 1680 4820 1740
rect 4880 1680 4920 1740
rect 4980 1680 5020 1740
rect 5080 1680 5120 1740
rect 5180 1680 5220 1740
rect 5280 1680 5320 1740
rect 5380 1680 5420 1740
rect 5480 1680 5520 1740
rect 5580 1680 5620 1740
rect 5680 1680 5720 1740
rect 5780 1680 5820 1740
rect 5880 1680 5920 1740
rect 5980 1680 6020 1740
rect 6080 1680 6120 1740
rect 6180 1680 6220 1740
rect 6280 1680 6320 1740
rect 6380 1680 6420 1740
rect 6480 1680 6520 1740
rect 6580 1680 6620 1740
rect 6680 1680 6700 1740
rect 1500 1620 6700 1680
rect 1500 1560 1520 1620
rect 1580 1560 1620 1620
rect 1680 1560 1720 1620
rect 1780 1560 1820 1620
rect 1880 1560 1920 1620
rect 1980 1560 2020 1620
rect 2080 1560 2120 1620
rect 2180 1560 2220 1620
rect 2280 1560 2320 1620
rect 2380 1560 2420 1620
rect 2480 1560 2520 1620
rect 2580 1560 2620 1620
rect 2680 1560 2720 1620
rect 2780 1560 2820 1620
rect 2880 1560 2920 1620
rect 2980 1560 3020 1620
rect 3080 1560 3120 1620
rect 3180 1560 3220 1620
rect 3280 1560 3320 1620
rect 3380 1560 3420 1620
rect 3480 1560 3520 1620
rect 3580 1560 3620 1620
rect 3680 1560 3720 1620
rect 3780 1560 3820 1620
rect 3880 1560 3920 1620
rect 3980 1560 4020 1620
rect 4080 1560 4120 1620
rect 4180 1560 4220 1620
rect 4280 1560 4320 1620
rect 4380 1560 4420 1620
rect 4480 1560 4520 1620
rect 4580 1560 4620 1620
rect 4680 1560 4720 1620
rect 4780 1560 4820 1620
rect 4880 1560 4920 1620
rect 4980 1560 5020 1620
rect 5080 1560 5120 1620
rect 5180 1560 5220 1620
rect 5280 1560 5320 1620
rect 5380 1560 5420 1620
rect 5480 1560 5520 1620
rect 5580 1560 5620 1620
rect 5680 1560 5720 1620
rect 5780 1560 5820 1620
rect 5880 1560 5920 1620
rect 5980 1560 6020 1620
rect 6080 1560 6120 1620
rect 6180 1560 6220 1620
rect 6280 1560 6320 1620
rect 6380 1560 6420 1620
rect 6480 1560 6520 1620
rect 6580 1560 6620 1620
rect 6680 1560 6700 1620
rect 1500 1500 6700 1560
rect 2080 300 2200 1500
rect 3900 1200 4300 1500
rect 3900 1140 4020 1200
rect 4080 1140 4120 1200
rect 4180 1140 4300 1200
rect 3280 140 3400 1120
rect 3900 1100 4300 1140
rect 3900 1040 4020 1100
rect 4080 1040 4120 1100
rect 4180 1040 4300 1100
rect 3900 1000 4300 1040
rect 3900 940 4020 1000
rect 4080 940 4120 1000
rect 4180 940 4300 1000
rect 3900 900 4300 940
rect 3900 840 4020 900
rect 4080 840 4120 900
rect 4180 840 4300 900
rect 3900 800 4300 840
rect 3900 740 4020 800
rect 4080 740 4120 800
rect 4180 740 4300 800
rect 3900 700 4300 740
rect 3900 640 4020 700
rect 4080 640 4120 700
rect 4180 640 4300 700
rect 3900 600 4300 640
rect 3900 540 4020 600
rect 4080 540 4120 600
rect 4180 540 4300 600
rect 3900 500 4300 540
rect 3900 440 4020 500
rect 4080 440 4120 500
rect 4180 440 4300 500
rect 3900 400 4300 440
rect 3900 340 4020 400
rect 4080 340 4120 400
rect 4180 340 4300 400
rect 3900 300 4300 340
rect 3900 240 4020 300
rect 4080 240 4120 300
rect 4180 240 4300 300
rect 3900 200 4300 240
rect 3900 140 4020 200
rect 4080 140 4120 200
rect 4180 140 4300 200
rect 4800 140 4920 1120
rect 5980 300 6100 1500
rect 3000 100 5200 140
rect 3000 40 4020 100
rect 4080 40 4120 100
rect 4180 40 5200 100
rect 3960 0 4240 40
rect 6800 2 6820 3300
rect 6480 0 6820 2
rect 1380 -30 3900 0
rect 1380 -70 1620 -30
rect 2680 -70 2820 -30
rect 3880 -70 3900 -30
rect 1380 -100 3900 -70
rect 3960 -60 4020 0
rect 4080 -60 4120 0
rect 4180 -60 4240 0
rect 3960 -100 4240 -60
rect 4300 -30 6820 0
rect 4300 -70 4320 -30
rect 5380 -70 5520 -30
rect 6580 -70 6820 -30
rect 4300 -100 6820 -70
rect 1380 -102 1720 -100
rect 1380 -190 1400 -102
rect 1300 -200 1400 -190
rect 6800 -190 6820 -100
rect 6880 -190 6900 3480
rect 6800 -200 6900 -190
rect 1300 -220 6900 -200
rect 1300 -280 1320 -220
rect 1380 -280 1400 -220
rect 6800 -280 6900 -220
rect 1300 -300 6900 -280
<< viali >>
rect 4020 3300 4080 3360
rect 4120 3300 4180 3360
rect 4020 3200 4080 3260
rect 4120 3200 4180 3260
rect 4020 3100 4080 3160
rect 4120 3100 4180 3160
rect 4020 3000 4080 3060
rect 4120 3000 4180 3060
rect 4020 2900 4080 2960
rect 4120 2900 4180 2960
rect 4020 2800 4080 2860
rect 4120 2800 4180 2860
rect 4020 2700 4080 2760
rect 4120 2700 4180 2760
rect 4020 2600 4080 2660
rect 4120 2600 4180 2660
rect 4020 2500 4080 2560
rect 4120 2500 4180 2560
rect 4020 2400 4080 2460
rect 4120 2400 4180 2460
rect 4020 2300 4080 2360
rect 4120 2300 4180 2360
rect 4020 2200 4080 2260
rect 4120 2200 4180 2260
rect 4020 2100 4080 2160
rect 4120 2100 4180 2160
rect 1520 1680 1580 1740
rect 1620 1680 1680 1740
rect 1720 1680 1780 1740
rect 1820 1680 1880 1740
rect 1920 1680 1980 1740
rect 2020 1680 2080 1740
rect 2120 1680 2180 1740
rect 2220 1680 2280 1740
rect 2320 1680 2380 1740
rect 2420 1680 2480 1740
rect 2520 1680 2580 1740
rect 2620 1680 2680 1740
rect 2720 1680 2780 1740
rect 2820 1680 2880 1740
rect 2920 1680 2980 1740
rect 3020 1680 3080 1740
rect 3120 1680 3180 1740
rect 3220 1680 3280 1740
rect 3320 1680 3380 1740
rect 3420 1680 3480 1740
rect 3520 1680 3580 1740
rect 3620 1680 3680 1740
rect 3720 1680 3780 1740
rect 3820 1680 3880 1740
rect 3920 1680 3980 1740
rect 4020 1680 4080 1740
rect 4120 1680 4180 1740
rect 4220 1680 4280 1740
rect 4320 1680 4380 1740
rect 4420 1680 4480 1740
rect 4520 1680 4580 1740
rect 4620 1680 4680 1740
rect 4720 1680 4780 1740
rect 4820 1680 4880 1740
rect 4920 1680 4980 1740
rect 5020 1680 5080 1740
rect 5120 1680 5180 1740
rect 5220 1680 5280 1740
rect 5320 1680 5380 1740
rect 5420 1680 5480 1740
rect 5520 1680 5580 1740
rect 5620 1680 5680 1740
rect 5720 1680 5780 1740
rect 5820 1680 5880 1740
rect 5920 1680 5980 1740
rect 6020 1680 6080 1740
rect 6120 1680 6180 1740
rect 6220 1680 6280 1740
rect 6320 1680 6380 1740
rect 6420 1680 6480 1740
rect 6520 1680 6580 1740
rect 6620 1680 6680 1740
rect 1520 1560 1580 1620
rect 1620 1560 1680 1620
rect 1720 1560 1780 1620
rect 1820 1560 1880 1620
rect 1920 1560 1980 1620
rect 2020 1560 2080 1620
rect 2120 1560 2180 1620
rect 2220 1560 2280 1620
rect 2320 1560 2380 1620
rect 2420 1560 2480 1620
rect 2520 1560 2580 1620
rect 2620 1560 2680 1620
rect 2720 1560 2780 1620
rect 2820 1560 2880 1620
rect 2920 1560 2980 1620
rect 3020 1560 3080 1620
rect 3120 1560 3180 1620
rect 3220 1560 3280 1620
rect 3320 1560 3380 1620
rect 3420 1560 3480 1620
rect 3520 1560 3580 1620
rect 3620 1560 3680 1620
rect 3720 1560 3780 1620
rect 3820 1560 3880 1620
rect 3920 1560 3980 1620
rect 4020 1560 4080 1620
rect 4120 1560 4180 1620
rect 4220 1560 4280 1620
rect 4320 1560 4380 1620
rect 4420 1560 4480 1620
rect 4520 1560 4580 1620
rect 4620 1560 4680 1620
rect 4720 1560 4780 1620
rect 4820 1560 4880 1620
rect 4920 1560 4980 1620
rect 5020 1560 5080 1620
rect 5120 1560 5180 1620
rect 5220 1560 5280 1620
rect 5320 1560 5380 1620
rect 5420 1560 5480 1620
rect 5520 1560 5580 1620
rect 5620 1560 5680 1620
rect 5720 1560 5780 1620
rect 5820 1560 5880 1620
rect 5920 1560 5980 1620
rect 6020 1560 6080 1620
rect 6120 1560 6180 1620
rect 6220 1560 6280 1620
rect 6320 1560 6380 1620
rect 6420 1560 6480 1620
rect 6520 1560 6580 1620
rect 6620 1560 6680 1620
rect 4020 1140 4080 1200
rect 4120 1140 4180 1200
rect 4020 1040 4080 1100
rect 4120 1040 4180 1100
rect 4020 940 4080 1000
rect 4120 940 4180 1000
rect 4020 840 4080 900
rect 4120 840 4180 900
rect 4020 740 4080 800
rect 4120 740 4180 800
rect 4020 640 4080 700
rect 4120 640 4180 700
rect 4020 540 4080 600
rect 4120 540 4180 600
rect 4020 440 4080 500
rect 4120 440 4180 500
rect 4020 340 4080 400
rect 4120 340 4180 400
rect 4020 240 4080 300
rect 4120 240 4180 300
rect 4020 140 4080 200
rect 4120 140 4180 200
rect 4020 40 4080 100
rect 4120 40 4180 100
rect 4020 -60 4080 0
rect 4120 -60 4180 0
rect 1320 -280 1380 -220
<< metal1 >>
rect 4000 3380 4200 3400
rect 2020 3360 2280 3380
rect 2020 3300 2040 3360
rect 2100 3300 2200 3360
rect 2260 3300 2280 3360
rect 2020 3260 2280 3300
rect 2020 3200 2040 3260
rect 2100 3200 2200 3260
rect 2260 3200 2280 3260
rect 1800 2880 1980 3140
rect 2020 3060 2280 3200
rect 1800 2820 1820 2880
rect 1880 2820 1980 2880
rect 1800 2780 1980 2820
rect 1800 2720 1820 2780
rect 1880 2720 1980 2780
rect 1800 2100 1980 2720
rect 2320 2880 2500 3140
rect 3000 2900 3180 3140
rect 2320 2820 2420 2880
rect 2480 2820 2500 2880
rect 2320 2780 2500 2820
rect 2320 2720 2420 2780
rect 2480 2720 2500 2780
rect 2320 2100 2500 2720
rect 2980 2700 3180 2900
rect 3000 2500 3180 2700
rect 2980 2480 3180 2500
rect 2980 2420 3000 2480
rect 3060 2420 3180 2480
rect 2980 2380 3180 2420
rect 2980 2320 3000 2380
rect 3060 2320 3180 2380
rect 2980 2300 3180 2320
rect 3000 2100 3180 2300
rect 3520 2480 3700 3140
rect 3520 2420 3620 2480
rect 3680 2420 3700 2480
rect 3520 2380 3700 2420
rect 3520 2320 3620 2380
rect 3680 2320 3700 2380
rect 3240 2140 3460 2160
rect 3220 2000 3480 2140
rect 3520 2100 3700 2320
rect 4000 3080 4020 3380
rect 4080 3080 4120 3380
rect 4180 3080 4200 3380
rect 5920 3360 6180 3380
rect 5920 3300 5940 3360
rect 6000 3300 6100 3360
rect 6160 3300 6180 3360
rect 5920 3260 6180 3300
rect 5920 3200 5940 3260
rect 6000 3200 6100 3260
rect 6160 3200 6180 3260
rect 4000 3060 4200 3080
rect 4000 3000 4020 3060
rect 4080 3000 4120 3060
rect 4180 3000 4200 3060
rect 4000 2980 4200 3000
rect 4000 2680 4020 2980
rect 4080 2680 4120 2980
rect 4180 2680 4200 2980
rect 4000 2660 4200 2680
rect 4000 2600 4020 2660
rect 4080 2600 4120 2660
rect 4180 2600 4200 2660
rect 4000 2580 4200 2600
rect 4000 2280 4020 2580
rect 4080 2280 4120 2580
rect 4180 2280 4200 2580
rect 4500 2500 4680 3140
rect 4480 2480 4680 2500
rect 4480 2420 4500 2480
rect 4560 2420 4680 2480
rect 4480 2380 4680 2420
rect 4480 2320 4500 2380
rect 4560 2320 4680 2380
rect 4480 2300 4680 2320
rect 4000 2260 4200 2280
rect 4000 2200 4020 2260
rect 4080 2200 4120 2260
rect 4180 2200 4200 2260
rect 4000 2180 4200 2200
rect 4000 2100 4020 2180
rect 4080 2100 4120 2180
rect 4180 2100 4200 2180
rect 4500 2100 4680 2300
rect 5020 2500 5180 3140
rect 5700 2900 5880 3160
rect 5920 3060 6180 3200
rect 5680 2880 5880 2900
rect 5680 2820 5700 2880
rect 5760 2820 5880 2880
rect 5680 2780 5880 2820
rect 5680 2720 5700 2780
rect 5760 2720 5880 2780
rect 5680 2700 5880 2720
rect 5020 2480 5200 2500
rect 5020 2420 5120 2480
rect 5180 2420 5200 2480
rect 5020 2380 5200 2420
rect 5020 2320 5120 2380
rect 5180 2320 5200 2380
rect 5020 2300 5200 2320
rect 4000 2080 4200 2100
rect 4720 2000 4980 2160
rect 5020 2100 5180 2300
rect 5700 2100 5880 2700
rect 6220 2880 6400 3160
rect 6220 2820 6320 2880
rect 6380 2820 6400 2880
rect 6220 2780 6400 2820
rect 6220 2720 6320 2780
rect 6380 2720 6400 2780
rect 6220 2100 6400 2720
rect 900 1980 7300 2000
rect 900 1920 1520 1980
rect 1580 1920 1620 1980
rect 1680 1920 6520 1980
rect 6580 1920 6620 1980
rect 6680 1920 7300 1980
rect 900 1880 7300 1920
rect 900 1820 1520 1880
rect 1580 1820 1620 1880
rect 1680 1820 6520 1880
rect 6580 1820 6620 1880
rect 6680 1820 7300 1880
rect 900 1800 7300 1820
rect 1500 1740 6700 1760
rect 1500 1680 1520 1740
rect 1580 1680 1620 1740
rect 1680 1680 1720 1740
rect 1780 1680 1820 1740
rect 1880 1680 1920 1740
rect 1980 1680 2020 1740
rect 2080 1680 2120 1740
rect 2180 1680 2220 1740
rect 2280 1680 2320 1740
rect 2380 1680 2420 1740
rect 2480 1680 2520 1740
rect 2580 1680 2620 1740
rect 2680 1680 2720 1740
rect 2780 1680 2820 1740
rect 2880 1680 2920 1740
rect 2980 1680 3020 1740
rect 3080 1680 3120 1740
rect 3180 1680 3220 1740
rect 3280 1680 3320 1740
rect 3380 1680 3420 1740
rect 3480 1680 3520 1740
rect 3580 1680 3620 1740
rect 3680 1680 3720 1740
rect 3780 1680 3820 1740
rect 3880 1680 3920 1740
rect 3980 1680 4020 1740
rect 4080 1680 4120 1740
rect 4180 1680 4220 1740
rect 4280 1680 4320 1740
rect 4380 1680 4420 1740
rect 4480 1680 4520 1740
rect 4580 1680 4620 1740
rect 4680 1680 4720 1740
rect 4780 1680 4820 1740
rect 4880 1680 4920 1740
rect 4980 1680 5020 1740
rect 5080 1680 5120 1740
rect 5180 1680 5220 1740
rect 5280 1680 5320 1740
rect 5380 1680 5420 1740
rect 5480 1680 5520 1740
rect 5580 1680 5620 1740
rect 5680 1680 5720 1740
rect 5780 1680 5820 1740
rect 5880 1680 5920 1740
rect 5980 1680 6020 1740
rect 6080 1680 6120 1740
rect 6180 1680 6220 1740
rect 6280 1680 6320 1740
rect 6380 1680 6420 1740
rect 6480 1680 6520 1740
rect 6580 1680 6620 1740
rect 6680 1680 6700 1740
rect 1500 1620 6700 1680
rect 1500 1560 1520 1620
rect 1580 1560 1620 1620
rect 1680 1560 1720 1620
rect 1780 1560 1820 1620
rect 1880 1560 1920 1620
rect 1980 1560 2020 1620
rect 2080 1560 2120 1620
rect 2180 1560 2220 1620
rect 2280 1560 2320 1620
rect 2380 1560 2420 1620
rect 2480 1560 2520 1620
rect 2580 1560 2620 1620
rect 2680 1560 2720 1620
rect 2780 1560 2820 1620
rect 2880 1560 2920 1620
rect 2980 1560 3020 1620
rect 3080 1560 3120 1620
rect 3180 1560 3220 1620
rect 3280 1560 3320 1620
rect 3380 1560 3420 1620
rect 3480 1560 3520 1620
rect 3580 1560 3620 1620
rect 3680 1560 3720 1620
rect 3780 1560 3820 1620
rect 3880 1560 3920 1620
rect 3980 1560 4020 1620
rect 4080 1560 4120 1620
rect 4180 1560 4220 1620
rect 4280 1560 4320 1620
rect 4380 1560 4420 1620
rect 4480 1560 4520 1620
rect 4580 1560 4620 1620
rect 4680 1560 4720 1620
rect 4780 1560 4820 1620
rect 4880 1560 4920 1620
rect 4980 1560 5020 1620
rect 5080 1560 5120 1620
rect 5180 1560 5220 1620
rect 5280 1560 5320 1620
rect 5380 1560 5420 1620
rect 5480 1560 5520 1620
rect 5580 1560 5620 1620
rect 5680 1560 5720 1620
rect 5780 1560 5820 1620
rect 5880 1560 5920 1620
rect 5980 1560 6020 1620
rect 6080 1560 6120 1620
rect 6180 1560 6220 1620
rect 6280 1560 6320 1620
rect 6380 1560 6420 1620
rect 6480 1560 6520 1620
rect 6580 1560 6620 1620
rect 6680 1560 6700 1620
rect 1500 1540 6700 1560
rect 900 1480 7300 1500
rect 900 1420 2620 1480
rect 2680 1420 2720 1480
rect 2780 1420 5420 1480
rect 5480 1420 5520 1480
rect 5580 1420 7300 1480
rect 900 1380 7300 1420
rect 900 1320 2620 1380
rect 2680 1320 2720 1380
rect 2780 1320 5420 1380
rect 5480 1320 5520 1380
rect 5580 1320 7300 1380
rect 900 1300 7300 1320
rect 1800 980 1980 1260
rect 1800 920 1820 980
rect 1880 920 1980 980
rect 1800 880 1980 920
rect 1800 820 1820 880
rect 1880 820 1980 880
rect 1800 200 1980 820
rect 2320 980 2500 1260
rect 2320 920 2400 980
rect 2460 920 2500 980
rect 2320 880 2500 920
rect 2320 820 2400 880
rect 2460 820 2500 880
rect 2020 100 2280 240
rect 2320 200 2500 820
rect 3000 580 3180 1260
rect 3220 1160 3480 1300
rect 3000 520 3020 580
rect 3080 520 3180 580
rect 3000 480 3180 520
rect 3000 420 3020 480
rect 3080 420 3180 480
rect 3000 200 3180 420
rect 3520 580 3700 1260
rect 3520 520 3600 580
rect 3660 520 3700 580
rect 3520 480 3700 520
rect 3520 420 3600 480
rect 3660 420 3700 480
rect 3520 200 3700 420
rect 4000 1200 4200 1220
rect 4000 1120 4020 1200
rect 4080 1120 4120 1200
rect 4180 1120 4200 1200
rect 4000 1100 4200 1120
rect 4000 1040 4020 1100
rect 4080 1040 4120 1100
rect 4180 1040 4200 1100
rect 4000 1020 4200 1040
rect 4000 720 4020 1020
rect 4080 720 4120 1020
rect 4180 720 4200 1020
rect 4000 700 4200 720
rect 4000 640 4020 700
rect 4080 640 4120 700
rect 4180 640 4200 700
rect 4000 620 4200 640
rect 4000 320 4020 620
rect 4080 320 4120 620
rect 4180 320 4200 620
rect 4000 300 4200 320
rect 4000 240 4020 300
rect 4080 240 4120 300
rect 4180 240 4200 300
rect 4000 220 4200 240
rect 2020 40 2040 100
rect 2100 40 2200 100
rect 2260 40 2280 100
rect 2020 0 2280 40
rect 2020 -60 2040 0
rect 2100 -60 2200 0
rect 2260 -60 2280 0
rect 2020 -80 2280 -60
rect 4000 -80 4020 220
rect 4080 -80 4120 220
rect 4180 -80 4200 220
rect 4500 580 4680 1260
rect 4720 1160 4980 1300
rect 4500 520 4520 580
rect 4580 520 4680 580
rect 4500 480 4680 520
rect 4500 420 4520 480
rect 4580 420 4680 480
rect 4500 200 4680 420
rect 5020 580 5200 1260
rect 5020 520 5100 580
rect 5160 520 5200 580
rect 5020 480 5200 520
rect 5020 420 5100 480
rect 5160 420 5200 480
rect 5020 200 5200 420
rect 5700 980 5880 1260
rect 5700 920 5720 980
rect 5780 920 5880 980
rect 5700 880 5880 920
rect 5700 820 5720 880
rect 5780 820 5880 880
rect 5700 200 5880 820
rect 6220 980 6400 1260
rect 6220 920 6300 980
rect 6360 920 6400 980
rect 6220 880 6400 920
rect 6220 820 6300 880
rect 6360 820 6400 880
rect 5920 100 6180 260
rect 6220 200 6400 820
rect 5920 40 5940 100
rect 6000 40 6100 100
rect 6160 40 6180 100
rect 5920 0 6180 40
rect 5920 -60 5940 0
rect 6000 -60 6100 0
rect 6160 -60 6180 0
rect 5920 -80 6180 -60
rect 4000 -100 4200 -80
rect 300 -120 500 -100
rect 300 -180 320 -120
rect 380 -180 420 -120
rect 480 -180 500 -120
rect 300 -220 500 -180
rect 300 -280 320 -220
rect 380 -280 420 -220
rect 480 -280 500 -220
rect 300 -300 500 -280
rect 600 -120 800 -100
rect 600 -180 620 -120
rect 680 -180 720 -120
rect 780 -180 800 -120
rect 600 -220 800 -180
rect 7400 -120 7600 -100
rect 7400 -180 7420 -120
rect 7480 -180 7520 -120
rect 7580 -180 7600 -120
rect 600 -280 620 -220
rect 680 -280 720 -220
rect 780 -280 800 -220
rect 600 -300 800 -280
rect 1300 -220 1400 -200
rect 1300 -280 1320 -220
rect 1380 -280 1400 -220
rect 1300 -300 1400 -280
rect 7400 -220 7600 -180
rect 7400 -280 7420 -220
rect 7480 -280 7520 -220
rect 7580 -280 7600 -220
rect 7400 -300 7600 -280
rect 7700 -120 7900 -100
rect 7700 -180 7720 -120
rect 7780 -180 7820 -120
rect 7880 -180 7900 -120
rect 7700 -220 7900 -180
rect 7700 -280 7720 -220
rect 7780 -280 7820 -220
rect 7880 -280 7900 -220
rect 7700 -300 7900 -280
rect 4000 -320 4200 -300
rect 4000 -380 4020 -320
rect 4080 -380 4120 -320
rect 4180 -380 4200 -320
rect 4000 -420 4200 -380
rect 4000 -480 4020 -420
rect 4080 -480 4120 -420
rect 4180 -480 4200 -420
rect 4000 -500 4200 -480
<< via1 >>
rect 2040 3300 2100 3360
rect 2200 3300 2260 3360
rect 2040 3200 2100 3260
rect 2200 3200 2260 3260
rect 1820 2820 1880 2880
rect 1820 2720 1880 2780
rect 2420 2820 2480 2880
rect 2420 2720 2480 2780
rect 3000 2420 3060 2480
rect 3000 2320 3060 2380
rect 3620 2420 3680 2480
rect 3620 2320 3680 2380
rect 4020 3360 4080 3380
rect 4020 3320 4080 3360
rect 4020 3260 4080 3300
rect 4020 3240 4080 3260
rect 4020 3200 4080 3220
rect 4020 3160 4080 3200
rect 4020 3100 4080 3140
rect 4020 3080 4080 3100
rect 4120 3360 4180 3380
rect 4120 3320 4180 3360
rect 4120 3260 4180 3300
rect 4120 3240 4180 3260
rect 4120 3200 4180 3220
rect 4120 3160 4180 3200
rect 4120 3100 4180 3140
rect 4120 3080 4180 3100
rect 5940 3300 6000 3360
rect 6100 3300 6160 3360
rect 5940 3200 6000 3260
rect 6100 3200 6160 3260
rect 4020 3000 4080 3060
rect 4120 3000 4180 3060
rect 4020 2960 4080 2980
rect 4020 2920 4080 2960
rect 4020 2860 4080 2900
rect 4020 2840 4080 2860
rect 4020 2800 4080 2820
rect 4020 2760 4080 2800
rect 4020 2700 4080 2740
rect 4020 2680 4080 2700
rect 4120 2960 4180 2980
rect 4120 2920 4180 2960
rect 4120 2860 4180 2900
rect 4120 2840 4180 2860
rect 4120 2800 4180 2820
rect 4120 2760 4180 2800
rect 4120 2700 4180 2740
rect 4120 2680 4180 2700
rect 4020 2600 4080 2660
rect 4120 2600 4180 2660
rect 4020 2560 4080 2580
rect 4020 2520 4080 2560
rect 4020 2460 4080 2500
rect 4020 2440 4080 2460
rect 4020 2400 4080 2420
rect 4020 2360 4080 2400
rect 4020 2300 4080 2340
rect 4020 2280 4080 2300
rect 4120 2560 4180 2580
rect 4120 2520 4180 2560
rect 4120 2460 4180 2500
rect 4120 2440 4180 2460
rect 4120 2400 4180 2420
rect 4120 2360 4180 2400
rect 4120 2300 4180 2340
rect 4120 2280 4180 2300
rect 4500 2420 4560 2480
rect 4500 2320 4560 2380
rect 4020 2200 4080 2260
rect 4120 2200 4180 2260
rect 4020 2160 4080 2180
rect 4020 2120 4080 2160
rect 4120 2160 4180 2180
rect 4120 2120 4180 2160
rect 5700 2820 5760 2880
rect 5700 2720 5760 2780
rect 5120 2420 5180 2480
rect 5120 2320 5180 2380
rect 6320 2820 6380 2880
rect 6320 2720 6380 2780
rect 1520 1920 1580 1980
rect 1620 1920 1680 1980
rect 6520 1920 6580 1980
rect 6620 1920 6680 1980
rect 1520 1820 1580 1880
rect 1620 1820 1680 1880
rect 6520 1820 6580 1880
rect 6620 1820 6680 1880
rect 4020 1680 4080 1740
rect 4120 1680 4180 1740
rect 4020 1560 4080 1620
rect 4120 1560 4180 1620
rect 2620 1420 2680 1480
rect 2720 1420 2780 1480
rect 5420 1420 5480 1480
rect 5520 1420 5580 1480
rect 2620 1320 2680 1380
rect 2720 1320 2780 1380
rect 5420 1320 5480 1380
rect 5520 1320 5580 1380
rect 1820 920 1880 980
rect 1820 820 1880 880
rect 2400 920 2460 980
rect 2400 820 2460 880
rect 3020 520 3080 580
rect 3020 420 3080 480
rect 3600 520 3660 580
rect 3600 420 3660 480
rect 4020 1140 4080 1180
rect 4020 1120 4080 1140
rect 4120 1140 4180 1180
rect 4120 1120 4180 1140
rect 4020 1040 4080 1100
rect 4120 1040 4180 1100
rect 4020 1000 4080 1020
rect 4020 960 4080 1000
rect 4020 900 4080 940
rect 4020 880 4080 900
rect 4020 840 4080 860
rect 4020 800 4080 840
rect 4020 740 4080 780
rect 4020 720 4080 740
rect 4120 1000 4180 1020
rect 4120 960 4180 1000
rect 4120 900 4180 940
rect 4120 880 4180 900
rect 4120 840 4180 860
rect 4120 800 4180 840
rect 4120 740 4180 780
rect 4120 720 4180 740
rect 4020 640 4080 700
rect 4120 640 4180 700
rect 4020 600 4080 620
rect 4020 560 4080 600
rect 4020 500 4080 540
rect 4020 480 4080 500
rect 4020 440 4080 460
rect 4020 400 4080 440
rect 4020 340 4080 380
rect 4020 320 4080 340
rect 4120 600 4180 620
rect 4120 560 4180 600
rect 4120 500 4180 540
rect 4120 480 4180 500
rect 4120 440 4180 460
rect 4120 400 4180 440
rect 4120 340 4180 380
rect 4120 320 4180 340
rect 4020 240 4080 300
rect 4120 240 4180 300
rect 2040 40 2100 100
rect 2200 40 2260 100
rect 2040 -60 2100 0
rect 2200 -60 2260 0
rect 4020 200 4080 220
rect 4020 160 4080 200
rect 4020 100 4080 140
rect 4020 80 4080 100
rect 4020 40 4080 60
rect 4020 0 4080 40
rect 4020 -60 4080 -20
rect 4020 -80 4080 -60
rect 4120 200 4180 220
rect 4120 160 4180 200
rect 4120 100 4180 140
rect 4120 80 4180 100
rect 4120 40 4180 60
rect 4120 0 4180 40
rect 4120 -60 4180 -20
rect 4120 -80 4180 -60
rect 4520 520 4580 580
rect 4520 420 4580 480
rect 5100 520 5160 580
rect 5100 420 5160 480
rect 5720 920 5780 980
rect 5720 820 5780 880
rect 6300 920 6360 980
rect 6300 820 6360 880
rect 5940 40 6000 100
rect 6100 40 6160 100
rect 5940 -60 6000 0
rect 6100 -60 6160 0
rect 320 -180 380 -120
rect 420 -180 480 -120
rect 320 -280 380 -220
rect 420 -280 480 -220
rect 620 -180 680 -120
rect 720 -180 780 -120
rect 7420 -180 7480 -120
rect 7520 -180 7580 -120
rect 620 -280 680 -220
rect 720 -280 780 -220
rect 7420 -280 7480 -220
rect 7520 -280 7580 -220
rect 7720 -180 7780 -120
rect 7820 -180 7880 -120
rect 7720 -280 7780 -220
rect 7820 -280 7880 -220
rect 4020 -380 4080 -320
rect 4120 -380 4180 -320
rect 4020 -480 4080 -420
rect 4120 -480 4180 -420
<< metal2 >>
rect 300 2480 500 3600
rect 300 2420 320 2480
rect 380 2420 420 2480
rect 480 2420 500 2480
rect 300 2380 500 2420
rect 300 2320 320 2380
rect 380 2320 420 2380
rect 480 2320 500 2380
rect 300 980 500 2320
rect 300 920 320 980
rect 380 920 420 980
rect 480 920 500 980
rect 300 880 500 920
rect 300 820 320 880
rect 380 820 420 880
rect 480 820 500 880
rect 300 -120 500 820
rect 300 -180 320 -120
rect 380 -180 420 -120
rect 480 -180 500 -120
rect 300 -220 500 -180
rect 300 -280 320 -220
rect 380 -280 420 -220
rect 480 -280 500 -220
rect 300 -300 500 -280
rect 600 2880 800 3600
rect 4000 3380 4200 3400
rect 2000 3360 2800 3380
rect 2000 3300 2040 3360
rect 2100 3300 2200 3360
rect 2260 3300 2800 3360
rect 2000 3260 2800 3300
rect 2000 3200 2040 3260
rect 2100 3200 2200 3260
rect 2260 3200 2800 3260
rect 2000 3180 2800 3200
rect 600 2820 620 2880
rect 680 2820 720 2880
rect 780 2820 800 2880
rect 600 2780 800 2820
rect 600 2720 620 2780
rect 680 2720 720 2780
rect 780 2720 800 2780
rect 600 580 800 2720
rect 1800 2880 1900 2900
rect 1800 2820 1820 2880
rect 1880 2820 1900 2880
rect 1800 2780 1900 2820
rect 1800 2720 1820 2780
rect 1880 2720 1900 2780
rect 1800 2700 1900 2720
rect 2400 2880 2500 2900
rect 2400 2820 2420 2880
rect 2480 2820 2500 2880
rect 2400 2780 2500 2820
rect 2400 2720 2420 2780
rect 2480 2720 2500 2780
rect 2400 2700 2500 2720
rect 600 520 620 580
rect 680 520 720 580
rect 780 520 800 580
rect 600 480 800 520
rect 600 420 620 480
rect 680 420 720 480
rect 780 420 800 480
rect 600 -120 800 420
rect 1500 1980 1700 2000
rect 1500 1920 1520 1980
rect 1580 1920 1620 1980
rect 1680 1920 1700 1980
rect 1500 1880 1700 1920
rect 1500 1820 1520 1880
rect 1580 1820 1620 1880
rect 1680 1820 1700 1880
rect 1500 120 1700 1820
rect 2600 1480 2800 3180
rect 4000 3320 4020 3380
rect 4080 3320 4120 3380
rect 4180 3320 4200 3380
rect 4000 3300 4200 3320
rect 4000 3240 4020 3300
rect 4080 3240 4120 3300
rect 4180 3240 4200 3300
rect 4000 3220 4200 3240
rect 4000 3160 4020 3220
rect 4080 3160 4120 3220
rect 4180 3160 4200 3220
rect 4000 3140 4200 3160
rect 4000 3080 4020 3140
rect 4080 3080 4120 3140
rect 4180 3080 4200 3140
rect 4000 3060 4200 3080
rect 4000 3000 4020 3060
rect 4080 3000 4120 3060
rect 4180 3000 4200 3060
rect 4000 2980 4200 3000
rect 4000 2920 4020 2980
rect 4080 2920 4120 2980
rect 4180 2920 4200 2980
rect 4000 2900 4200 2920
rect 4000 2840 4020 2900
rect 4080 2840 4120 2900
rect 4180 2840 4200 2900
rect 4000 2820 4200 2840
rect 4000 2760 4020 2820
rect 4080 2760 4120 2820
rect 4180 2760 4200 2820
rect 4000 2740 4200 2760
rect 4000 2680 4020 2740
rect 4080 2680 4120 2740
rect 4180 2680 4200 2740
rect 4000 2660 4200 2680
rect 4000 2600 4020 2660
rect 4080 2600 4120 2660
rect 4180 2600 4200 2660
rect 4000 2580 4200 2600
rect 4000 2520 4020 2580
rect 4080 2520 4120 2580
rect 4180 2520 4200 2580
rect 4000 2500 4200 2520
rect 5400 3360 6200 3380
rect 5400 3300 5940 3360
rect 6000 3300 6100 3360
rect 6160 3300 6200 3360
rect 5400 3260 6200 3300
rect 5400 3200 5940 3260
rect 6000 3200 6100 3260
rect 6160 3200 6200 3260
rect 5400 3180 6200 3200
rect 2980 2480 3080 2500
rect 2980 2420 3000 2480
rect 3060 2420 3080 2480
rect 2980 2380 3080 2420
rect 2980 2320 3000 2380
rect 3060 2320 3080 2380
rect 2980 2300 3080 2320
rect 3600 2480 3700 2500
rect 3600 2420 3620 2480
rect 3680 2420 3700 2480
rect 3600 2380 3700 2420
rect 3600 2320 3620 2380
rect 3680 2320 3700 2380
rect 3600 2300 3700 2320
rect 4000 2440 4020 2500
rect 4080 2440 4120 2500
rect 4180 2440 4200 2500
rect 4000 2420 4200 2440
rect 4000 2360 4020 2420
rect 4080 2360 4120 2420
rect 4180 2360 4200 2420
rect 4000 2340 4200 2360
rect 2600 1420 2620 1480
rect 2680 1420 2720 1480
rect 2780 1420 2800 1480
rect 2600 1380 2800 1420
rect 2600 1320 2620 1380
rect 2680 1320 2720 1380
rect 2780 1320 2800 1380
rect 2600 1300 2800 1320
rect 4000 2280 4020 2340
rect 4080 2280 4120 2340
rect 4180 2280 4200 2340
rect 4480 2480 4580 2500
rect 4480 2420 4500 2480
rect 4560 2420 4580 2480
rect 4480 2380 4580 2420
rect 4480 2320 4500 2380
rect 4560 2320 4580 2380
rect 4480 2300 4580 2320
rect 5100 2480 5200 2500
rect 5100 2420 5120 2480
rect 5180 2420 5200 2480
rect 5100 2380 5200 2420
rect 5100 2320 5120 2380
rect 5180 2320 5200 2380
rect 5100 2300 5200 2320
rect 4000 2260 4200 2280
rect 4000 2200 4020 2260
rect 4080 2200 4120 2260
rect 4180 2200 4200 2260
rect 4000 2180 4200 2200
rect 4000 2120 4020 2180
rect 4080 2120 4120 2180
rect 4180 2120 4200 2180
rect 4000 1740 4200 2120
rect 4000 1680 4020 1740
rect 4080 1680 4120 1740
rect 4180 1680 4200 1740
rect 4000 1620 4200 1680
rect 4000 1560 4020 1620
rect 4080 1560 4120 1620
rect 4180 1560 4200 1620
rect 4000 1180 4200 1560
rect 5400 1480 5600 3180
rect 5680 2880 5780 2900
rect 5680 2820 5700 2880
rect 5760 2820 5780 2880
rect 5680 2780 5780 2820
rect 5680 2720 5700 2780
rect 5760 2720 5780 2780
rect 5680 2700 5780 2720
rect 6300 2880 6400 2900
rect 6300 2820 6320 2880
rect 6380 2820 6400 2880
rect 6300 2780 6400 2820
rect 6300 2720 6320 2780
rect 6380 2720 6400 2780
rect 6300 2700 6400 2720
rect 7400 2880 7600 3600
rect 7400 2820 7420 2880
rect 7480 2820 7520 2880
rect 7580 2820 7600 2880
rect 7400 2780 7600 2820
rect 7400 2720 7420 2780
rect 7480 2720 7520 2780
rect 7580 2720 7600 2780
rect 5400 1420 5420 1480
rect 5480 1420 5520 1480
rect 5580 1420 5600 1480
rect 5400 1380 5600 1420
rect 5400 1320 5420 1380
rect 5480 1320 5520 1380
rect 5580 1320 5600 1380
rect 5400 1300 5600 1320
rect 6500 1980 6700 2000
rect 6500 1920 6520 1980
rect 6580 1920 6620 1980
rect 6680 1920 6700 1980
rect 6500 1880 6700 1920
rect 6500 1820 6520 1880
rect 6580 1820 6620 1880
rect 6680 1820 6700 1880
rect 4000 1120 4020 1180
rect 4080 1120 4120 1180
rect 4180 1120 4200 1180
rect 4000 1100 4200 1120
rect 4000 1040 4020 1100
rect 4080 1040 4120 1100
rect 4180 1040 4200 1100
rect 4000 1020 4200 1040
rect 1800 980 1900 1000
rect 1800 920 1820 980
rect 1880 920 1900 980
rect 1800 880 1900 920
rect 1800 820 1820 880
rect 1880 820 1900 880
rect 1800 800 1900 820
rect 2380 980 2480 1000
rect 2380 920 2400 980
rect 2460 920 2480 980
rect 2380 880 2480 920
rect 2380 820 2400 880
rect 2460 820 2480 880
rect 2380 800 2480 820
rect 4000 960 4020 1020
rect 4080 960 4120 1020
rect 4180 960 4200 1020
rect 4000 940 4200 960
rect 4000 880 4020 940
rect 4080 880 4120 940
rect 4180 880 4200 940
rect 4000 860 4200 880
rect 4000 800 4020 860
rect 4080 800 4120 860
rect 4180 800 4200 860
rect 5700 980 5800 1000
rect 5700 920 5720 980
rect 5780 920 5800 980
rect 5700 880 5800 920
rect 5700 820 5720 880
rect 5780 820 5800 880
rect 5700 800 5800 820
rect 6280 980 6380 1000
rect 6280 920 6300 980
rect 6360 920 6380 980
rect 6280 880 6380 920
rect 6280 820 6300 880
rect 6360 820 6380 880
rect 6280 800 6380 820
rect 4000 780 4200 800
rect 4000 720 4020 780
rect 4080 720 4120 780
rect 4180 720 4200 780
rect 4000 700 4200 720
rect 4000 640 4020 700
rect 4080 640 4120 700
rect 4180 640 4200 700
rect 4000 620 4200 640
rect 3000 580 3100 600
rect 3000 520 3020 580
rect 3080 520 3100 580
rect 3000 480 3100 520
rect 3000 420 3020 480
rect 3080 420 3100 480
rect 3000 400 3100 420
rect 3580 580 3680 600
rect 3580 520 3600 580
rect 3660 520 3680 580
rect 3580 480 3680 520
rect 3580 420 3600 480
rect 3660 420 3680 480
rect 3580 400 3680 420
rect 4000 560 4020 620
rect 4080 560 4120 620
rect 4180 560 4200 620
rect 4000 540 4200 560
rect 4000 480 4020 540
rect 4080 480 4120 540
rect 4180 480 4200 540
rect 4000 460 4200 480
rect 4000 400 4020 460
rect 4080 400 4120 460
rect 4180 400 4200 460
rect 4500 580 4600 600
rect 4500 520 4520 580
rect 4580 520 4600 580
rect 4500 480 4600 520
rect 4500 420 4520 480
rect 4580 420 4600 480
rect 4500 400 4600 420
rect 5080 580 5180 600
rect 5080 520 5100 580
rect 5160 520 5180 580
rect 5080 480 5180 520
rect 5080 420 5100 480
rect 5160 420 5180 480
rect 5080 400 5180 420
rect 4000 380 4200 400
rect 4000 320 4020 380
rect 4080 320 4120 380
rect 4180 320 4200 380
rect 4000 300 4200 320
rect 4000 240 4020 300
rect 4080 240 4120 300
rect 4180 240 4200 300
rect 4000 220 4200 240
rect 4000 160 4020 220
rect 4080 160 4120 220
rect 4180 160 4200 220
rect 4000 140 4200 160
rect 1500 100 2300 120
rect 1500 40 2040 100
rect 2100 40 2200 100
rect 2260 40 2300 100
rect 1500 0 2300 40
rect 1500 -60 2040 0
rect 2100 -60 2200 0
rect 2260 -60 2300 0
rect 1500 -80 2300 -60
rect 4000 80 4020 140
rect 4080 80 4120 140
rect 4180 80 4200 140
rect 6500 120 6700 1820
rect 4000 60 4200 80
rect 4000 0 4020 60
rect 4080 0 4120 60
rect 4180 0 4200 60
rect 4000 -20 4200 0
rect 4000 -80 4020 -20
rect 4080 -80 4120 -20
rect 4180 -80 4200 -20
rect 5900 100 6700 120
rect 5900 40 5940 100
rect 6000 40 6100 100
rect 6160 40 6700 100
rect 5900 0 6700 40
rect 5900 -60 5940 0
rect 6000 -60 6100 0
rect 6160 -60 6700 0
rect 5900 -80 6700 -60
rect 7400 580 7600 2720
rect 7400 520 7420 580
rect 7480 520 7520 580
rect 7580 520 7600 580
rect 7400 480 7600 520
rect 7400 420 7420 480
rect 7480 420 7520 480
rect 7580 420 7600 480
rect 600 -180 620 -120
rect 680 -180 720 -120
rect 780 -180 800 -120
rect 600 -220 800 -180
rect 600 -280 620 -220
rect 680 -280 720 -220
rect 780 -280 800 -220
rect 600 -300 800 -280
rect 4000 -320 4200 -80
rect 7400 -120 7600 420
rect 7400 -180 7420 -120
rect 7480 -180 7520 -120
rect 7580 -180 7600 -120
rect 7400 -220 7600 -180
rect 7400 -280 7420 -220
rect 7480 -280 7520 -220
rect 7580 -280 7600 -220
rect 7400 -300 7600 -280
rect 7700 2480 7900 3600
rect 7700 2420 7720 2480
rect 7780 2420 7820 2480
rect 7880 2420 7900 2480
rect 7700 2380 7900 2420
rect 7700 2320 7720 2380
rect 7780 2320 7820 2380
rect 7880 2320 7900 2380
rect 7700 980 7900 2320
rect 7700 920 7720 980
rect 7780 920 7820 980
rect 7880 920 7900 980
rect 7700 880 7900 920
rect 7700 820 7720 880
rect 7780 820 7820 880
rect 7880 820 7900 880
rect 7700 -120 7900 820
rect 7700 -180 7720 -120
rect 7780 -180 7820 -120
rect 7880 -180 7900 -120
rect 7700 -220 7900 -180
rect 7700 -280 7720 -220
rect 7780 -280 7820 -220
rect 7880 -280 7900 -220
rect 7700 -300 7900 -280
rect 4000 -380 4020 -320
rect 4080 -380 4120 -320
rect 4180 -380 4200 -320
rect 4000 -420 4200 -380
rect 4000 -480 4020 -420
rect 4080 -480 4120 -420
rect 4180 -480 4200 -420
rect 4000 -500 4200 -480
<< via2 >>
rect 320 2420 380 2480
rect 420 2420 480 2480
rect 320 2320 380 2380
rect 420 2320 480 2380
rect 320 920 380 980
rect 420 920 480 980
rect 320 820 380 880
rect 420 820 480 880
rect 620 2820 680 2880
rect 720 2820 780 2880
rect 620 2720 680 2780
rect 720 2720 780 2780
rect 1820 2820 1880 2880
rect 1820 2720 1880 2780
rect 2420 2820 2480 2880
rect 2420 2720 2480 2780
rect 620 520 680 580
rect 720 520 780 580
rect 620 420 680 480
rect 720 420 780 480
rect 3000 2420 3060 2480
rect 3000 2320 3060 2380
rect 3620 2420 3680 2480
rect 3620 2320 3680 2380
rect 4500 2420 4560 2480
rect 4500 2320 4560 2380
rect 5120 2420 5180 2480
rect 5120 2320 5180 2380
rect 5700 2820 5760 2880
rect 5700 2720 5760 2780
rect 6320 2820 6380 2880
rect 6320 2720 6380 2780
rect 7420 2820 7480 2880
rect 7520 2820 7580 2880
rect 7420 2720 7480 2780
rect 7520 2720 7580 2780
rect 1820 920 1880 980
rect 1820 820 1880 880
rect 2400 920 2460 980
rect 2400 820 2460 880
rect 5720 920 5780 980
rect 5720 820 5780 880
rect 6300 920 6360 980
rect 6300 820 6360 880
rect 3020 520 3080 580
rect 3020 420 3080 480
rect 3600 520 3660 580
rect 3600 420 3660 480
rect 4520 520 4580 580
rect 4520 420 4580 480
rect 5100 520 5160 580
rect 5100 420 5160 480
rect 7420 520 7480 580
rect 7520 520 7580 580
rect 7420 420 7480 480
rect 7520 420 7580 480
rect 7720 2420 7780 2480
rect 7820 2420 7880 2480
rect 7720 2320 7780 2380
rect 7820 2320 7880 2380
rect 7720 920 7780 980
rect 7820 920 7880 980
rect 7720 820 7780 880
rect 7820 820 7880 880
<< metal3 >>
rect 300 2880 7900 2900
rect 300 2820 620 2880
rect 680 2820 720 2880
rect 780 2820 1820 2880
rect 1880 2820 2420 2880
rect 2480 2820 5700 2880
rect 5760 2820 6320 2880
rect 6380 2820 7420 2880
rect 7480 2820 7520 2880
rect 7580 2820 7900 2880
rect 300 2780 7900 2820
rect 300 2720 620 2780
rect 680 2720 720 2780
rect 780 2720 1820 2780
rect 1880 2720 2420 2780
rect 2480 2720 5700 2780
rect 5760 2720 6320 2780
rect 6380 2720 7420 2780
rect 7480 2720 7520 2780
rect 7580 2720 7900 2780
rect 300 2700 7900 2720
rect 300 2480 7900 2500
rect 300 2420 320 2480
rect 380 2420 420 2480
rect 480 2420 3000 2480
rect 3060 2420 3620 2480
rect 3680 2420 4500 2480
rect 4560 2420 5120 2480
rect 5180 2420 7720 2480
rect 7780 2420 7820 2480
rect 7880 2420 7900 2480
rect 300 2380 7900 2420
rect 300 2320 320 2380
rect 380 2320 420 2380
rect 480 2320 3000 2380
rect 3060 2320 3620 2380
rect 3680 2320 4500 2380
rect 4560 2320 5120 2380
rect 5180 2320 7720 2380
rect 7780 2320 7820 2380
rect 7880 2320 7900 2380
rect 300 2300 7900 2320
rect 300 980 7900 1000
rect 300 920 320 980
rect 380 920 420 980
rect 480 920 1820 980
rect 1880 920 2400 980
rect 2460 920 5720 980
rect 5780 920 6300 980
rect 6360 920 7720 980
rect 7780 920 7820 980
rect 7880 920 7900 980
rect 300 880 7900 920
rect 300 820 320 880
rect 380 820 420 880
rect 480 820 1820 880
rect 1880 820 2400 880
rect 2460 820 5720 880
rect 5780 820 6300 880
rect 6360 820 7720 880
rect 7780 820 7820 880
rect 7880 820 7900 880
rect 300 800 7900 820
rect 300 580 7900 600
rect 300 520 620 580
rect 680 520 720 580
rect 780 520 3020 580
rect 3080 520 3600 580
rect 3660 520 4520 580
rect 4580 520 5100 580
rect 5160 520 7420 580
rect 7480 520 7520 580
rect 7580 520 7900 580
rect 300 480 7900 520
rect 300 420 620 480
rect 680 420 720 480
rect 780 420 3020 480
rect 3080 420 3600 480
rect 3660 420 4520 480
rect 4580 420 5100 480
rect 5160 420 7420 480
rect 7480 420 7520 480
rect 7580 420 7900 480
rect 300 400 7900 420
use sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH  sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_0
timestamp 1769952370
transform 1 0 3345 0 1 2632
box -345 -532 345 532
use sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH  sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_1
timestamp 1769952370
transform 1 0 6045 0 1 732
box -345 -532 345 532
use sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH  sky130_fd_pr__nfet_g5v0d10v5_CQ6KSH_2
timestamp 1769952370
transform 1 0 2145 0 1 732
box -345 -532 345 532
use sky130_fd_pr__nfet_g5v0d10v5_SNDLS5  sky130_fd_pr__nfet_g5v0d10v5_SNDLS5_0
timestamp 1769952370
transform 1 0 4845 0 1 2632
box -345 -532 345 532
use sky130_fd_pr__nfet_g5v0d10v5_X57ESK  sky130_fd_pr__nfet_g5v0d10v5_X57ESK_0
timestamp 1769952370
transform 1 0 2145 0 1 2632
box -345 -532 345 532
use sky130_fd_pr__nfet_g5v0d10v5_X57ESK  sky130_fd_pr__nfet_g5v0d10v5_X57ESK_1
timestamp 1769952370
transform 1 0 6045 0 1 2632
box -345 -532 345 532
use sky130_fd_pr__nfet_g5v0d10v5_X57ESK  sky130_fd_pr__nfet_g5v0d10v5_X57ESK_2
timestamp 1769952370
transform 1 0 4845 0 1 732
box -345 -532 345 532
use sky130_fd_pr__nfet_g5v0d10v5_X57ESK  sky130_fd_pr__nfet_g5v0d10v5_X57ESK_3
timestamp 1769952370
transform 1 0 3345 0 1 732
box -345 -532 345 532
<< labels >>
flabel metal1 900 1300 1100 1500 0 FreeSans 256 0 0 0 VP
port 0 nsew
flabel metal1 900 1800 1100 2000 0 FreeSans 256 0 0 0 VN
port 1 nsew
flabel metal1 640 -300 740 -200 0 FreeSans 256 0 0 0 D1
port 4 nsew
flabel metal1 320 -300 420 -200 0 FreeSans 256 0 0 0 D2
port 3 nsew
flabel metal1 4060 -460 4160 -360 0 FreeSans 256 0 0 0 S
port 2 nsew
flabel metal1 1300 -300 1400 -200 0 FreeSans 256 0 0 0 VSS
port 5 nsew
<< end >>
