magic
tech sky130A
magscale 1 2
timestamp 1768989049
<< nwell >>
rect -705 -797 705 797
<< mvpmos >>
rect -447 -500 -267 500
rect -209 -500 -29 500
rect 29 -500 209 500
rect 267 -500 447 500
<< mvpdiff >>
rect -505 488 -447 500
rect -505 -488 -493 488
rect -459 -488 -447 488
rect -505 -500 -447 -488
rect -267 488 -209 500
rect -267 -488 -255 488
rect -221 -488 -209 488
rect -267 -500 -209 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 209 488 267 500
rect 209 -488 221 488
rect 255 -488 267 488
rect 209 -500 267 -488
rect 447 488 505 500
rect 447 -488 459 488
rect 493 -488 505 488
rect 447 -500 505 -488
<< mvpdiffc >>
rect -493 -488 -459 488
rect -255 -488 -221 488
rect -17 -488 17 488
rect 221 -488 255 488
rect 459 -488 493 488
<< mvnsubdiff >>
rect -639 719 639 731
rect -639 685 -531 719
rect 531 685 639 719
rect -639 673 639 685
rect -639 623 -581 673
rect -639 -623 -627 623
rect -593 -623 -581 623
rect 581 623 639 673
rect -639 -673 -581 -623
rect 581 -623 593 623
rect 627 -623 639 623
rect 581 -673 639 -623
rect -639 -685 639 -673
rect -639 -719 -531 -685
rect 531 -719 639 -685
rect -639 -731 639 -719
<< mvnsubdiffcont >>
rect -531 685 531 719
rect -627 -623 -593 623
rect 593 -623 627 623
rect -531 -719 531 -685
<< poly >>
rect -447 581 -267 597
rect -447 547 -431 581
rect -283 547 -267 581
rect -447 500 -267 547
rect -209 581 -29 597
rect -209 547 -193 581
rect -45 547 -29 581
rect -209 500 -29 547
rect 29 581 209 597
rect 29 547 45 581
rect 193 547 209 581
rect 29 500 209 547
rect 267 581 447 597
rect 267 547 283 581
rect 431 547 447 581
rect 267 500 447 547
rect -447 -547 -267 -500
rect -447 -581 -431 -547
rect -283 -581 -267 -547
rect -447 -597 -267 -581
rect -209 -547 -29 -500
rect -209 -581 -193 -547
rect -45 -581 -29 -547
rect -209 -597 -29 -581
rect 29 -547 209 -500
rect 29 -581 45 -547
rect 193 -581 209 -547
rect 29 -597 209 -581
rect 267 -547 447 -500
rect 267 -581 283 -547
rect 431 -581 447 -547
rect 267 -597 447 -581
<< polycont >>
rect -431 547 -283 581
rect -193 547 -45 581
rect 45 547 193 581
rect 283 547 431 581
rect -431 -581 -283 -547
rect -193 -581 -45 -547
rect 45 -581 193 -547
rect 283 -581 431 -547
<< locali >>
rect -627 685 -531 719
rect 531 685 627 719
rect -627 623 -593 685
rect 593 623 627 685
rect -447 547 -431 581
rect -283 547 -267 581
rect -209 547 -193 581
rect -45 547 -29 581
rect 29 547 45 581
rect 193 547 209 581
rect 267 547 283 581
rect 431 547 447 581
rect -493 488 -459 504
rect -493 -504 -459 -488
rect -255 488 -221 504
rect -255 -504 -221 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 221 488 255 504
rect 221 -504 255 -488
rect 459 488 493 504
rect 459 -504 493 -488
rect -447 -581 -431 -547
rect -283 -581 -267 -547
rect -209 -581 -193 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 193 -581 209 -547
rect 267 -581 283 -547
rect 431 -581 447 -547
rect -627 -685 -593 -623
rect 593 -685 627 -623
rect -627 -719 -531 -685
rect 531 -719 627 -685
<< viali >>
rect -431 547 -283 581
rect -193 547 -45 581
rect 45 547 193 581
rect 283 547 431 581
rect -493 -488 -459 488
rect -255 -488 -221 488
rect -17 -488 17 488
rect 221 -488 255 488
rect 459 -488 493 488
rect -431 -581 -283 -547
rect -193 -581 -45 -547
rect 45 -581 193 -547
rect 283 -581 431 -547
<< metal1 >>
rect -443 581 -271 587
rect -443 547 -431 581
rect -283 547 -271 581
rect -443 541 -271 547
rect -205 581 -33 587
rect -205 547 -193 581
rect -45 547 -33 581
rect -205 541 -33 547
rect 33 581 205 587
rect 33 547 45 581
rect 193 547 205 581
rect 33 541 205 547
rect 271 581 443 587
rect 271 547 283 581
rect 431 547 443 581
rect 271 541 443 547
rect -499 488 -453 500
rect -499 -488 -493 488
rect -459 -488 -453 488
rect -499 -500 -453 -488
rect -261 488 -215 500
rect -261 -488 -255 488
rect -221 -488 -215 488
rect -261 -500 -215 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 215 488 261 500
rect 215 -488 221 488
rect 255 -488 261 488
rect 215 -500 261 -488
rect 453 488 499 500
rect 453 -488 459 488
rect 493 -488 499 488
rect 453 -500 499 -488
rect -443 -547 -271 -541
rect -443 -581 -431 -547
rect -283 -581 -271 -547
rect -443 -587 -271 -581
rect -205 -547 -33 -541
rect -205 -581 -193 -547
rect -45 -581 -33 -547
rect -205 -587 -33 -581
rect 33 -547 205 -541
rect 33 -581 45 -547
rect 193 -581 205 -547
rect 33 -587 205 -581
rect 271 -547 443 -541
rect 271 -581 283 -547
rect 431 -581 443 -547
rect 271 -587 443 -581
<< properties >>
string FIXED_BBOX -610 -702 610 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.9 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
