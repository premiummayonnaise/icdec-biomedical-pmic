magic
tech sky130A
magscale 1 2
timestamp 1768759310
<< error_p >>
rect -891 341 891 345
rect -891 -273 -861 341
rect -825 275 -459 279
rect -397 275 -31 279
rect 31 275 397 279
rect 459 275 825 279
rect -825 -207 -795 275
rect 795 -207 825 275
rect 861 -273 891 341
<< nwell >>
rect -861 -307 861 341
<< mvpmos >>
rect -767 -207 -517 279
rect -339 -207 -89 279
rect 89 -207 339 279
rect 517 -207 767 279
<< mvpdiff >>
rect -825 267 -767 279
rect -825 -195 -813 267
rect -779 -195 -767 267
rect -825 -207 -767 -195
rect -517 267 -459 279
rect -517 -195 -505 267
rect -471 -195 -459 267
rect -517 -207 -459 -195
rect -397 267 -339 279
rect -397 -195 -385 267
rect -351 -195 -339 267
rect -397 -207 -339 -195
rect -89 267 -31 279
rect -89 -195 -77 267
rect -43 -195 -31 267
rect -89 -207 -31 -195
rect 31 267 89 279
rect 31 -195 43 267
rect 77 -195 89 267
rect 31 -207 89 -195
rect 339 267 397 279
rect 339 -195 351 267
rect 385 -195 397 267
rect 339 -207 397 -195
rect 459 267 517 279
rect 459 -195 471 267
rect 505 -195 517 267
rect 459 -207 517 -195
rect 767 267 825 279
rect 767 -195 779 267
rect 813 -195 825 267
rect 767 -207 825 -195
<< mvpdiffc >>
rect -813 -195 -779 267
rect -505 -195 -471 267
rect -385 -195 -351 267
rect -77 -195 -43 267
rect 43 -195 77 267
rect 351 -195 385 267
rect 471 -195 505 267
rect 779 -195 813 267
<< poly >>
rect -767 279 -517 305
rect -339 279 -89 305
rect 89 279 339 305
rect 517 279 767 305
rect -767 -254 -517 -207
rect -767 -288 -751 -254
rect -533 -288 -517 -254
rect -767 -304 -517 -288
rect -339 -254 -89 -207
rect -339 -288 -323 -254
rect -105 -288 -89 -254
rect -339 -304 -89 -288
rect 89 -254 339 -207
rect 89 -288 105 -254
rect 323 -288 339 -254
rect 89 -304 339 -288
rect 517 -254 767 -207
rect 517 -288 533 -254
rect 751 -288 767 -254
rect 517 -304 767 -288
<< polycont >>
rect -751 -288 -533 -254
rect -323 -288 -105 -254
rect 105 -288 323 -254
rect 533 -288 751 -254
<< locali >>
rect -813 267 -779 283
rect -813 -211 -779 -195
rect -505 267 -471 283
rect -505 -211 -471 -195
rect -385 267 -351 283
rect -385 -211 -351 -195
rect -77 267 -43 283
rect -77 -211 -43 -195
rect 43 267 77 283
rect 43 -211 77 -195
rect 351 267 385 283
rect 351 -211 385 -195
rect 471 267 505 283
rect 471 -211 505 -195
rect 779 267 813 283
rect 779 -211 813 -195
rect -767 -288 -751 -254
rect -533 -288 -517 -254
rect -339 -288 -323 -254
rect -105 -288 -89 -254
rect 89 -288 105 -254
rect 323 -288 339 -254
rect 517 -288 533 -254
rect 751 -288 767 -254
<< viali >>
rect -813 -195 -779 267
rect -505 -195 -471 267
rect -385 -195 -351 267
rect -77 -195 -43 267
rect 43 -195 77 267
rect 351 -195 385 267
rect 471 -195 505 267
rect 779 -195 813 267
rect -751 -288 -533 -254
rect -323 -288 -105 -254
rect 105 -288 323 -254
rect 533 -288 751 -254
<< metal1 >>
rect -819 267 -773 279
rect -819 -195 -813 267
rect -779 -195 -773 267
rect -819 -207 -773 -195
rect -511 267 -465 279
rect -511 -195 -505 267
rect -471 -195 -465 267
rect -511 -207 -465 -195
rect -391 267 -345 279
rect -391 -195 -385 267
rect -351 -195 -345 267
rect -391 -207 -345 -195
rect -83 267 -37 279
rect -83 -195 -77 267
rect -43 -195 -37 267
rect -83 -207 -37 -195
rect 37 267 83 279
rect 37 -195 43 267
rect 77 -195 83 267
rect 37 -207 83 -195
rect 345 267 391 279
rect 345 -195 351 267
rect 385 -195 391 267
rect 345 -207 391 -195
rect 465 267 511 279
rect 465 -195 471 267
rect 505 -195 511 267
rect 465 -207 511 -195
rect 773 267 819 279
rect 773 -195 779 267
rect 813 -195 819 267
rect 773 -207 819 -195
rect -763 -254 -521 -248
rect -763 -288 -751 -254
rect -533 -288 -521 -254
rect -763 -294 -521 -288
rect -335 -254 -93 -248
rect -335 -288 -323 -254
rect -105 -288 -93 -254
rect -335 -294 -93 -288
rect 93 -254 335 -248
rect 93 -288 105 -254
rect 323 -288 335 -254
rect 93 -294 335 -288
rect 521 -254 763 -248
rect 521 -288 533 -254
rect 751 -288 763 -254
rect 521 -294 763 -288
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.425 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
