magic
tech sky130A
magscale 1 2
timestamp 1769135993
<< nmos >>
rect -458 -139 -358 201
rect -186 -139 -86 201
rect 86 -139 186 201
rect 358 -139 458 201
<< ndiff >>
rect -516 189 -458 201
rect -516 -127 -504 189
rect -470 -127 -458 189
rect -516 -139 -458 -127
rect -358 189 -300 201
rect -358 -127 -346 189
rect -312 -127 -300 189
rect -358 -139 -300 -127
rect -244 189 -186 201
rect -244 -127 -232 189
rect -198 -127 -186 189
rect -244 -139 -186 -127
rect -86 189 -28 201
rect -86 -127 -74 189
rect -40 -127 -28 189
rect -86 -139 -28 -127
rect 28 189 86 201
rect 28 -127 40 189
rect 74 -127 86 189
rect 28 -139 86 -127
rect 186 189 244 201
rect 186 -127 198 189
rect 232 -127 244 189
rect 186 -139 244 -127
rect 300 189 358 201
rect 300 -127 312 189
rect 346 -127 358 189
rect 300 -139 358 -127
rect 458 189 516 201
rect 458 -127 470 189
rect 504 -127 516 189
rect 458 -139 516 -127
<< ndiffc >>
rect -504 -127 -470 189
rect -346 -127 -312 189
rect -232 -127 -198 189
rect -74 -127 -40 189
rect 40 -127 74 189
rect 198 -127 232 189
rect 312 -127 346 189
rect 470 -127 504 189
<< poly >>
rect -458 201 -358 227
rect -186 201 -86 227
rect 86 201 186 227
rect 358 201 458 227
rect -458 -177 -358 -139
rect -458 -211 -442 -177
rect -374 -211 -358 -177
rect -458 -227 -358 -211
rect -186 -177 -86 -139
rect -186 -211 -170 -177
rect -102 -211 -86 -177
rect -186 -227 -86 -211
rect 86 -177 186 -139
rect 86 -211 102 -177
rect 170 -211 186 -177
rect 86 -227 186 -211
rect 358 -177 458 -139
rect 358 -211 374 -177
rect 442 -211 458 -177
rect 358 -227 458 -211
<< polycont >>
rect -442 -211 -374 -177
rect -170 -211 -102 -177
rect 102 -211 170 -177
rect 374 -211 442 -177
<< locali >>
rect -504 189 -470 205
rect -504 -143 -470 -127
rect -346 189 -312 205
rect -346 -143 -312 -127
rect -232 189 -198 205
rect -232 -143 -198 -127
rect -74 189 -40 205
rect -74 -143 -40 -127
rect 40 189 74 205
rect 40 -143 74 -127
rect 198 189 232 205
rect 198 -143 232 -127
rect 312 189 346 205
rect 312 -143 346 -127
rect 470 189 504 205
rect 470 -143 504 -127
rect -458 -211 -442 -177
rect -374 -211 -358 -177
rect -186 -211 -170 -177
rect -102 -211 -86 -177
rect 86 -211 102 -177
rect 170 -211 186 -177
rect 358 -211 374 -177
rect 442 -211 458 -177
<< viali >>
rect -504 -127 -470 189
rect -346 -127 -312 189
rect -232 -127 -198 189
rect -74 -127 -40 189
rect 40 -127 74 189
rect 198 -127 232 189
rect 312 -127 346 189
rect 470 -127 504 189
rect -442 -211 -374 -177
rect -170 -211 -102 -177
rect 102 -211 170 -177
rect 374 -211 442 -177
<< metal1 >>
rect -510 189 -464 201
rect -510 -127 -504 189
rect -470 -127 -464 189
rect -510 -139 -464 -127
rect -352 189 -306 201
rect -352 -127 -346 189
rect -312 -127 -306 189
rect -352 -139 -306 -127
rect -238 189 -192 201
rect -238 -127 -232 189
rect -198 -127 -192 189
rect -238 -139 -192 -127
rect -80 189 -34 201
rect -80 -127 -74 189
rect -40 -127 -34 189
rect -80 -139 -34 -127
rect 34 189 80 201
rect 34 -127 40 189
rect 74 -127 80 189
rect 34 -139 80 -127
rect 192 189 238 201
rect 192 -127 198 189
rect 232 -127 238 189
rect 192 -139 238 -127
rect 306 189 352 201
rect 306 -127 312 189
rect 346 -127 352 189
rect 306 -139 352 -127
rect 464 189 510 201
rect 464 -127 470 189
rect 504 -127 510 189
rect 464 -139 510 -127
rect -454 -177 -362 -171
rect -454 -211 -442 -177
rect -374 -211 -362 -177
rect -454 -217 -362 -211
rect -182 -177 -90 -171
rect -182 -211 -170 -177
rect -102 -211 -90 -177
rect -182 -217 -90 -211
rect 90 -177 182 -171
rect 90 -211 102 -177
rect 170 -211 182 -177
rect 90 -217 182 -211
rect 362 -177 454 -171
rect 362 -211 374 -177
rect 442 -211 454 -177
rect 362 -217 454 -211
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.7 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
