magic
tech sky130A
magscale 1 2
timestamp 1769076474
<< nwell >>
rect -437 -601 437 601
<< mvpmos >>
rect -179 -375 -29 375
rect 29 -375 179 375
<< mvpdiff >>
rect -237 363 -179 375
rect -237 -363 -225 363
rect -191 -363 -179 363
rect -237 -375 -179 -363
rect -29 363 29 375
rect -29 -363 -17 363
rect 17 -363 29 363
rect -29 -375 29 -363
rect 179 363 237 375
rect 179 -363 191 363
rect 225 -363 237 363
rect 179 -375 237 -363
<< mvpdiffc >>
rect -225 -363 -191 363
rect -17 -363 17 363
rect 191 -363 225 363
<< mvnsubdiff >>
rect -371 523 371 535
rect -371 489 -263 523
rect 263 489 371 523
rect -371 477 371 489
rect -371 427 -313 477
rect -371 -427 -359 427
rect -325 -427 -313 427
rect 313 427 371 477
rect -371 -477 -313 -427
rect 313 -427 325 427
rect 359 -427 371 427
rect 313 -477 371 -427
rect -371 -489 371 -477
rect -371 -523 -263 -489
rect 263 -523 371 -489
rect -371 -535 371 -523
<< mvnsubdiffcont >>
rect -263 489 263 523
rect -359 -427 -325 427
rect 325 -427 359 427
rect -263 -523 263 -489
<< poly >>
rect -179 375 -29 401
rect 29 375 179 401
rect -179 -401 -29 -375
rect 29 -401 179 -375
<< locali >>
rect -359 489 -263 523
rect 263 489 359 523
rect -359 427 -325 489
rect 325 427 359 489
rect -225 363 -191 379
rect -225 -379 -191 -363
rect -17 363 17 379
rect -17 -379 17 -363
rect 191 363 225 379
rect 191 -379 225 -363
rect -359 -489 -325 -427
rect 325 -489 359 -427
rect -359 -523 -263 -489
rect 263 -523 359 -489
<< viali >>
rect -225 -363 -191 363
rect -17 -363 17 363
rect 191 -363 225 363
<< metal1 >>
rect -231 363 -185 375
rect -231 -363 -225 363
rect -191 -363 -185 363
rect -231 -375 -185 -363
rect -23 363 23 375
rect -23 -363 -17 363
rect 17 -363 23 363
rect -23 -375 23 -363
rect 185 363 231 375
rect 185 -363 191 363
rect 225 -363 231 363
rect 185 -375 231 -363
<< properties >>
string FIXED_BBOX -342 -506 342 506
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3.75 l 0.75 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
