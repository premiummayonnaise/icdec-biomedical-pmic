magic
tech sky130A
magscale 1 2
timestamp 1769529800
<< pwell >>
rect -815 -1008 815 1008
<< mvnmos >>
rect -587 -750 -337 750
rect -279 -750 -29 750
rect 29 -750 279 750
rect 337 -750 587 750
<< mvndiff >>
rect -645 738 -587 750
rect -645 -738 -633 738
rect -599 -738 -587 738
rect -645 -750 -587 -738
rect -337 738 -279 750
rect -337 -738 -325 738
rect -291 -738 -279 738
rect -337 -750 -279 -738
rect -29 738 29 750
rect -29 -738 -17 738
rect 17 -738 29 738
rect -29 -750 29 -738
rect 279 738 337 750
rect 279 -738 291 738
rect 325 -738 337 738
rect 279 -750 337 -738
rect 587 738 645 750
rect 587 -738 599 738
rect 633 -738 645 738
rect 587 -750 645 -738
<< mvndiffc >>
rect -633 -738 -599 738
rect -325 -738 -291 738
rect -17 -738 17 738
rect 291 -738 325 738
rect 599 -738 633 738
<< mvpsubdiff >>
rect -779 960 779 972
rect -779 926 -671 960
rect 671 926 779 960
rect -779 914 779 926
rect -779 864 -721 914
rect -779 -864 -767 864
rect -733 -864 -721 864
rect 721 864 779 914
rect -779 -914 -721 -864
rect 721 -864 733 864
rect 767 -864 779 864
rect 721 -914 779 -864
rect -779 -926 779 -914
rect -779 -960 -671 -926
rect 671 -960 779 -926
rect -779 -972 779 -960
<< mvpsubdiffcont >>
rect -671 926 671 960
rect -767 -864 -733 864
rect 733 -864 767 864
rect -671 -960 671 -926
<< poly >>
rect -587 822 -337 838
rect -587 788 -571 822
rect -353 788 -337 822
rect -587 750 -337 788
rect -279 822 -29 838
rect -279 788 -263 822
rect -45 788 -29 822
rect -279 750 -29 788
rect 29 822 279 838
rect 29 788 45 822
rect 263 788 279 822
rect 29 750 279 788
rect 337 822 587 838
rect 337 788 353 822
rect 571 788 587 822
rect 337 750 587 788
rect -587 -788 -337 -750
rect -587 -822 -571 -788
rect -353 -822 -337 -788
rect -587 -838 -337 -822
rect -279 -788 -29 -750
rect -279 -822 -263 -788
rect -45 -822 -29 -788
rect -279 -838 -29 -822
rect 29 -788 279 -750
rect 29 -822 45 -788
rect 263 -822 279 -788
rect 29 -838 279 -822
rect 337 -788 587 -750
rect 337 -822 353 -788
rect 571 -822 587 -788
rect 337 -838 587 -822
<< polycont >>
rect -571 788 -353 822
rect -263 788 -45 822
rect 45 788 263 822
rect 353 788 571 822
rect -571 -822 -353 -788
rect -263 -822 -45 -788
rect 45 -822 263 -788
rect 353 -822 571 -788
<< locali >>
rect -767 926 -671 960
rect 671 926 767 960
rect -767 864 -733 926
rect 733 864 767 926
rect -587 788 -571 822
rect -353 788 -337 822
rect -279 788 -263 822
rect -45 788 -29 822
rect 29 788 45 822
rect 263 788 279 822
rect 337 788 353 822
rect 571 788 587 822
rect -633 738 -599 754
rect -633 -754 -599 -738
rect -325 738 -291 754
rect -325 -754 -291 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 291 738 325 754
rect 291 -754 325 -738
rect 599 738 633 754
rect 599 -754 633 -738
rect -587 -822 -571 -788
rect -353 -822 -337 -788
rect -279 -822 -263 -788
rect -45 -822 -29 -788
rect 29 -822 45 -788
rect 263 -822 279 -788
rect 337 -822 353 -788
rect 571 -822 587 -788
rect -767 -926 -733 -864
rect 733 -926 767 -864
rect -767 -960 -671 -926
rect 671 -960 767 -926
<< viali >>
rect -571 788 -353 822
rect -263 788 -45 822
rect 45 788 263 822
rect 353 788 571 822
rect -633 -738 -599 738
rect -325 -738 -291 738
rect -17 -738 17 738
rect 291 -738 325 738
rect 599 -738 633 738
rect -571 -822 -353 -788
rect -263 -822 -45 -788
rect 45 -822 263 -788
rect 353 -822 571 -788
<< metal1 >>
rect -583 822 -341 828
rect -583 788 -571 822
rect -353 788 -341 822
rect -583 782 -341 788
rect -275 822 -33 828
rect -275 788 -263 822
rect -45 788 -33 822
rect -275 782 -33 788
rect 33 822 275 828
rect 33 788 45 822
rect 263 788 275 822
rect 33 782 275 788
rect 341 822 583 828
rect 341 788 353 822
rect 571 788 583 822
rect 341 782 583 788
rect -639 738 -593 750
rect -639 -738 -633 738
rect -599 -738 -593 738
rect -639 -750 -593 -738
rect -331 738 -285 750
rect -331 -738 -325 738
rect -291 -738 -285 738
rect -331 -750 -285 -738
rect -23 738 23 750
rect -23 -738 -17 738
rect 17 -738 23 738
rect -23 -750 23 -738
rect 285 738 331 750
rect 285 -738 291 738
rect 325 -738 331 738
rect 285 -750 331 -738
rect 593 738 639 750
rect 593 -738 599 738
rect 633 -738 639 738
rect 593 -750 639 -738
rect -583 -788 -341 -782
rect -583 -822 -571 -788
rect -353 -822 -341 -788
rect -583 -828 -341 -822
rect -275 -788 -33 -782
rect -275 -822 -263 -788
rect -45 -822 -33 -788
rect -275 -828 -33 -822
rect 33 -788 275 -782
rect 33 -822 45 -788
rect 263 -822 275 -788
rect 33 -828 275 -822
rect 341 -788 583 -782
rect 341 -822 353 -788
rect 571 -822 583 -788
rect 341 -828 583 -822
<< properties >>
string FIXED_BBOX -750 -943 750 943
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
