magic
tech sky130A
magscale 1 2
timestamp 1769417084
<< error_p >>
rect -571 598 571 602
rect -571 -530 -541 598
rect -505 532 505 536
rect -505 -464 -475 532
rect 475 -464 505 532
rect 541 -530 571 598
<< nwell >>
rect -541 -564 541 598
<< mvpmos >>
rect -447 -464 -267 536
rect -209 -464 -29 536
rect 29 -464 209 536
rect 267 -464 447 536
<< mvpdiff >>
rect -505 524 -447 536
rect -505 -452 -493 524
rect -459 -452 -447 524
rect -505 -464 -447 -452
rect -267 524 -209 536
rect -267 -452 -255 524
rect -221 -452 -209 524
rect -267 -464 -209 -452
rect -29 524 29 536
rect -29 -452 -17 524
rect 17 -452 29 524
rect -29 -464 29 -452
rect 209 524 267 536
rect 209 -452 221 524
rect 255 -452 267 524
rect 209 -464 267 -452
rect 447 524 505 536
rect 447 -452 459 524
rect 493 -452 505 524
rect 447 -464 505 -452
<< mvpdiffc >>
rect -493 -452 -459 524
rect -255 -452 -221 524
rect -17 -452 17 524
rect 221 -452 255 524
rect 459 -452 493 524
<< poly >>
rect -447 536 -267 562
rect -209 536 -29 562
rect 29 536 209 562
rect 267 536 447 562
rect -447 -511 -267 -464
rect -447 -545 -431 -511
rect -283 -545 -267 -511
rect -447 -561 -267 -545
rect -209 -511 -29 -464
rect -209 -545 -193 -511
rect -45 -545 -29 -511
rect -209 -561 -29 -545
rect 29 -511 209 -464
rect 29 -545 45 -511
rect 193 -545 209 -511
rect 29 -561 209 -545
rect 267 -511 447 -464
rect 267 -545 283 -511
rect 431 -545 447 -511
rect 267 -561 447 -545
<< polycont >>
rect -431 -545 -283 -511
rect -193 -545 -45 -511
rect 45 -545 193 -511
rect 283 -545 431 -511
<< locali >>
rect -493 524 -459 540
rect -493 -468 -459 -452
rect -255 524 -221 540
rect -255 -468 -221 -452
rect -17 524 17 540
rect -17 -468 17 -452
rect 221 524 255 540
rect 221 -468 255 -452
rect 459 524 493 540
rect 459 -468 493 -452
rect -447 -545 -431 -511
rect -283 -545 -267 -511
rect -209 -545 -193 -511
rect -45 -545 -29 -511
rect 29 -545 45 -511
rect 193 -545 209 -511
rect 267 -545 283 -511
rect 431 -545 447 -511
<< viali >>
rect -493 -452 -459 524
rect -255 -452 -221 524
rect -17 -452 17 524
rect 221 -452 255 524
rect 459 -452 493 524
rect -431 -545 -283 -511
rect -193 -545 -45 -511
rect 45 -545 193 -511
rect 283 -545 431 -511
<< metal1 >>
rect -499 524 -453 536
rect -499 -452 -493 524
rect -459 -452 -453 524
rect -499 -464 -453 -452
rect -261 524 -215 536
rect -261 -452 -255 524
rect -221 -452 -215 524
rect -261 -464 -215 -452
rect -23 524 23 536
rect -23 -452 -17 524
rect 17 -452 23 524
rect -23 -464 23 -452
rect 215 524 261 536
rect 215 -452 221 524
rect 255 -452 261 524
rect 215 -464 261 -452
rect 453 524 499 536
rect 453 -452 459 524
rect 493 -452 499 524
rect 453 -464 499 -452
rect -443 -511 -271 -505
rect -443 -545 -431 -511
rect -283 -545 -271 -511
rect -443 -551 -271 -545
rect -205 -511 -33 -505
rect -205 -545 -193 -511
rect -45 -545 -33 -511
rect -205 -551 -33 -545
rect 33 -511 205 -505
rect 33 -545 45 -511
rect 193 -545 205 -511
rect 33 -551 205 -545
rect 271 -511 443 -505
rect 271 -545 283 -511
rect 431 -545 443 -511
rect 271 -551 443 -545
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.9 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
