magic
tech sky130A
magscale 1 2
timestamp 1768989364
<< nwell >>
rect -645 -672 645 672
<< mvpmos >>
rect -387 -375 -237 375
rect -179 -375 -29 375
rect 29 -375 179 375
rect 237 -375 387 375
<< mvpdiff >>
rect -445 363 -387 375
rect -445 -363 -433 363
rect -399 -363 -387 363
rect -445 -375 -387 -363
rect -237 363 -179 375
rect -237 -363 -225 363
rect -191 -363 -179 363
rect -237 -375 -179 -363
rect -29 363 29 375
rect -29 -363 -17 363
rect 17 -363 29 363
rect -29 -375 29 -363
rect 179 363 237 375
rect 179 -363 191 363
rect 225 -363 237 363
rect 179 -375 237 -363
rect 387 363 445 375
rect 387 -363 399 363
rect 433 -363 445 363
rect 387 -375 445 -363
<< mvpdiffc >>
rect -433 -363 -399 363
rect -225 -363 -191 363
rect -17 -363 17 363
rect 191 -363 225 363
rect 399 -363 433 363
<< mvnsubdiff >>
rect -579 594 579 606
rect -579 560 -471 594
rect 471 560 579 594
rect -579 548 579 560
rect -579 498 -521 548
rect -579 -498 -567 498
rect -533 -498 -521 498
rect 521 498 579 548
rect -579 -548 -521 -498
rect 521 -498 533 498
rect 567 -498 579 498
rect 521 -548 579 -498
rect -579 -560 579 -548
rect -579 -594 -471 -560
rect 471 -594 579 -560
rect -579 -606 579 -594
<< mvnsubdiffcont >>
rect -471 560 471 594
rect -567 -498 -533 498
rect 533 -498 567 498
rect -471 -594 471 -560
<< poly >>
rect -387 456 -237 472
rect -387 422 -371 456
rect -253 422 -237 456
rect -387 375 -237 422
rect -179 456 -29 472
rect -179 422 -163 456
rect -45 422 -29 456
rect -179 375 -29 422
rect 29 456 179 472
rect 29 422 45 456
rect 163 422 179 456
rect 29 375 179 422
rect 237 456 387 472
rect 237 422 253 456
rect 371 422 387 456
rect 237 375 387 422
rect -387 -422 -237 -375
rect -387 -456 -371 -422
rect -253 -456 -237 -422
rect -387 -472 -237 -456
rect -179 -422 -29 -375
rect -179 -456 -163 -422
rect -45 -456 -29 -422
rect -179 -472 -29 -456
rect 29 -422 179 -375
rect 29 -456 45 -422
rect 163 -456 179 -422
rect 29 -472 179 -456
rect 237 -422 387 -375
rect 237 -456 253 -422
rect 371 -456 387 -422
rect 237 -472 387 -456
<< polycont >>
rect -371 422 -253 456
rect -163 422 -45 456
rect 45 422 163 456
rect 253 422 371 456
rect -371 -456 -253 -422
rect -163 -456 -45 -422
rect 45 -456 163 -422
rect 253 -456 371 -422
<< locali >>
rect -567 560 -471 594
rect 471 560 567 594
rect -567 498 -533 560
rect 533 498 567 560
rect -387 422 -371 456
rect -253 422 -237 456
rect -179 422 -163 456
rect -45 422 -29 456
rect 29 422 45 456
rect 163 422 179 456
rect 237 422 253 456
rect 371 422 387 456
rect -433 363 -399 379
rect -433 -379 -399 -363
rect -225 363 -191 379
rect -225 -379 -191 -363
rect -17 363 17 379
rect -17 -379 17 -363
rect 191 363 225 379
rect 191 -379 225 -363
rect 399 363 433 379
rect 399 -379 433 -363
rect -387 -456 -371 -422
rect -253 -456 -237 -422
rect -179 -456 -163 -422
rect -45 -456 -29 -422
rect 29 -456 45 -422
rect 163 -456 179 -422
rect 237 -456 253 -422
rect 371 -456 387 -422
rect -567 -560 -533 -498
rect 533 -560 567 -498
rect -567 -594 -471 -560
rect 471 -594 567 -560
<< viali >>
rect -371 422 -253 456
rect -163 422 -45 456
rect 45 422 163 456
rect 253 422 371 456
rect -433 -363 -399 363
rect -225 -363 -191 363
rect -17 -363 17 363
rect 191 -363 225 363
rect 399 -363 433 363
rect -371 -456 -253 -422
rect -163 -456 -45 -422
rect 45 -456 163 -422
rect 253 -456 371 -422
<< metal1 >>
rect -383 456 -241 462
rect -383 422 -371 456
rect -253 422 -241 456
rect -383 416 -241 422
rect -175 456 -33 462
rect -175 422 -163 456
rect -45 422 -33 456
rect -175 416 -33 422
rect 33 456 175 462
rect 33 422 45 456
rect 163 422 175 456
rect 33 416 175 422
rect 241 456 383 462
rect 241 422 253 456
rect 371 422 383 456
rect 241 416 383 422
rect -439 363 -393 375
rect -439 -363 -433 363
rect -399 -363 -393 363
rect -439 -375 -393 -363
rect -231 363 -185 375
rect -231 -363 -225 363
rect -191 -363 -185 363
rect -231 -375 -185 -363
rect -23 363 23 375
rect -23 -363 -17 363
rect 17 -363 23 363
rect -23 -375 23 -363
rect 185 363 231 375
rect 185 -363 191 363
rect 225 -363 231 363
rect 185 -375 231 -363
rect 393 363 439 375
rect 393 -363 399 363
rect 433 -363 439 363
rect 393 -375 439 -363
rect -383 -422 -241 -416
rect -383 -456 -371 -422
rect -253 -456 -241 -422
rect -383 -462 -241 -456
rect -175 -422 -33 -416
rect -175 -456 -163 -422
rect -45 -456 -33 -422
rect -175 -462 -33 -456
rect 33 -422 175 -416
rect 33 -456 45 -422
rect 163 -456 175 -422
rect 33 -462 175 -456
rect 241 -422 383 -416
rect 241 -456 253 -422
rect 371 -456 383 -422
rect 241 -462 383 -456
<< labels >>
rlabel mvnsubdiffcont 0 -577 0 -577 0 B
port 1 nsew
rlabel mvpdiffc -416 0 -416 0 0 D0
port 2 nsew
rlabel polycont -312 439 -312 439 0 G0
port 3 nsew
rlabel mvpdiffc -208 0 -208 0 0 S1
port 4 nsew
rlabel polycont -104 439 -104 439 0 G1
port 5 nsew
rlabel mvpdiffc 0 0 0 0 0 D2
port 6 nsew
rlabel polycont 104 439 104 439 0 G2
port 7 nsew
rlabel mvpdiffc 208 0 208 0 0 S3
port 8 nsew
rlabel polycont 312 439 312 439 0 G3
port 9 nsew
<< properties >>
string FIXED_BBOX -550 -577 550 577
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3.75 l 0.75 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
