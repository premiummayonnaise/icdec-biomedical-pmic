magic
tech sky130A
magscale 1 2
timestamp 1768761814
<< nwell >>
rect 1200 -500 5000 1000
<< pwell >>
rect 1200 -3400 5000 -500
<< psubdiff >>
rect 2300 -550 3960 -540
rect 2300 -590 2360 -550
rect 2480 -590 2520 -550
rect 2640 -590 2680 -550
rect 2800 -590 2840 -550
rect 2960 -590 3000 -550
rect 3120 -590 3160 -550
rect 3260 -590 3300 -550
rect 3420 -590 3460 -550
rect 3580 -590 3620 -550
rect 3740 -590 3780 -550
rect 3900 -590 3960 -550
rect 2300 -600 3960 -590
rect 2300 -1340 2360 -600
rect 3900 -1340 3960 -600
rect 2300 -1350 3960 -1340
rect 2300 -1390 2310 -1350
rect 2430 -1390 3830 -1350
rect 3950 -1390 3960 -1350
rect 2300 -1400 3960 -1390
rect 2300 -2160 2360 -1400
rect 3900 -2160 3960 -1400
rect 2300 -2220 3960 -2160
rect 2520 -2860 2580 -2220
rect 3660 -2860 3720 -2220
rect 2520 -2870 3720 -2860
rect 2520 -2910 2580 -2870
rect 2660 -2910 2700 -2870
rect 2780 -2910 2820 -2870
rect 2900 -2910 2940 -2870
rect 3020 -2910 3060 -2870
rect 3140 -2910 3180 -2870
rect 3260 -2910 3300 -2870
rect 3380 -2910 3420 -2870
rect 3540 -2910 3580 -2870
rect 3660 -2910 3720 -2870
rect 2520 -2920 3720 -2910
<< nsubdiff >>
rect 2100 380 4160 440
rect 2100 -360 2160 380
rect 4100 -360 4160 380
rect 2100 -420 4160 -360
<< psubdiffcont >>
rect 2360 -590 2480 -550
rect 2520 -590 2640 -550
rect 2680 -590 2800 -550
rect 2840 -590 2960 -550
rect 3000 -590 3120 -550
rect 3160 -590 3260 -550
rect 3300 -590 3420 -550
rect 3460 -590 3580 -550
rect 3620 -590 3740 -550
rect 3780 -590 3900 -550
rect 2310 -1390 2430 -1350
rect 3830 -1390 3950 -1350
rect 2580 -2910 2660 -2870
rect 2700 -2910 2780 -2870
rect 2820 -2910 2900 -2870
rect 2940 -2910 3020 -2870
rect 3060 -2910 3140 -2870
rect 3180 -2910 3260 -2870
rect 3300 -2910 3380 -2870
rect 3420 -2910 3540 -2870
rect 3580 -2910 3660 -2870
<< locali >>
rect 1200 400 5000 1000
rect 2100 380 4160 400
rect 2100 -360 2160 380
rect 4100 -360 4160 380
rect 2100 -420 4160 -360
rect 2300 -550 3960 -540
rect 2300 -590 2360 -550
rect 2480 -590 2520 -550
rect 2640 -590 2680 -550
rect 2800 -590 2840 -550
rect 2960 -590 3000 -550
rect 3120 -590 3160 -550
rect 3260 -590 3300 -550
rect 3420 -590 3460 -550
rect 3580 -590 3620 -550
rect 3740 -590 3780 -550
rect 3900 -590 3960 -550
rect 2300 -600 3960 -590
rect 2300 -1340 2360 -600
rect 3900 -1340 3960 -600
rect 2300 -1350 3960 -1340
rect 2300 -1390 2310 -1350
rect 2430 -1390 3830 -1350
rect 3950 -1390 3960 -1350
rect 2300 -1400 3960 -1390
rect 2300 -2160 2360 -1400
rect 3900 -2160 3960 -1400
rect 2300 -2220 3960 -2160
rect 2520 -2800 2580 -2220
rect 3660 -2800 3720 -2220
rect 1200 -2870 5000 -2800
rect 1200 -2910 2580 -2870
rect 2660 -2910 2700 -2870
rect 2780 -2910 2820 -2870
rect 2900 -2910 2940 -2870
rect 3020 -2910 3060 -2870
rect 3140 -2910 3180 -2870
rect 3260 -2910 3300 -2870
rect 3380 -2910 3420 -2870
rect 3540 -2910 3580 -2870
rect 3660 -2910 5000 -2870
rect 1200 -3400 5000 -2910
<< metal1 >>
rect 1201 10397 3201 10398
rect 1201 1000 5006 10397
rect 1200 400 5006 1000
rect 1201 398 5006 400
rect 3006 397 5006 398
rect 1500 -1340 4000 -1240
rect 4500 -1400 4600 -1300
rect 1500 -1500 4000 -1400
rect 1500 -2300 4000 -2200
rect 1200 -3400 5000 -2800
use sky130_fd_pr__nfet_g5v0d10v5_NDYTJY  sky130_fd_pr__nfet_g5v0d10v5_NDYTJY_0
timestamp 1768760819
transform 1 0 3125 0 1 -1830
box -625 -270 625 270
use sky130_fd_pr__nfet_g5v0d10v5_64ZTJY  XM2
timestamp 1768760819
transform 1 0 3125 0 1 -930
box -625 -270 625 270
use sky130_fd_pr__nfet_g5v0d10v5_TNU6Q5  XM3
timestamp 1768760819
transform 1 0 3117 0 1 -2545
box -397 -215 397 215
use sky130_fd_pr__pfet_g5v0d10v5_HRLS9E  XM5
timestamp 1768759310
transform 1 0 3126 0 1 2
box -891 -307 891 345
<< labels >>
flabel metal1 1900 500 2100 700 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1900 -3100 2100 -2900 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 4500 -1400 4600 -1300 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 1500 -1340 1600 -1240 0 FreeSans 256 0 0 0 VN
port 3 nsew
flabel metal1 1500 -1500 1600 -1400 0 FreeSans 256 0 0 0 VP
port 4 nsew
flabel metal1 1500 -2300 1600 -2200 0 FreeSans 256 0 0 0 IBIAS
port 2 nsew
<< end >>
