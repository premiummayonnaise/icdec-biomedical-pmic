magic
tech sky130A
magscale 1 2
timestamp 1769616064
<< error_p >>
rect -521 -220 -463 -214
rect -193 -220 -135 -214
rect 135 -220 193 -214
rect 463 -220 521 -214
rect -521 -254 -509 -220
rect -193 -254 -181 -220
rect 135 -254 147 -220
rect 463 -254 475 -220
rect -521 -260 -463 -254
rect -193 -260 -135 -254
rect 135 -260 193 -254
rect 463 -260 521 -254
<< pwell >>
rect -795 -440 795 440
<< mvnmos >>
rect -567 -182 -417 244
rect -239 -182 -89 244
rect 89 -182 239 244
rect 417 -182 567 244
<< mvndiff >>
rect -625 232 -567 244
rect -625 -170 -613 232
rect -579 -170 -567 232
rect -625 -182 -567 -170
rect -417 232 -359 244
rect -417 -170 -405 232
rect -371 -170 -359 232
rect -417 -182 -359 -170
rect -297 232 -239 244
rect -297 -170 -285 232
rect -251 -170 -239 232
rect -297 -182 -239 -170
rect -89 232 -31 244
rect -89 -170 -77 232
rect -43 -170 -31 232
rect -89 -182 -31 -170
rect 31 232 89 244
rect 31 -170 43 232
rect 77 -170 89 232
rect 31 -182 89 -170
rect 239 232 297 244
rect 239 -170 251 232
rect 285 -170 297 232
rect 239 -182 297 -170
rect 359 232 417 244
rect 359 -170 371 232
rect 405 -170 417 232
rect 359 -182 417 -170
rect 567 232 625 244
rect 567 -170 579 232
rect 613 -170 625 232
rect 567 -182 625 -170
<< mvndiffc >>
rect -613 -170 -579 232
rect -405 -170 -371 232
rect -285 -170 -251 232
rect -77 -170 -43 232
rect 43 -170 77 232
rect 251 -170 285 232
rect 371 -170 405 232
rect 579 -170 613 232
<< mvpsubdiff >>
rect -759 346 759 404
rect -759 296 -701 346
rect -759 -296 -747 296
rect -713 -296 -701 296
rect 701 296 759 346
rect -759 -346 -701 -296
rect 701 -296 713 296
rect 747 -296 759 296
rect 701 -346 759 -296
rect -759 -404 759 -346
<< mvpsubdiffcont >>
rect -747 -296 -713 296
rect 713 -296 747 296
<< poly >>
rect -567 244 -417 270
rect -239 244 -89 270
rect 89 244 239 270
rect 417 244 567 270
rect -567 -220 -417 -182
rect -567 -237 -509 -220
rect -525 -254 -509 -237
rect -475 -237 -417 -220
rect -239 -220 -89 -182
rect -239 -237 -181 -220
rect -475 -254 -459 -237
rect -525 -270 -459 -254
rect -197 -254 -181 -237
rect -147 -237 -89 -220
rect 89 -220 239 -182
rect 89 -237 147 -220
rect -147 -254 -131 -237
rect -197 -270 -131 -254
rect 131 -254 147 -237
rect 181 -237 239 -220
rect 417 -220 567 -182
rect 417 -237 475 -220
rect 181 -254 197 -237
rect 131 -270 197 -254
rect 459 -254 475 -237
rect 509 -237 567 -220
rect 509 -254 525 -237
rect 459 -270 525 -254
<< polycont >>
rect -509 -254 -475 -220
rect -181 -254 -147 -220
rect 147 -254 181 -220
rect 475 -254 509 -220
<< locali >>
rect -747 296 -713 312
rect 713 296 747 312
rect -613 232 -579 248
rect -613 -186 -579 -170
rect -405 232 -371 248
rect -405 -186 -371 -170
rect -285 232 -251 248
rect -285 -186 -251 -170
rect -77 232 -43 248
rect -77 -186 -43 -170
rect 43 232 77 248
rect 43 -186 77 -170
rect 251 232 285 248
rect 251 -186 285 -170
rect 371 232 405 248
rect 371 -186 405 -170
rect 579 232 613 248
rect 579 -186 613 -170
rect -525 -254 -509 -220
rect -475 -254 -459 -220
rect -197 -254 -181 -220
rect -147 -254 -131 -220
rect 131 -254 147 -220
rect 181 -254 197 -220
rect 459 -254 475 -220
rect 509 -254 525 -220
rect -747 -312 -713 -296
rect 713 -312 747 -296
<< viali >>
rect -613 -170 -579 232
rect -405 -170 -371 232
rect -285 -170 -251 232
rect -77 -170 -43 232
rect 43 -170 77 232
rect 251 -170 285 232
rect 371 -170 405 232
rect 579 -170 613 232
rect -509 -254 -475 -220
rect -181 -254 -147 -220
rect 147 -254 181 -220
rect 475 -254 509 -220
<< metal1 >>
rect -619 232 -573 244
rect -619 -170 -613 232
rect -579 -170 -573 232
rect -619 -182 -573 -170
rect -411 232 -365 244
rect -411 -170 -405 232
rect -371 -170 -365 232
rect -411 -182 -365 -170
rect -291 232 -245 244
rect -291 -170 -285 232
rect -251 -170 -245 232
rect -291 -182 -245 -170
rect -83 232 -37 244
rect -83 -170 -77 232
rect -43 -170 -37 232
rect -83 -182 -37 -170
rect 37 232 83 244
rect 37 -170 43 232
rect 77 -170 83 232
rect 37 -182 83 -170
rect 245 232 291 244
rect 245 -170 251 232
rect 285 -170 291 232
rect 245 -182 291 -170
rect 365 232 411 244
rect 365 -170 371 232
rect 405 -170 411 232
rect 365 -182 411 -170
rect 573 232 619 244
rect 573 -170 579 232
rect 613 -170 619 232
rect 573 -182 619 -170
rect -521 -220 -463 -214
rect -521 -254 -509 -220
rect -475 -254 -463 -220
rect -521 -260 -463 -254
rect -193 -220 -135 -214
rect -193 -254 -181 -220
rect -147 -254 -135 -220
rect -193 -260 -135 -254
rect 135 -220 193 -214
rect 135 -254 147 -220
rect 181 -254 193 -220
rect 135 -260 193 -254
rect 463 -220 521 -214
rect 463 -254 475 -220
rect 509 -254 521 -220
rect 463 -260 521 -254
<< properties >>
string FIXED_BBOX -730 -375 730 375
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.125 l 0.75 m 1 nf 4 diffcov 100 polycov 20 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
